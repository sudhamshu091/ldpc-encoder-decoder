module ldpc_encoder
  ( input  [1722:0] uncoded_block
  , output [2047:0] coded_block
  );
  wire _0 = uncoded_block[1] ^ uncoded_block[2];
  wire _1 = uncoded_block[3] ^ uncoded_block[4];
  wire _2 = _0 ^ _1;
  wire _3 = uncoded_block[5] ^ uncoded_block[7];
  wire _4 = uncoded_block[9] ^ uncoded_block[10];
  wire _5 = _3 ^ _4;
  wire _6 = _2 ^ _5;
  wire _7 = uncoded_block[11] ^ uncoded_block[12];
  wire _8 = uncoded_block[13] ^ uncoded_block[17];
  wire _9 = _7 ^ _8;
  wire _10 = uncoded_block[21] ^ uncoded_block[24];
  wire _11 = uncoded_block[30] ^ uncoded_block[31];
  wire _12 = _10 ^ _11;
  wire _13 = _9 ^ _12;
  wire _14 = _6 ^ _13;
  wire _15 = uncoded_block[32] ^ uncoded_block[33];
  wire _16 = uncoded_block[34] ^ uncoded_block[35];
  wire _17 = _15 ^ _16;
  wire _18 = uncoded_block[37] ^ uncoded_block[38];
  wire _19 = uncoded_block[39] ^ uncoded_block[40];
  wire _20 = _18 ^ _19;
  wire _21 = _17 ^ _20;
  wire _22 = uncoded_block[43] ^ uncoded_block[44];
  wire _23 = uncoded_block[45] ^ uncoded_block[46];
  wire _24 = _22 ^ _23;
  wire _25 = uncoded_block[53] ^ uncoded_block[56];
  wire _26 = uncoded_block[58] ^ uncoded_block[59];
  wire _27 = _25 ^ _26;
  wire _28 = _24 ^ _27;
  wire _29 = _21 ^ _28;
  wire _30 = _14 ^ _29;
  wire _31 = uncoded_block[60] ^ uncoded_block[62];
  wire _32 = uncoded_block[63] ^ uncoded_block[65];
  wire _33 = _31 ^ _32;
  wire _34 = uncoded_block[66] ^ uncoded_block[67];
  wire _35 = uncoded_block[68] ^ uncoded_block[69];
  wire _36 = _34 ^ _35;
  wire _37 = _33 ^ _36;
  wire _38 = uncoded_block[71] ^ uncoded_block[74];
  wire _39 = uncoded_block[76] ^ uncoded_block[77];
  wire _40 = _38 ^ _39;
  wire _41 = uncoded_block[82] ^ uncoded_block[83];
  wire _42 = uncoded_block[87] ^ uncoded_block[91];
  wire _43 = _41 ^ _42;
  wire _44 = _40 ^ _43;
  wire _45 = _37 ^ _44;
  wire _46 = uncoded_block[95] ^ uncoded_block[96];
  wire _47 = uncoded_block[97] ^ uncoded_block[98];
  wire _48 = _46 ^ _47;
  wire _49 = uncoded_block[101] ^ uncoded_block[103];
  wire _50 = uncoded_block[105] ^ uncoded_block[108];
  wire _51 = _49 ^ _50;
  wire _52 = _48 ^ _51;
  wire _53 = uncoded_block[109] ^ uncoded_block[114];
  wire _54 = uncoded_block[116] ^ uncoded_block[117];
  wire _55 = _53 ^ _54;
  wire _56 = uncoded_block[121] ^ uncoded_block[123];
  wire _57 = uncoded_block[127] ^ uncoded_block[129];
  wire _58 = _56 ^ _57;
  wire _59 = _55 ^ _58;
  wire _60 = _52 ^ _59;
  wire _61 = _45 ^ _60;
  wire _62 = _30 ^ _61;
  wire _63 = uncoded_block[132] ^ uncoded_block[136];
  wire _64 = uncoded_block[138] ^ uncoded_block[139];
  wire _65 = _63 ^ _64;
  wire _66 = uncoded_block[141] ^ uncoded_block[145];
  wire _67 = uncoded_block[146] ^ uncoded_block[148];
  wire _68 = _66 ^ _67;
  wire _69 = _65 ^ _68;
  wire _70 = uncoded_block[150] ^ uncoded_block[151];
  wire _71 = uncoded_block[152] ^ uncoded_block[154];
  wire _72 = _70 ^ _71;
  wire _73 = uncoded_block[157] ^ uncoded_block[158];
  wire _74 = uncoded_block[161] ^ uncoded_block[162];
  wire _75 = _73 ^ _74;
  wire _76 = _72 ^ _75;
  wire _77 = _69 ^ _76;
  wire _78 = uncoded_block[163] ^ uncoded_block[165];
  wire _79 = uncoded_block[167] ^ uncoded_block[168];
  wire _80 = _78 ^ _79;
  wire _81 = uncoded_block[170] ^ uncoded_block[172];
  wire _82 = uncoded_block[176] ^ uncoded_block[177];
  wire _83 = _81 ^ _82;
  wire _84 = _80 ^ _83;
  wire _85 = uncoded_block[178] ^ uncoded_block[179];
  wire _86 = uncoded_block[183] ^ uncoded_block[184];
  wire _87 = _85 ^ _86;
  wire _88 = uncoded_block[185] ^ uncoded_block[191];
  wire _89 = uncoded_block[193] ^ uncoded_block[194];
  wire _90 = _88 ^ _89;
  wire _91 = _87 ^ _90;
  wire _92 = _84 ^ _91;
  wire _93 = _77 ^ _92;
  wire _94 = uncoded_block[196] ^ uncoded_block[197];
  wire _95 = uncoded_block[200] ^ uncoded_block[202];
  wire _96 = _94 ^ _95;
  wire _97 = uncoded_block[208] ^ uncoded_block[209];
  wire _98 = uncoded_block[210] ^ uncoded_block[212];
  wire _99 = _97 ^ _98;
  wire _100 = _96 ^ _99;
  wire _101 = uncoded_block[215] ^ uncoded_block[217];
  wire _102 = uncoded_block[219] ^ uncoded_block[220];
  wire _103 = _101 ^ _102;
  wire _104 = uncoded_block[221] ^ uncoded_block[223];
  wire _105 = uncoded_block[224] ^ uncoded_block[226];
  wire _106 = _104 ^ _105;
  wire _107 = _103 ^ _106;
  wire _108 = _100 ^ _107;
  wire _109 = uncoded_block[227] ^ uncoded_block[228];
  wire _110 = uncoded_block[230] ^ uncoded_block[237];
  wire _111 = _109 ^ _110;
  wire _112 = uncoded_block[239] ^ uncoded_block[241];
  wire _113 = uncoded_block[242] ^ uncoded_block[244];
  wire _114 = _112 ^ _113;
  wire _115 = _111 ^ _114;
  wire _116 = uncoded_block[247] ^ uncoded_block[249];
  wire _117 = uncoded_block[252] ^ uncoded_block[257];
  wire _118 = _116 ^ _117;
  wire _119 = uncoded_block[259] ^ uncoded_block[260];
  wire _120 = uncoded_block[261] ^ uncoded_block[264];
  wire _121 = _119 ^ _120;
  wire _122 = _118 ^ _121;
  wire _123 = _115 ^ _122;
  wire _124 = _108 ^ _123;
  wire _125 = _93 ^ _124;
  wire _126 = _62 ^ _125;
  wire _127 = uncoded_block[267] ^ uncoded_block[269];
  wire _128 = uncoded_block[270] ^ uncoded_block[272];
  wire _129 = _127 ^ _128;
  wire _130 = uncoded_block[273] ^ uncoded_block[275];
  wire _131 = uncoded_block[278] ^ uncoded_block[284];
  wire _132 = _130 ^ _131;
  wire _133 = _129 ^ _132;
  wire _134 = uncoded_block[286] ^ uncoded_block[287];
  wire _135 = uncoded_block[288] ^ uncoded_block[290];
  wire _136 = _134 ^ _135;
  wire _137 = uncoded_block[295] ^ uncoded_block[296];
  wire _138 = uncoded_block[297] ^ uncoded_block[300];
  wire _139 = _137 ^ _138;
  wire _140 = _136 ^ _139;
  wire _141 = _133 ^ _140;
  wire _142 = uncoded_block[301] ^ uncoded_block[302];
  wire _143 = uncoded_block[303] ^ uncoded_block[306];
  wire _144 = _142 ^ _143;
  wire _145 = uncoded_block[313] ^ uncoded_block[314];
  wire _146 = uncoded_block[315] ^ uncoded_block[316];
  wire _147 = _145 ^ _146;
  wire _148 = _144 ^ _147;
  wire _149 = uncoded_block[317] ^ uncoded_block[319];
  wire _150 = uncoded_block[320] ^ uncoded_block[323];
  wire _151 = _149 ^ _150;
  wire _152 = uncoded_block[325] ^ uncoded_block[326];
  wire _153 = uncoded_block[328] ^ uncoded_block[335];
  wire _154 = _152 ^ _153;
  wire _155 = _151 ^ _154;
  wire _156 = _148 ^ _155;
  wire _157 = _141 ^ _156;
  wire _158 = uncoded_block[339] ^ uncoded_block[342];
  wire _159 = uncoded_block[345] ^ uncoded_block[346];
  wire _160 = _158 ^ _159;
  wire _161 = uncoded_block[347] ^ uncoded_block[349];
  wire _162 = uncoded_block[352] ^ uncoded_block[353];
  wire _163 = _161 ^ _162;
  wire _164 = _160 ^ _163;
  wire _165 = uncoded_block[354] ^ uncoded_block[358];
  wire _166 = uncoded_block[360] ^ uncoded_block[361];
  wire _167 = _165 ^ _166;
  wire _168 = uncoded_block[364] ^ uncoded_block[366];
  wire _169 = uncoded_block[369] ^ uncoded_block[371];
  wire _170 = _168 ^ _169;
  wire _171 = _167 ^ _170;
  wire _172 = _164 ^ _171;
  wire _173 = uncoded_block[373] ^ uncoded_block[376];
  wire _174 = uncoded_block[377] ^ uncoded_block[384];
  wire _175 = _173 ^ _174;
  wire _176 = uncoded_block[388] ^ uncoded_block[390];
  wire _177 = uncoded_block[393] ^ uncoded_block[395];
  wire _178 = _176 ^ _177;
  wire _179 = _175 ^ _178;
  wire _180 = uncoded_block[396] ^ uncoded_block[399];
  wire _181 = uncoded_block[400] ^ uncoded_block[401];
  wire _182 = _180 ^ _181;
  wire _183 = uncoded_block[402] ^ uncoded_block[404];
  wire _184 = uncoded_block[406] ^ uncoded_block[407];
  wire _185 = _183 ^ _184;
  wire _186 = _182 ^ _185;
  wire _187 = _179 ^ _186;
  wire _188 = _172 ^ _187;
  wire _189 = _157 ^ _188;
  wire _190 = uncoded_block[408] ^ uncoded_block[409];
  wire _191 = uncoded_block[410] ^ uncoded_block[413];
  wire _192 = _190 ^ _191;
  wire _193 = uncoded_block[416] ^ uncoded_block[418];
  wire _194 = uncoded_block[421] ^ uncoded_block[423];
  wire _195 = _193 ^ _194;
  wire _196 = _192 ^ _195;
  wire _197 = uncoded_block[425] ^ uncoded_block[427];
  wire _198 = uncoded_block[428] ^ uncoded_block[430];
  wire _199 = _197 ^ _198;
  wire _200 = uncoded_block[432] ^ uncoded_block[434];
  wire _201 = uncoded_block[435] ^ uncoded_block[437];
  wire _202 = _200 ^ _201;
  wire _203 = _199 ^ _202;
  wire _204 = _196 ^ _203;
  wire _205 = uncoded_block[441] ^ uncoded_block[442];
  wire _206 = uncoded_block[443] ^ uncoded_block[444];
  wire _207 = _205 ^ _206;
  wire _208 = uncoded_block[449] ^ uncoded_block[451];
  wire _209 = uncoded_block[452] ^ uncoded_block[454];
  wire _210 = _208 ^ _209;
  wire _211 = _207 ^ _210;
  wire _212 = uncoded_block[455] ^ uncoded_block[456];
  wire _213 = uncoded_block[457] ^ uncoded_block[458];
  wire _214 = _212 ^ _213;
  wire _215 = uncoded_block[459] ^ uncoded_block[464];
  wire _216 = uncoded_block[466] ^ uncoded_block[472];
  wire _217 = _215 ^ _216;
  wire _218 = _214 ^ _217;
  wire _219 = _211 ^ _218;
  wire _220 = _204 ^ _219;
  wire _221 = uncoded_block[473] ^ uncoded_block[475];
  wire _222 = uncoded_block[476] ^ uncoded_block[482];
  wire _223 = _221 ^ _222;
  wire _224 = uncoded_block[486] ^ uncoded_block[488];
  wire _225 = uncoded_block[490] ^ uncoded_block[495];
  wire _226 = _224 ^ _225;
  wire _227 = _223 ^ _226;
  wire _228 = uncoded_block[499] ^ uncoded_block[500];
  wire _229 = uncoded_block[502] ^ uncoded_block[504];
  wire _230 = _228 ^ _229;
  wire _231 = uncoded_block[508] ^ uncoded_block[510];
  wire _232 = uncoded_block[514] ^ uncoded_block[515];
  wire _233 = _231 ^ _232;
  wire _234 = _230 ^ _233;
  wire _235 = _227 ^ _234;
  wire _236 = uncoded_block[516] ^ uncoded_block[519];
  wire _237 = uncoded_block[521] ^ uncoded_block[523];
  wire _238 = _236 ^ _237;
  wire _239 = uncoded_block[524] ^ uncoded_block[528];
  wire _240 = uncoded_block[530] ^ uncoded_block[533];
  wire _241 = _239 ^ _240;
  wire _242 = _238 ^ _241;
  wire _243 = uncoded_block[535] ^ uncoded_block[537];
  wire _244 = uncoded_block[543] ^ uncoded_block[545];
  wire _245 = _243 ^ _244;
  wire _246 = uncoded_block[546] ^ uncoded_block[549];
  wire _247 = uncoded_block[550] ^ uncoded_block[551];
  wire _248 = _246 ^ _247;
  wire _249 = _245 ^ _248;
  wire _250 = _242 ^ _249;
  wire _251 = _235 ^ _250;
  wire _252 = _220 ^ _251;
  wire _253 = _189 ^ _252;
  wire _254 = _126 ^ _253;
  wire _255 = uncoded_block[552] ^ uncoded_block[557];
  wire _256 = uncoded_block[558] ^ uncoded_block[560];
  wire _257 = _255 ^ _256;
  wire _258 = uncoded_block[562] ^ uncoded_block[564];
  wire _259 = uncoded_block[566] ^ uncoded_block[570];
  wire _260 = _258 ^ _259;
  wire _261 = _257 ^ _260;
  wire _262 = uncoded_block[573] ^ uncoded_block[574];
  wire _263 = uncoded_block[577] ^ uncoded_block[578];
  wire _264 = _262 ^ _263;
  wire _265 = uncoded_block[579] ^ uncoded_block[581];
  wire _266 = uncoded_block[584] ^ uncoded_block[585];
  wire _267 = _265 ^ _266;
  wire _268 = _264 ^ _267;
  wire _269 = _261 ^ _268;
  wire _270 = uncoded_block[586] ^ uncoded_block[587];
  wire _271 = uncoded_block[588] ^ uncoded_block[591];
  wire _272 = _270 ^ _271;
  wire _273 = uncoded_block[592] ^ uncoded_block[596];
  wire _274 = uncoded_block[599] ^ uncoded_block[603];
  wire _275 = _273 ^ _274;
  wire _276 = _272 ^ _275;
  wire _277 = uncoded_block[606] ^ uncoded_block[607];
  wire _278 = uncoded_block[608] ^ uncoded_block[610];
  wire _279 = _277 ^ _278;
  wire _280 = uncoded_block[613] ^ uncoded_block[616];
  wire _281 = uncoded_block[617] ^ uncoded_block[619];
  wire _282 = _280 ^ _281;
  wire _283 = _279 ^ _282;
  wire _284 = _276 ^ _283;
  wire _285 = _269 ^ _284;
  wire _286 = uncoded_block[621] ^ uncoded_block[625];
  wire _287 = uncoded_block[626] ^ uncoded_block[628];
  wire _288 = _286 ^ _287;
  wire _289 = uncoded_block[629] ^ uncoded_block[632];
  wire _290 = uncoded_block[633] ^ uncoded_block[635];
  wire _291 = _289 ^ _290;
  wire _292 = _288 ^ _291;
  wire _293 = uncoded_block[636] ^ uncoded_block[639];
  wire _294 = uncoded_block[641] ^ uncoded_block[643];
  wire _295 = _293 ^ _294;
  wire _296 = uncoded_block[645] ^ uncoded_block[646];
  wire _297 = uncoded_block[648] ^ uncoded_block[649];
  wire _298 = _296 ^ _297;
  wire _299 = _295 ^ _298;
  wire _300 = _292 ^ _299;
  wire _301 = uncoded_block[650] ^ uncoded_block[651];
  wire _302 = uncoded_block[652] ^ uncoded_block[653];
  wire _303 = _301 ^ _302;
  wire _304 = uncoded_block[654] ^ uncoded_block[655];
  wire _305 = uncoded_block[657] ^ uncoded_block[659];
  wire _306 = _304 ^ _305;
  wire _307 = _303 ^ _306;
  wire _308 = uncoded_block[663] ^ uncoded_block[664];
  wire _309 = uncoded_block[666] ^ uncoded_block[667];
  wire _310 = _308 ^ _309;
  wire _311 = uncoded_block[669] ^ uncoded_block[670];
  wire _312 = uncoded_block[671] ^ uncoded_block[672];
  wire _313 = _311 ^ _312;
  wire _314 = _310 ^ _313;
  wire _315 = _307 ^ _314;
  wire _316 = _300 ^ _315;
  wire _317 = _285 ^ _316;
  wire _318 = uncoded_block[673] ^ uncoded_block[678];
  wire _319 = uncoded_block[680] ^ uncoded_block[682];
  wire _320 = _318 ^ _319;
  wire _321 = uncoded_block[684] ^ uncoded_block[685];
  wire _322 = uncoded_block[686] ^ uncoded_block[688];
  wire _323 = _321 ^ _322;
  wire _324 = _320 ^ _323;
  wire _325 = uncoded_block[689] ^ uncoded_block[690];
  wire _326 = uncoded_block[691] ^ uncoded_block[692];
  wire _327 = _325 ^ _326;
  wire _328 = uncoded_block[694] ^ uncoded_block[695];
  wire _329 = uncoded_block[696] ^ uncoded_block[699];
  wire _330 = _328 ^ _329;
  wire _331 = _327 ^ _330;
  wire _332 = _324 ^ _331;
  wire _333 = uncoded_block[700] ^ uncoded_block[701];
  wire _334 = uncoded_block[702] ^ uncoded_block[705];
  wire _335 = _333 ^ _334;
  wire _336 = uncoded_block[706] ^ uncoded_block[708];
  wire _337 = uncoded_block[712] ^ uncoded_block[714];
  wire _338 = _336 ^ _337;
  wire _339 = _335 ^ _338;
  wire _340 = uncoded_block[718] ^ uncoded_block[719];
  wire _341 = uncoded_block[720] ^ uncoded_block[721];
  wire _342 = _340 ^ _341;
  wire _343 = uncoded_block[722] ^ uncoded_block[723];
  wire _344 = uncoded_block[726] ^ uncoded_block[727];
  wire _345 = _343 ^ _344;
  wire _346 = _342 ^ _345;
  wire _347 = _339 ^ _346;
  wire _348 = _332 ^ _347;
  wire _349 = uncoded_block[731] ^ uncoded_block[734];
  wire _350 = uncoded_block[737] ^ uncoded_block[739];
  wire _351 = _349 ^ _350;
  wire _352 = uncoded_block[740] ^ uncoded_block[741];
  wire _353 = uncoded_block[744] ^ uncoded_block[746];
  wire _354 = _352 ^ _353;
  wire _355 = _351 ^ _354;
  wire _356 = uncoded_block[747] ^ uncoded_block[749];
  wire _357 = uncoded_block[750] ^ uncoded_block[756];
  wire _358 = _356 ^ _357;
  wire _359 = uncoded_block[758] ^ uncoded_block[759];
  wire _360 = uncoded_block[760] ^ uncoded_block[762];
  wire _361 = _359 ^ _360;
  wire _362 = _358 ^ _361;
  wire _363 = _355 ^ _362;
  wire _364 = uncoded_block[763] ^ uncoded_block[765];
  wire _365 = uncoded_block[766] ^ uncoded_block[767];
  wire _366 = _364 ^ _365;
  wire _367 = uncoded_block[768] ^ uncoded_block[774];
  wire _368 = uncoded_block[778] ^ uncoded_block[779];
  wire _369 = _367 ^ _368;
  wire _370 = _366 ^ _369;
  wire _371 = uncoded_block[785] ^ uncoded_block[786];
  wire _372 = uncoded_block[787] ^ uncoded_block[790];
  wire _373 = _371 ^ _372;
  wire _374 = uncoded_block[791] ^ uncoded_block[792];
  wire _375 = uncoded_block[794] ^ uncoded_block[795];
  wire _376 = _374 ^ _375;
  wire _377 = _373 ^ _376;
  wire _378 = _370 ^ _377;
  wire _379 = _363 ^ _378;
  wire _380 = _348 ^ _379;
  wire _381 = _317 ^ _380;
  wire _382 = uncoded_block[796] ^ uncoded_block[797];
  wire _383 = uncoded_block[798] ^ uncoded_block[799];
  wire _384 = _382 ^ _383;
  wire _385 = uncoded_block[800] ^ uncoded_block[801];
  wire _386 = uncoded_block[802] ^ uncoded_block[803];
  wire _387 = _385 ^ _386;
  wire _388 = _384 ^ _387;
  wire _389 = uncoded_block[804] ^ uncoded_block[805];
  wire _390 = uncoded_block[806] ^ uncoded_block[808];
  wire _391 = _389 ^ _390;
  wire _392 = uncoded_block[809] ^ uncoded_block[810];
  wire _393 = uncoded_block[815] ^ uncoded_block[818];
  wire _394 = _392 ^ _393;
  wire _395 = _391 ^ _394;
  wire _396 = _388 ^ _395;
  wire _397 = uncoded_block[821] ^ uncoded_block[823];
  wire _398 = uncoded_block[826] ^ uncoded_block[830];
  wire _399 = _397 ^ _398;
  wire _400 = uncoded_block[831] ^ uncoded_block[832];
  wire _401 = uncoded_block[835] ^ uncoded_block[836];
  wire _402 = _400 ^ _401;
  wire _403 = _399 ^ _402;
  wire _404 = uncoded_block[838] ^ uncoded_block[844];
  wire _405 = uncoded_block[845] ^ uncoded_block[848];
  wire _406 = _404 ^ _405;
  wire _407 = uncoded_block[850] ^ uncoded_block[857];
  wire _408 = uncoded_block[858] ^ uncoded_block[860];
  wire _409 = _407 ^ _408;
  wire _410 = _406 ^ _409;
  wire _411 = _403 ^ _410;
  wire _412 = _396 ^ _411;
  wire _413 = uncoded_block[862] ^ uncoded_block[863];
  wire _414 = uncoded_block[865] ^ uncoded_block[866];
  wire _415 = _413 ^ _414;
  wire _416 = uncoded_block[871] ^ uncoded_block[872];
  wire _417 = uncoded_block[874] ^ uncoded_block[875];
  wire _418 = _416 ^ _417;
  wire _419 = _415 ^ _418;
  wire _420 = uncoded_block[877] ^ uncoded_block[879];
  wire _421 = uncoded_block[880] ^ uncoded_block[882];
  wire _422 = _420 ^ _421;
  wire _423 = uncoded_block[884] ^ uncoded_block[885];
  wire _424 = uncoded_block[886] ^ uncoded_block[894];
  wire _425 = _423 ^ _424;
  wire _426 = _422 ^ _425;
  wire _427 = _419 ^ _426;
  wire _428 = uncoded_block[897] ^ uncoded_block[898];
  wire _429 = uncoded_block[900] ^ uncoded_block[901];
  wire _430 = _428 ^ _429;
  wire _431 = uncoded_block[905] ^ uncoded_block[907];
  wire _432 = uncoded_block[908] ^ uncoded_block[910];
  wire _433 = _431 ^ _432;
  wire _434 = _430 ^ _433;
  wire _435 = uncoded_block[911] ^ uncoded_block[913];
  wire _436 = uncoded_block[914] ^ uncoded_block[916];
  wire _437 = _435 ^ _436;
  wire _438 = uncoded_block[917] ^ uncoded_block[919];
  wire _439 = uncoded_block[920] ^ uncoded_block[921];
  wire _440 = _438 ^ _439;
  wire _441 = _437 ^ _440;
  wire _442 = _434 ^ _441;
  wire _443 = _427 ^ _442;
  wire _444 = _412 ^ _443;
  wire _445 = uncoded_block[922] ^ uncoded_block[923];
  wire _446 = uncoded_block[927] ^ uncoded_block[928];
  wire _447 = _445 ^ _446;
  wire _448 = uncoded_block[930] ^ uncoded_block[931];
  wire _449 = uncoded_block[933] ^ uncoded_block[935];
  wire _450 = _448 ^ _449;
  wire _451 = _447 ^ _450;
  wire _452 = uncoded_block[937] ^ uncoded_block[938];
  wire _453 = uncoded_block[940] ^ uncoded_block[941];
  wire _454 = _452 ^ _453;
  wire _455 = uncoded_block[943] ^ uncoded_block[945];
  wire _456 = uncoded_block[946] ^ uncoded_block[947];
  wire _457 = _455 ^ _456;
  wire _458 = _454 ^ _457;
  wire _459 = _451 ^ _458;
  wire _460 = uncoded_block[948] ^ uncoded_block[950];
  wire _461 = uncoded_block[954] ^ uncoded_block[955];
  wire _462 = _460 ^ _461;
  wire _463 = uncoded_block[956] ^ uncoded_block[959];
  wire _464 = uncoded_block[960] ^ uncoded_block[963];
  wire _465 = _463 ^ _464;
  wire _466 = _462 ^ _465;
  wire _467 = uncoded_block[967] ^ uncoded_block[970];
  wire _468 = uncoded_block[971] ^ uncoded_block[972];
  wire _469 = _467 ^ _468;
  wire _470 = uncoded_block[974] ^ uncoded_block[975];
  wire _471 = uncoded_block[977] ^ uncoded_block[979];
  wire _472 = _470 ^ _471;
  wire _473 = _469 ^ _472;
  wire _474 = _466 ^ _473;
  wire _475 = _459 ^ _474;
  wire _476 = uncoded_block[981] ^ uncoded_block[982];
  wire _477 = uncoded_block[985] ^ uncoded_block[991];
  wire _478 = _476 ^ _477;
  wire _479 = uncoded_block[994] ^ uncoded_block[995];
  wire _480 = uncoded_block[996] ^ uncoded_block[998];
  wire _481 = _479 ^ _480;
  wire _482 = _478 ^ _481;
  wire _483 = uncoded_block[1001] ^ uncoded_block[1003];
  wire _484 = uncoded_block[1004] ^ uncoded_block[1005];
  wire _485 = _483 ^ _484;
  wire _486 = uncoded_block[1006] ^ uncoded_block[1008];
  wire _487 = uncoded_block[1009] ^ uncoded_block[1011];
  wire _488 = _486 ^ _487;
  wire _489 = _485 ^ _488;
  wire _490 = _482 ^ _489;
  wire _491 = uncoded_block[1012] ^ uncoded_block[1014];
  wire _492 = uncoded_block[1016] ^ uncoded_block[1018];
  wire _493 = _491 ^ _492;
  wire _494 = uncoded_block[1019] ^ uncoded_block[1023];
  wire _495 = uncoded_block[1025] ^ uncoded_block[1026];
  wire _496 = _494 ^ _495;
  wire _497 = _493 ^ _496;
  wire _498 = uncoded_block[1027] ^ uncoded_block[1028];
  wire _499 = uncoded_block[1031] ^ uncoded_block[1032];
  wire _500 = _498 ^ _499;
  wire _501 = uncoded_block[1034] ^ uncoded_block[1035];
  wire _502 = uncoded_block[1036] ^ uncoded_block[1038];
  wire _503 = _501 ^ _502;
  wire _504 = _500 ^ _503;
  wire _505 = _497 ^ _504;
  wire _506 = _490 ^ _505;
  wire _507 = _475 ^ _506;
  wire _508 = _444 ^ _507;
  wire _509 = _381 ^ _508;
  wire _510 = _254 ^ _509;
  wire _511 = uncoded_block[1039] ^ uncoded_block[1041];
  wire _512 = uncoded_block[1042] ^ uncoded_block[1043];
  wire _513 = _511 ^ _512;
  wire _514 = uncoded_block[1044] ^ uncoded_block[1045];
  wire _515 = uncoded_block[1047] ^ uncoded_block[1048];
  wire _516 = _514 ^ _515;
  wire _517 = _513 ^ _516;
  wire _518 = uncoded_block[1050] ^ uncoded_block[1051];
  wire _519 = uncoded_block[1056] ^ uncoded_block[1057];
  wire _520 = _518 ^ _519;
  wire _521 = uncoded_block[1059] ^ uncoded_block[1061];
  wire _522 = uncoded_block[1062] ^ uncoded_block[1063];
  wire _523 = _521 ^ _522;
  wire _524 = _520 ^ _523;
  wire _525 = _517 ^ _524;
  wire _526 = uncoded_block[1065] ^ uncoded_block[1068];
  wire _527 = uncoded_block[1071] ^ uncoded_block[1072];
  wire _528 = _526 ^ _527;
  wire _529 = uncoded_block[1074] ^ uncoded_block[1076];
  wire _530 = uncoded_block[1080] ^ uncoded_block[1081];
  wire _531 = _529 ^ _530;
  wire _532 = _528 ^ _531;
  wire _533 = uncoded_block[1083] ^ uncoded_block[1084];
  wire _534 = uncoded_block[1085] ^ uncoded_block[1088];
  wire _535 = _533 ^ _534;
  wire _536 = uncoded_block[1090] ^ uncoded_block[1092];
  wire _537 = uncoded_block[1093] ^ uncoded_block[1094];
  wire _538 = _536 ^ _537;
  wire _539 = _535 ^ _538;
  wire _540 = _532 ^ _539;
  wire _541 = _525 ^ _540;
  wire _542 = uncoded_block[1095] ^ uncoded_block[1096];
  wire _543 = uncoded_block[1098] ^ uncoded_block[1099];
  wire _544 = _542 ^ _543;
  wire _545 = uncoded_block[1100] ^ uncoded_block[1101];
  wire _546 = uncoded_block[1102] ^ uncoded_block[1105];
  wire _547 = _545 ^ _546;
  wire _548 = _544 ^ _547;
  wire _549 = uncoded_block[1107] ^ uncoded_block[1108];
  wire _550 = uncoded_block[1109] ^ uncoded_block[1111];
  wire _551 = _549 ^ _550;
  wire _552 = uncoded_block[1112] ^ uncoded_block[1115];
  wire _553 = uncoded_block[1116] ^ uncoded_block[1119];
  wire _554 = _552 ^ _553;
  wire _555 = _551 ^ _554;
  wire _556 = _548 ^ _555;
  wire _557 = uncoded_block[1121] ^ uncoded_block[1124];
  wire _558 = uncoded_block[1126] ^ uncoded_block[1129];
  wire _559 = _557 ^ _558;
  wire _560 = uncoded_block[1130] ^ uncoded_block[1131];
  wire _561 = uncoded_block[1132] ^ uncoded_block[1133];
  wire _562 = _560 ^ _561;
  wire _563 = _559 ^ _562;
  wire _564 = uncoded_block[1135] ^ uncoded_block[1137];
  wire _565 = uncoded_block[1138] ^ uncoded_block[1139];
  wire _566 = _564 ^ _565;
  wire _567 = uncoded_block[1140] ^ uncoded_block[1141];
  wire _568 = uncoded_block[1142] ^ uncoded_block[1143];
  wire _569 = _567 ^ _568;
  wire _570 = _566 ^ _569;
  wire _571 = _563 ^ _570;
  wire _572 = _556 ^ _571;
  wire _573 = _541 ^ _572;
  wire _574 = uncoded_block[1144] ^ uncoded_block[1146];
  wire _575 = uncoded_block[1147] ^ uncoded_block[1151];
  wire _576 = _574 ^ _575;
  wire _577 = uncoded_block[1152] ^ uncoded_block[1154];
  wire _578 = uncoded_block[1158] ^ uncoded_block[1159];
  wire _579 = _577 ^ _578;
  wire _580 = _576 ^ _579;
  wire _581 = uncoded_block[1160] ^ uncoded_block[1162];
  wire _582 = uncoded_block[1163] ^ uncoded_block[1167];
  wire _583 = _581 ^ _582;
  wire _584 = uncoded_block[1170] ^ uncoded_block[1174];
  wire _585 = uncoded_block[1175] ^ uncoded_block[1176];
  wire _586 = _584 ^ _585;
  wire _587 = _583 ^ _586;
  wire _588 = _580 ^ _587;
  wire _589 = uncoded_block[1177] ^ uncoded_block[1178];
  wire _590 = uncoded_block[1180] ^ uncoded_block[1181];
  wire _591 = _589 ^ _590;
  wire _592 = uncoded_block[1182] ^ uncoded_block[1183];
  wire _593 = uncoded_block[1187] ^ uncoded_block[1191];
  wire _594 = _592 ^ _593;
  wire _595 = _591 ^ _594;
  wire _596 = uncoded_block[1193] ^ uncoded_block[1195];
  wire _597 = uncoded_block[1196] ^ uncoded_block[1198];
  wire _598 = _596 ^ _597;
  wire _599 = uncoded_block[1199] ^ uncoded_block[1201];
  wire _600 = uncoded_block[1205] ^ uncoded_block[1214];
  wire _601 = _599 ^ _600;
  wire _602 = _598 ^ _601;
  wire _603 = _595 ^ _602;
  wire _604 = _588 ^ _603;
  wire _605 = uncoded_block[1216] ^ uncoded_block[1217];
  wire _606 = uncoded_block[1218] ^ uncoded_block[1219];
  wire _607 = _605 ^ _606;
  wire _608 = uncoded_block[1220] ^ uncoded_block[1222];
  wire _609 = uncoded_block[1223] ^ uncoded_block[1224];
  wire _610 = _608 ^ _609;
  wire _611 = _607 ^ _610;
  wire _612 = uncoded_block[1226] ^ uncoded_block[1227];
  wire _613 = uncoded_block[1228] ^ uncoded_block[1231];
  wire _614 = _612 ^ _613;
  wire _615 = uncoded_block[1232] ^ uncoded_block[1236];
  wire _616 = uncoded_block[1237] ^ uncoded_block[1242];
  wire _617 = _615 ^ _616;
  wire _618 = _614 ^ _617;
  wire _619 = _611 ^ _618;
  wire _620 = uncoded_block[1243] ^ uncoded_block[1247];
  wire _621 = uncoded_block[1249] ^ uncoded_block[1251];
  wire _622 = _620 ^ _621;
  wire _623 = uncoded_block[1252] ^ uncoded_block[1255];
  wire _624 = uncoded_block[1257] ^ uncoded_block[1260];
  wire _625 = _623 ^ _624;
  wire _626 = _622 ^ _625;
  wire _627 = uncoded_block[1265] ^ uncoded_block[1266];
  wire _628 = uncoded_block[1271] ^ uncoded_block[1272];
  wire _629 = _627 ^ _628;
  wire _630 = uncoded_block[1275] ^ uncoded_block[1277];
  wire _631 = uncoded_block[1279] ^ uncoded_block[1280];
  wire _632 = _630 ^ _631;
  wire _633 = _629 ^ _632;
  wire _634 = _626 ^ _633;
  wire _635 = _619 ^ _634;
  wire _636 = _604 ^ _635;
  wire _637 = _573 ^ _636;
  wire _638 = uncoded_block[1283] ^ uncoded_block[1284];
  wire _639 = uncoded_block[1286] ^ uncoded_block[1287];
  wire _640 = _638 ^ _639;
  wire _641 = uncoded_block[1289] ^ uncoded_block[1291];
  wire _642 = uncoded_block[1292] ^ uncoded_block[1295];
  wire _643 = _641 ^ _642;
  wire _644 = _640 ^ _643;
  wire _645 = uncoded_block[1296] ^ uncoded_block[1298];
  wire _646 = uncoded_block[1300] ^ uncoded_block[1302];
  wire _647 = _645 ^ _646;
  wire _648 = uncoded_block[1305] ^ uncoded_block[1306];
  wire _649 = uncoded_block[1307] ^ uncoded_block[1309];
  wire _650 = _648 ^ _649;
  wire _651 = _647 ^ _650;
  wire _652 = _644 ^ _651;
  wire _653 = uncoded_block[1310] ^ uncoded_block[1316];
  wire _654 = uncoded_block[1319] ^ uncoded_block[1321];
  wire _655 = _653 ^ _654;
  wire _656 = uncoded_block[1325] ^ uncoded_block[1326];
  wire _657 = uncoded_block[1327] ^ uncoded_block[1330];
  wire _658 = _656 ^ _657;
  wire _659 = _655 ^ _658;
  wire _660 = uncoded_block[1331] ^ uncoded_block[1334];
  wire _661 = uncoded_block[1335] ^ uncoded_block[1337];
  wire _662 = _660 ^ _661;
  wire _663 = uncoded_block[1338] ^ uncoded_block[1343];
  wire _664 = uncoded_block[1346] ^ uncoded_block[1347];
  wire _665 = _663 ^ _664;
  wire _666 = _662 ^ _665;
  wire _667 = _659 ^ _666;
  wire _668 = _652 ^ _667;
  wire _669 = uncoded_block[1348] ^ uncoded_block[1349];
  wire _670 = uncoded_block[1351] ^ uncoded_block[1352];
  wire _671 = _669 ^ _670;
  wire _672 = uncoded_block[1353] ^ uncoded_block[1355];
  wire _673 = uncoded_block[1356] ^ uncoded_block[1358];
  wire _674 = _672 ^ _673;
  wire _675 = _671 ^ _674;
  wire _676 = uncoded_block[1359] ^ uncoded_block[1362];
  wire _677 = uncoded_block[1363] ^ uncoded_block[1364];
  wire _678 = _676 ^ _677;
  wire _679 = uncoded_block[1365] ^ uncoded_block[1367];
  wire _680 = uncoded_block[1369] ^ uncoded_block[1371];
  wire _681 = _679 ^ _680;
  wire _682 = _678 ^ _681;
  wire _683 = _675 ^ _682;
  wire _684 = uncoded_block[1372] ^ uncoded_block[1373];
  wire _685 = uncoded_block[1374] ^ uncoded_block[1378];
  wire _686 = _684 ^ _685;
  wire _687 = uncoded_block[1381] ^ uncoded_block[1383];
  wire _688 = uncoded_block[1385] ^ uncoded_block[1387];
  wire _689 = _687 ^ _688;
  wire _690 = _686 ^ _689;
  wire _691 = uncoded_block[1388] ^ uncoded_block[1389];
  wire _692 = uncoded_block[1390] ^ uncoded_block[1393];
  wire _693 = _691 ^ _692;
  wire _694 = uncoded_block[1394] ^ uncoded_block[1395];
  wire _695 = uncoded_block[1397] ^ uncoded_block[1402];
  wire _696 = _694 ^ _695;
  wire _697 = _693 ^ _696;
  wire _698 = _690 ^ _697;
  wire _699 = _683 ^ _698;
  wire _700 = _668 ^ _699;
  wire _701 = uncoded_block[1406] ^ uncoded_block[1408];
  wire _702 = uncoded_block[1411] ^ uncoded_block[1413];
  wire _703 = _701 ^ _702;
  wire _704 = uncoded_block[1414] ^ uncoded_block[1416];
  wire _705 = uncoded_block[1417] ^ uncoded_block[1418];
  wire _706 = _704 ^ _705;
  wire _707 = _703 ^ _706;
  wire _708 = uncoded_block[1420] ^ uncoded_block[1423];
  wire _709 = uncoded_block[1424] ^ uncoded_block[1425];
  wire _710 = _708 ^ _709;
  wire _711 = uncoded_block[1427] ^ uncoded_block[1436];
  wire _712 = uncoded_block[1437] ^ uncoded_block[1440];
  wire _713 = _711 ^ _712;
  wire _714 = _710 ^ _713;
  wire _715 = _707 ^ _714;
  wire _716 = uncoded_block[1443] ^ uncoded_block[1445];
  wire _717 = uncoded_block[1447] ^ uncoded_block[1449];
  wire _718 = _716 ^ _717;
  wire _719 = uncoded_block[1452] ^ uncoded_block[1453];
  wire _720 = uncoded_block[1454] ^ uncoded_block[1456];
  wire _721 = _719 ^ _720;
  wire _722 = _718 ^ _721;
  wire _723 = uncoded_block[1457] ^ uncoded_block[1458];
  wire _724 = uncoded_block[1459] ^ uncoded_block[1460];
  wire _725 = _723 ^ _724;
  wire _726 = uncoded_block[1461] ^ uncoded_block[1462];
  wire _727 = uncoded_block[1466] ^ uncoded_block[1467];
  wire _728 = _726 ^ _727;
  wire _729 = _725 ^ _728;
  wire _730 = _722 ^ _729;
  wire _731 = _715 ^ _730;
  wire _732 = uncoded_block[1469] ^ uncoded_block[1471];
  wire _733 = uncoded_block[1474] ^ uncoded_block[1475];
  wire _734 = _732 ^ _733;
  wire _735 = uncoded_block[1476] ^ uncoded_block[1477];
  wire _736 = uncoded_block[1478] ^ uncoded_block[1482];
  wire _737 = _735 ^ _736;
  wire _738 = _734 ^ _737;
  wire _739 = uncoded_block[1486] ^ uncoded_block[1487];
  wire _740 = uncoded_block[1488] ^ uncoded_block[1489];
  wire _741 = _739 ^ _740;
  wire _742 = uncoded_block[1490] ^ uncoded_block[1495];
  wire _743 = uncoded_block[1496] ^ uncoded_block[1497];
  wire _744 = _742 ^ _743;
  wire _745 = _741 ^ _744;
  wire _746 = _738 ^ _745;
  wire _747 = uncoded_block[1499] ^ uncoded_block[1500];
  wire _748 = uncoded_block[1501] ^ uncoded_block[1506];
  wire _749 = _747 ^ _748;
  wire _750 = uncoded_block[1509] ^ uncoded_block[1511];
  wire _751 = uncoded_block[1514] ^ uncoded_block[1517];
  //https://github.com/bigdot123456/LPDC5G
  wire _752 = _750 ^ _751;
  wire _753 = _749 ^ _752;
  wire _754 = uncoded_block[1518] ^ uncoded_block[1520];
  wire _755 = uncoded_block[1523] ^ uncoded_block[1525];
  wire _756 = _754 ^ _755;
  wire _757 = uncoded_block[1529] ^ uncoded_block[1538];
  wire _758 = uncoded_block[1539] ^ uncoded_block[1541];
  wire _759 = _757 ^ _758;
  wire _760 = _756 ^ _759;
  wire _761 = _753 ^ _760;
  wire _762 = _746 ^ _761;
  wire _763 = _731 ^ _762;
  wire _764 = _700 ^ _763;
  wire _765 = _637 ^ _764;
  wire _766 = uncoded_block[1547] ^ uncoded_block[1550];
  wire _767 = uncoded_block[1551] ^ uncoded_block[1552];
  wire _768 = _766 ^ _767;
  wire _769 = uncoded_block[1553] ^ uncoded_block[1554];
  wire _770 = uncoded_block[1555] ^ uncoded_block[1557];
  wire _771 = _769 ^ _770;
  wire _772 = _768 ^ _771;
  wire _773 = uncoded_block[1558] ^ uncoded_block[1560];
  wire _774 = uncoded_block[1561] ^ uncoded_block[1562];
  wire _775 = _773 ^ _774;
  wire _776 = uncoded_block[1563] ^ uncoded_block[1565];
  wire _777 = uncoded_block[1566] ^ uncoded_block[1570];
  wire _778 = _776 ^ _777;
  wire _779 = _775 ^ _778;
  wire _780 = _772 ^ _779;
  wire _781 = uncoded_block[1574] ^ uncoded_block[1575];
  wire _782 = uncoded_block[1576] ^ uncoded_block[1577];
  wire _783 = _781 ^ _782;
  wire _784 = uncoded_block[1580] ^ uncoded_block[1581];
  wire _785 = uncoded_block[1583] ^ uncoded_block[1584];
  wire _786 = _784 ^ _785;
  wire _787 = _783 ^ _786;
  wire _788 = uncoded_block[1585] ^ uncoded_block[1587];
  wire _789 = uncoded_block[1589] ^ uncoded_block[1591];
  wire _790 = _788 ^ _789;
  wire _791 = uncoded_block[1592] ^ uncoded_block[1593];
  wire _792 = uncoded_block[1595] ^ uncoded_block[1596];
  wire _793 = _791 ^ _792;
  wire _794 = _790 ^ _793;
  wire _795 = _787 ^ _794;
  wire _796 = _780 ^ _795;
  wire _797 = uncoded_block[1598] ^ uncoded_block[1600];
  wire _798 = uncoded_block[1602] ^ uncoded_block[1604];
  wire _799 = _797 ^ _798;
  wire _800 = uncoded_block[1606] ^ uncoded_block[1607];
  wire _801 = uncoded_block[1611] ^ uncoded_block[1612];
  wire _802 = _800 ^ _801;
  wire _803 = _799 ^ _802;
  wire _804 = uncoded_block[1617] ^ uncoded_block[1618];
  wire _805 = uncoded_block[1619] ^ uncoded_block[1622];
  wire _806 = _804 ^ _805;
  wire _807 = uncoded_block[1625] ^ uncoded_block[1626];
  wire _808 = uncoded_block[1628] ^ uncoded_block[1630];
  wire _809 = _807 ^ _808;
  wire _810 = _806 ^ _809;
  wire _811 = _803 ^ _810;
  wire _812 = uncoded_block[1632] ^ uncoded_block[1633];
  wire _813 = uncoded_block[1634] ^ uncoded_block[1639];
  wire _814 = _812 ^ _813;
  wire _815 = uncoded_block[1642] ^ uncoded_block[1644];
  wire _816 = uncoded_block[1645] ^ uncoded_block[1646];
  wire _817 = _815 ^ _816;
  wire _818 = _814 ^ _817;
  wire _819 = uncoded_block[1648] ^ uncoded_block[1651];
  wire _820 = uncoded_block[1654] ^ uncoded_block[1656];
  wire _821 = _819 ^ _820;
  wire _822 = uncoded_block[1657] ^ uncoded_block[1659];
  wire _823 = uncoded_block[1661] ^ uncoded_block[1662];
  wire _824 = _822 ^ _823;
  wire _825 = _821 ^ _824;
  wire _826 = _818 ^ _825;
  wire _827 = _811 ^ _826;
  wire _828 = _796 ^ _827;
  wire _829 = uncoded_block[1663] ^ uncoded_block[1672];
  wire _830 = uncoded_block[1674] ^ uncoded_block[1675];
  wire _831 = _829 ^ _830;
  wire _832 = uncoded_block[1676] ^ uncoded_block[1678];
  wire _833 = uncoded_block[1679] ^ uncoded_block[1681];
  wire _834 = _832 ^ _833;
  wire _835 = _831 ^ _834;
  wire _836 = uncoded_block[1683] ^ uncoded_block[1687];
  wire _837 = uncoded_block[1688] ^ uncoded_block[1689];
  wire _838 = _836 ^ _837;
  wire _839 = uncoded_block[1690] ^ uncoded_block[1693];
  wire _840 = uncoded_block[1694] ^ uncoded_block[1695];
  wire _841 = _839 ^ _840;
  wire _842 = _838 ^ _841;
  wire _843 = _835 ^ _842;
  wire _844 = uncoded_block[1696] ^ uncoded_block[1699];
  wire _845 = uncoded_block[1700] ^ uncoded_block[1703];
  wire _846 = _844 ^ _845;
  wire _847 = uncoded_block[1704] ^ uncoded_block[1706];
  wire _848 = uncoded_block[1707] ^ uncoded_block[1708];
  wire _849 = _847 ^ _848;
  wire _850 = _846 ^ _849;
  wire _851 = uncoded_block[1709] ^ uncoded_block[1710];
  wire _852 = uncoded_block[1712] ^ uncoded_block[1713];
  wire _853 = _851 ^ _852;
  wire _854 = uncoded_block[1714] ^ uncoded_block[1715];
  wire _855 = uncoded_block[1716] ^ uncoded_block[1718];
  wire _856 = _854 ^ _855;
  wire _857 = _853 ^ _856;
  wire _858 = _850 ^ _857;
  wire _859 = _843 ^ _858;
  wire _860 = uncoded_block[1719] ^ uncoded_block[1720];
  wire _861 = _860 ^ uncoded_block[1721];
  wire _862 = _859 ^ _861;
  wire _863 = _828 ^ _862;
  wire _864 = _765 ^ _863;
  wire _865 = _510 ^ _864;
  wire _866 = uncoded_block[3] ^ uncoded_block[6];
  wire _867 = _866 ^ _4;
  wire _868 = uncoded_block[14] ^ uncoded_block[15];
  wire _869 = _7 ^ _868;
  wire _870 = _867 ^ _869;
  wire _871 = uncoded_block[16] ^ uncoded_block[17];
  wire _872 = uncoded_block[20] ^ uncoded_block[25];
  wire _873 = _871 ^ _872;
  wire _874 = uncoded_block[28] ^ uncoded_block[30];
  wire _875 = uncoded_block[31] ^ uncoded_block[32];
  wire _876 = _874 ^ _875;
  wire _877 = _873 ^ _876;
  wire _878 = _870 ^ _877;
  wire _879 = uncoded_block[35] ^ uncoded_block[36];
  wire _880 = uncoded_block[37] ^ uncoded_block[39];
  wire _881 = _879 ^ _880;
  wire _882 = uncoded_block[40] ^ uncoded_block[42];
  wire _883 = _882 ^ _23;
  wire _884 = _881 ^ _883;
  wire _885 = uncoded_block[47] ^ uncoded_block[49];
  wire _886 = uncoded_block[51] ^ uncoded_block[53];
  wire _887 = _885 ^ _886;
  wire _888 = uncoded_block[55] ^ uncoded_block[56];
  wire _889 = uncoded_block[58] ^ uncoded_block[60];
  wire _890 = _888 ^ _889;
  wire _891 = _887 ^ _890;
  wire _892 = _884 ^ _891;
  wire _893 = _878 ^ _892;
  wire _894 = uncoded_block[62] ^ uncoded_block[64];
  wire _895 = _894 ^ _34;
  wire _896 = uncoded_block[69] ^ uncoded_block[71];
  wire _897 = uncoded_block[72] ^ uncoded_block[73];
  wire _898 = _896 ^ _897;
  wire _899 = _895 ^ _898;
  wire _900 = uncoded_block[74] ^ uncoded_block[76];
  wire _901 = uncoded_block[77] ^ uncoded_block[78];
  wire _902 = _900 ^ _901;
  wire _903 = uncoded_block[90] ^ uncoded_block[91];
  wire _904 = _41 ^ _903;
  wire _905 = _902 ^ _904;
  wire _906 = _899 ^ _905;
  wire _907 = uncoded_block[92] ^ uncoded_block[93];
  wire _908 = uncoded_block[94] ^ uncoded_block[97];
  wire _909 = _907 ^ _908;
  wire _910 = uncoded_block[99] ^ uncoded_block[101];
  wire _911 = uncoded_block[106] ^ uncoded_block[108];
  wire _912 = _910 ^ _911;
  wire _913 = _909 ^ _912;
  wire _914 = uncoded_block[112] ^ uncoded_block[114];
  wire _915 = uncoded_block[115] ^ uncoded_block[117];
  wire _916 = _914 ^ _915;
  wire _917 = uncoded_block[126] ^ uncoded_block[128];
  wire _918 = _56 ^ _917;
  wire _919 = _916 ^ _918;
  wire _920 = _913 ^ _919;
  wire _921 = _906 ^ _920;
  wire _922 = _893 ^ _921;
  wire _923 = uncoded_block[129] ^ uncoded_block[130];
  wire _924 = uncoded_block[132] ^ uncoded_block[133];
  wire _925 = _923 ^ _924;
  wire _926 = uncoded_block[134] ^ uncoded_block[135];
  wire _927 = uncoded_block[137] ^ uncoded_block[140];
  wire _928 = _926 ^ _927;
  wire _929 = _925 ^ _928;
  wire _930 = uncoded_block[141] ^ uncoded_block[151];
  wire _931 = _930 ^ _71;
  wire _932 = uncoded_block[155] ^ uncoded_block[157];
  wire _933 = uncoded_block[159] ^ uncoded_block[164];
  wire _934 = _932 ^ _933;
  wire _935 = _931 ^ _934;
  wire _936 = _929 ^ _935;
  wire _937 = uncoded_block[165] ^ uncoded_block[171];
  wire _938 = uncoded_block[172] ^ uncoded_block[173];
  wire _939 = _937 ^ _938;
  wire _940 = uncoded_block[177] ^ uncoded_block[178];
  wire _941 = uncoded_block[180] ^ uncoded_block[182];
  wire _942 = _940 ^ _941;
  wire _943 = _939 ^ _942;
  wire _944 = uncoded_block[183] ^ uncoded_block[185];
  wire _945 = uncoded_block[187] ^ uncoded_block[188];
  wire _946 = _944 ^ _945;
  wire _947 = uncoded_block[189] ^ uncoded_block[191];
  wire _948 = _947 ^ _94;
  wire _949 = _946 ^ _948;
  wire _950 = _943 ^ _949;
  wire _951 = _936 ^ _950;
  wire _952 = uncoded_block[198] ^ uncoded_block[201];
  wire _953 = uncoded_block[202] ^ uncoded_block[206];
  wire _954 = _952 ^ _953;
  wire _955 = uncoded_block[209] ^ uncoded_block[210];
  wire _956 = uncoded_block[211] ^ uncoded_block[212];
  wire _957 = _955 ^ _956;
  wire _958 = _954 ^ _957;
  wire _959 = uncoded_block[213] ^ uncoded_block[214];
  wire _960 = uncoded_block[217] ^ uncoded_block[218];
  wire _961 = _959 ^ _960;
  wire _962 = uncoded_block[219] ^ uncoded_block[224];
  wire _963 = uncoded_block[225] ^ uncoded_block[231];
  wire _964 = _962 ^ _963;
  wire _965 = _961 ^ _964;
  wire _966 = _958 ^ _965;
  wire _967 = uncoded_block[232] ^ uncoded_block[233];
  wire _968 = uncoded_block[234] ^ uncoded_block[235];
  wire _969 = _967 ^ _968;
  wire _970 = uncoded_block[237] ^ uncoded_block[238];
  wire _971 = uncoded_block[243] ^ uncoded_block[246];
  wire _972 = _970 ^ _971;
  wire _973 = _969 ^ _972;
  wire _974 = uncoded_block[247] ^ uncoded_block[250];
  wire _975 = _974 ^ _117;
  wire _976 = uncoded_block[258] ^ uncoded_block[263];
  wire _977 = uncoded_block[264] ^ uncoded_block[265];
  wire _978 = _976 ^ _977;
  wire _979 = _975 ^ _978;
  wire _980 = _973 ^ _979;
  wire _981 = _966 ^ _980;
  wire _982 = _951 ^ _981;
  wire _983 = _922 ^ _982;
  wire _984 = uncoded_block[266] ^ uncoded_block[267];
  wire _985 = uncoded_block[268] ^ uncoded_block[269];
  wire _986 = _984 ^ _985;
  wire _987 = uncoded_block[271] ^ uncoded_block[280];
  wire _988 = uncoded_block[281] ^ uncoded_block[283];
  wire _989 = _987 ^ _988;
  wire _990 = _986 ^ _989;
  wire _991 = uncoded_block[285] ^ uncoded_block[287];
  wire _992 = uncoded_block[288] ^ uncoded_block[289];
  wire _993 = _991 ^ _992;
  wire _994 = uncoded_block[291] ^ uncoded_block[292];
  wire _995 = uncoded_block[293] ^ uncoded_block[294];
  wire _996 = _994 ^ _995;
  wire _997 = _993 ^ _996;
  wire _998 = _990 ^ _997;
  wire _999 = uncoded_block[300] ^ uncoded_block[303];
  wire _1000 = uncoded_block[304] ^ uncoded_block[305];
  wire _1001 = _999 ^ _1000;
  wire _1002 = uncoded_block[306] ^ uncoded_block[308];
  wire _1003 = uncoded_block[310] ^ uncoded_block[312];
  wire _1004 = _1002 ^ _1003;
  wire _1005 = _1001 ^ _1004;
  wire _1006 = uncoded_block[315] ^ uncoded_block[317];
  wire _1007 = _145 ^ _1006;
  wire _1008 = uncoded_block[319] ^ uncoded_block[320];
  wire _1009 = uncoded_block[321] ^ uncoded_block[324];
  wire _1010 = _1008 ^ _1009;
  wire _1011 = _1007 ^ _1010;
  wire _1012 = _1005 ^ _1011;
  wire _1013 = _998 ^ _1012;
  wire _1014 = uncoded_block[326] ^ uncoded_block[327];
  wire _1015 = uncoded_block[329] ^ uncoded_block[332];
  wire _1016 = _1014 ^ _1015;
  wire _1017 = uncoded_block[334] ^ uncoded_block[336];
  wire _1018 = uncoded_block[337] ^ uncoded_block[340];
  wire _1019 = _1017 ^ _1018;
  wire _1020 = _1016 ^ _1019;
  wire _1021 = uncoded_block[341] ^ uncoded_block[342];
  wire _1022 = _1021 ^ _159;
  wire _1023 = uncoded_block[347] ^ uncoded_block[348];
  wire _1024 = uncoded_block[351] ^ uncoded_block[352];
  wire _1025 = _1023 ^ _1024;
  wire _1026 = _1022 ^ _1025;
  wire _1027 = _1020 ^ _1026;
  wire _1028 = uncoded_block[353] ^ uncoded_block[354];
  wire _1029 = uncoded_block[357] ^ uncoded_block[359];
  wire _1030 = _1028 ^ _1029;
  wire _1031 = uncoded_block[361] ^ uncoded_block[363];
  wire _1032 = uncoded_block[364] ^ uncoded_block[367];
  wire _1033 = _1031 ^ _1032;
  wire _1034 = _1030 ^ _1033;
  wire _1035 = uncoded_block[370] ^ uncoded_block[372];
  wire _1036 = uncoded_block[374] ^ uncoded_block[375];
  wire _1037 = _1035 ^ _1036;
  wire _1038 = uncoded_block[381] ^ uncoded_block[382];
  wire _1039 = uncoded_block[384] ^ uncoded_block[385];
  wire _1040 = _1038 ^ _1039;
  wire _1041 = _1037 ^ _1040;
  wire _1042 = _1034 ^ _1041;
  wire _1043 = _1027 ^ _1042;
  wire _1044 = _1013 ^ _1043;
  wire _1045 = uncoded_block[387] ^ uncoded_block[391];
  wire _1046 = uncoded_block[392] ^ uncoded_block[397];
  wire _1047 = _1045 ^ _1046;
  wire _1048 = uncoded_block[398] ^ uncoded_block[399];
  wire _1049 = _1048 ^ _181;
  wire _1050 = _1047 ^ _1049;
  wire _1051 = uncoded_block[405] ^ uncoded_block[407];
  wire _1052 = uncoded_block[408] ^ uncoded_block[410];
  wire _1053 = _1051 ^ _1052;
  wire _1054 = uncoded_block[412] ^ uncoded_block[413];
  wire _1055 = uncoded_block[414] ^ uncoded_block[415];
  wire _1056 = _1054 ^ _1055;
  wire _1057 = _1053 ^ _1056;
  wire _1058 = _1050 ^ _1057;
  wire _1059 = uncoded_block[419] ^ uncoded_block[422];
  wire _1060 = uncoded_block[423] ^ uncoded_block[425];
  wire _1061 = _1059 ^ _1060;
  wire _1062 = uncoded_block[426] ^ uncoded_block[427];
  wire _1063 = uncoded_block[429] ^ uncoded_block[432];
  wire _1064 = _1062 ^ _1063;
  wire _1065 = _1061 ^ _1064;
  wire _1066 = uncoded_block[433] ^ uncoded_block[436];
  wire _1067 = uncoded_block[439] ^ uncoded_block[444];
  wire _1068 = _1066 ^ _1067;
  wire _1069 = uncoded_block[446] ^ uncoded_block[449];
  wire _1070 = uncoded_block[450] ^ uncoded_block[452];
  wire _1071 = _1069 ^ _1070;
  wire _1072 = _1068 ^ _1071;
  wire _1073 = _1065 ^ _1072;
  wire _1074 = _1058 ^ _1073;
  wire _1075 = uncoded_block[453] ^ uncoded_block[454];
  wire _1076 = uncoded_block[455] ^ uncoded_block[458];
  wire _1077 = _1075 ^ _1076;
  wire _1078 = uncoded_block[459] ^ uncoded_block[465];
  wire _1079 = uncoded_block[466] ^ uncoded_block[467];
  wire _1080 = _1078 ^ _1079;
  wire _1081 = _1077 ^ _1080;
  wire _1082 = uncoded_block[471] ^ uncoded_block[472];
  wire _1083 = uncoded_block[473] ^ uncoded_block[474];
  wire _1084 = _1082 ^ _1083;
  wire _1085 = uncoded_block[479] ^ uncoded_block[480];
  wire _1086 = uncoded_block[482] ^ uncoded_block[483];
  wire _1087 = _1085 ^ _1086;
  wire _1088 = _1084 ^ _1087;
  wire _1089 = _1081 ^ _1088;
  wire _1090 = uncoded_block[485] ^ uncoded_block[486];
  wire _1091 = uncoded_block[487] ^ uncoded_block[492];
  wire _1092 = _1090 ^ _1091;
  wire _1093 = uncoded_block[494] ^ uncoded_block[495];
  wire _1094 = uncoded_block[496] ^ uncoded_block[498];
  wire _1095 = _1093 ^ _1094;
  wire _1096 = _1092 ^ _1095;
  wire _1097 = uncoded_block[499] ^ uncoded_block[501];
  wire _1098 = _1097 ^ _229;
  wire _1099 = uncoded_block[508] ^ uncoded_block[515];
  wire _1100 = _1099 ^ _236;
  wire _1101 = _1098 ^ _1100;
  wire _1102 = _1096 ^ _1101;
  wire _1103 = _1089 ^ _1102;
  wire _1104 = _1074 ^ _1103;
  wire _1105 = _1044 ^ _1104;
  wire _1106 = _983 ^ _1105;
  wire _1107 = uncoded_block[520] ^ uncoded_block[521];
  wire _1108 = uncoded_block[522] ^ uncoded_block[523];
  wire _1109 = _1107 ^ _1108;
  wire _1110 = uncoded_block[524] ^ uncoded_block[527];
  wire _1111 = uncoded_block[530] ^ uncoded_block[531];
  wire _1112 = _1110 ^ _1111;
  wire _1113 = _1109 ^ _1112;
  wire _1114 = uncoded_block[533] ^ uncoded_block[535];
  wire _1115 = uncoded_block[537] ^ uncoded_block[540];
  wire _1116 = _1114 ^ _1115;
  wire _1117 = uncoded_block[544] ^ uncoded_block[545];
  wire _1118 = uncoded_block[547] ^ uncoded_block[550];
  wire _1119 = _1117 ^ _1118;
  wire _1120 = _1116 ^ _1119;
  wire _1121 = _1113 ^ _1120;
  wire _1122 = uncoded_block[554] ^ uncoded_block[555];
  wire _1123 = uncoded_block[556] ^ uncoded_block[557];
  wire _1124 = _1122 ^ _1123;
  wire _1125 = uncoded_block[558] ^ uncoded_block[564];
  wire _1126 = uncoded_block[565] ^ uncoded_block[566];
  wire _1127 = _1125 ^ _1126;
  wire _1128 = _1124 ^ _1127;
  wire _1129 = uncoded_block[567] ^ uncoded_block[570];
  wire _1130 = uncoded_block[572] ^ uncoded_block[575];
  wire _1131 = _1129 ^ _1130;
  wire _1132 = uncoded_block[576] ^ uncoded_block[577];
  wire _1133 = uncoded_block[578] ^ uncoded_block[579];
  wire _1134 = _1132 ^ _1133;
  wire _1135 = _1131 ^ _1134;
  wire _1136 = _1128 ^ _1135;
  wire _1137 = _1121 ^ _1136;
  wire _1138 = uncoded_block[580] ^ uncoded_block[582];
  wire _1139 = uncoded_block[585] ^ uncoded_block[586];
  wire _1140 = _1138 ^ _1139;
  wire _1141 = uncoded_block[589] ^ uncoded_block[590];
  wire _1142 = uncoded_block[598] ^ uncoded_block[600];
  wire _1143 = _1141 ^ _1142;
  wire _1144 = _1140 ^ _1143;
  wire _1145 = uncoded_block[601] ^ uncoded_block[604];
  wire _1146 = uncoded_block[605] ^ uncoded_block[607];
  wire _1147 = _1145 ^ _1146;
  wire _1148 = uncoded_block[610] ^ uncoded_block[614];
  wire _1149 = uncoded_block[615] ^ uncoded_block[616];
  wire _1150 = _1148 ^ _1149;
  wire _1151 = _1147 ^ _1150;
  wire _1152 = _1144 ^ _1151;
  wire _1153 = uncoded_block[617] ^ uncoded_block[624];
  wire _1154 = uncoded_block[626] ^ uncoded_block[627];
  wire _1155 = _1153 ^ _1154;
  wire _1156 = uncoded_block[628] ^ uncoded_block[630];
  wire _1157 = uncoded_block[632] ^ uncoded_block[635];
  wire _1158 = _1156 ^ _1157;
  wire _1159 = _1155 ^ _1158;
  wire _1160 = uncoded_block[636] ^ uncoded_block[637];
  wire _1161 = uncoded_block[638] ^ uncoded_block[639];
  wire _1162 = _1160 ^ _1161;
  wire _1163 = uncoded_block[640] ^ uncoded_block[641];
  wire _1164 = uncoded_block[645] ^ uncoded_block[647];
  wire _1165 = _1163 ^ _1164;
  wire _1166 = _1162 ^ _1165;
  wire _1167 = _1159 ^ _1166;
  wire _1168 = _1152 ^ _1167;
  wire _1169 = _1137 ^ _1168;
  wire _1170 = uncoded_block[650] ^ uncoded_block[654];
  wire _1171 = uncoded_block[655] ^ uncoded_block[664];
  wire _1172 = _1170 ^ _1171;
  wire _1173 = uncoded_block[665] ^ uncoded_block[666];
  wire _1174 = uncoded_block[668] ^ uncoded_block[669];
  wire _1175 = _1173 ^ _1174;
  wire _1176 = _1172 ^ _1175;
  wire _1177 = uncoded_block[670] ^ uncoded_block[671];
  wire _1178 = uncoded_block[672] ^ uncoded_block[673];
  wire _1179 = _1177 ^ _1178;
  wire _1180 = uncoded_block[675] ^ uncoded_block[677];
  wire _1181 = uncoded_block[679] ^ uncoded_block[681];
  wire _1182 = _1180 ^ _1181;
  wire _1183 = _1179 ^ _1182;
  wire _1184 = _1176 ^ _1183;
  wire _1185 = uncoded_block[683] ^ uncoded_block[687];
  wire _1186 = uncoded_block[690] ^ uncoded_block[693];
  wire _1187 = _1185 ^ _1186;
  wire _1188 = uncoded_block[697] ^ uncoded_block[703];
  wire _1189 = _328 ^ _1188;
  wire _1190 = _1187 ^ _1189;
  wire _1191 = uncoded_block[705] ^ uncoded_block[708];
  wire _1192 = uncoded_block[710] ^ uncoded_block[711];
  wire _1193 = _1191 ^ _1192;
  wire _1194 = uncoded_block[714] ^ uncoded_block[715];
  wire _1195 = uncoded_block[716] ^ uncoded_block[717];
  wire _1196 = _1194 ^ _1195;
  wire _1197 = _1193 ^ _1196;
  wire _1198 = _1190 ^ _1197;
  wire _1199 = _1184 ^ _1198;
  wire _1200 = uncoded_block[718] ^ uncoded_block[722];
  wire _1201 = _1200 ^ _344;
  wire _1202 = uncoded_block[729] ^ uncoded_block[733];
  wire _1203 = uncoded_block[734] ^ uncoded_block[735];
  wire _1204 = _1202 ^ _1203;
  wire _1205 = _1201 ^ _1204;
  wire _1206 = uncoded_block[736] ^ uncoded_block[737];
  wire _1207 = uncoded_block[740] ^ uncoded_block[742];
  wire _1208 = _1206 ^ _1207;
  wire _1209 = uncoded_block[744] ^ uncoded_block[747];
  wire _1210 = uncoded_block[749] ^ uncoded_block[750];
  wire _1211 = _1209 ^ _1210;
  wire _1212 = _1208 ^ _1211;
  wire _1213 = _1205 ^ _1212;
  wire _1214 = uncoded_block[752] ^ uncoded_block[753];
  wire _1215 = uncoded_block[755] ^ uncoded_block[758];
  wire _1216 = _1214 ^ _1215;
  wire _1217 = uncoded_block[763] ^ uncoded_block[764];
  wire _1218 = uncoded_block[769] ^ uncoded_block[770];
  wire _1219 = _1217 ^ _1218;
  wire _1220 = _1216 ^ _1219;
  wire _1221 = uncoded_block[772] ^ uncoded_block[773];
  wire _1222 = uncoded_block[774] ^ uncoded_block[781];
  wire _1223 = _1221 ^ _1222;
  wire _1224 = uncoded_block[786] ^ uncoded_block[787];
  wire _1225 = uncoded_block[789] ^ uncoded_block[791];
  wire _1226 = _1224 ^ _1225;
  wire _1227 = _1223 ^ _1226;
  wire _1228 = _1220 ^ _1227;
  wire _1229 = _1213 ^ _1228;
  wire _1230 = _1199 ^ _1229;
  wire _1231 = _1169 ^ _1230;
  wire _1232 = uncoded_block[792] ^ uncoded_block[794];
  wire _1233 = uncoded_block[795] ^ uncoded_block[797];
  wire _1234 = _1232 ^ _1233;
  wire _1235 = uncoded_block[803] ^ uncoded_block[805];
  wire _1236 = _383 ^ _1235;
  wire _1237 = _1234 ^ _1236;
  wire _1238 = uncoded_block[807] ^ uncoded_block[808];
  wire _1239 = uncoded_block[813] ^ uncoded_block[816];
  wire _1240 = _1238 ^ _1239;
  wire _1241 = uncoded_block[817] ^ uncoded_block[818];
  wire _1242 = uncoded_block[819] ^ uncoded_block[820];
  wire _1243 = _1241 ^ _1242;
  wire _1244 = _1240 ^ _1243;
  wire _1245 = _1237 ^ _1244;
  wire _1246 = uncoded_block[824] ^ uncoded_block[825];
  wire _1247 = uncoded_block[826] ^ uncoded_block[828];
  wire _1248 = _1246 ^ _1247;
  wire _1249 = uncoded_block[829] ^ uncoded_block[831];
  wire _1250 = uncoded_block[833] ^ uncoded_block[834];
  wire _1251 = _1249 ^ _1250;
  wire _1252 = _1248 ^ _1251;
  wire _1253 = uncoded_block[835] ^ uncoded_block[837];
  wire _1254 = uncoded_block[839] ^ uncoded_block[841];
  wire _1255 = _1253 ^ _1254;
  wire _1256 = uncoded_block[843] ^ uncoded_block[844];
  wire _1257 = uncoded_block[846] ^ uncoded_block[847];
  wire _1258 = _1256 ^ _1257;
  wire _1259 = _1255 ^ _1258;
  wire _1260 = _1252 ^ _1259;
  wire _1261 = _1245 ^ _1260;
  wire _1262 = uncoded_block[850] ^ uncoded_block[854];
  wire _1263 = uncoded_block[855] ^ uncoded_block[860];
  wire _1264 = _1262 ^ _1263;
  wire _1265 = uncoded_block[862] ^ uncoded_block[866];
  wire _1266 = uncoded_block[867] ^ uncoded_block[868];
  wire _1267 = _1265 ^ _1266;
  wire _1268 = _1264 ^ _1267;
  wire _1269 = uncoded_block[872] ^ uncoded_block[873];
  wire _1270 = uncoded_block[876] ^ uncoded_block[883];
  wire _1271 = _1269 ^ _1270;
  wire _1272 = uncoded_block[884] ^ uncoded_block[887];
  wire _1273 = uncoded_block[888] ^ uncoded_block[890];
  wire _1274 = _1272 ^ _1273;
  wire _1275 = _1271 ^ _1274;
  wire _1276 = _1268 ^ _1275;
  wire _1277 = uncoded_block[893] ^ uncoded_block[895];
  wire _1278 = uncoded_block[898] ^ uncoded_block[899];
  wire _1279 = _1277 ^ _1278;
  wire _1280 = uncoded_block[902] ^ uncoded_block[904];
  wire _1281 = uncoded_block[905] ^ uncoded_block[906];
  wire _1282 = _1280 ^ _1281;
  wire _1283 = _1279 ^ _1282;
  wire _1284 = uncoded_block[907] ^ uncoded_block[908];
  wire _1285 = uncoded_block[909] ^ uncoded_block[911];
  wire _1286 = _1284 ^ _1285;
  wire _1287 = uncoded_block[913] ^ uncoded_block[914];
  wire _1288 = uncoded_block[915] ^ uncoded_block[919];
  wire _1289 = _1287 ^ _1288;
  wire _1290 = _1286 ^ _1289;
  wire _1291 = _1283 ^ _1290;
  wire _1292 = _1276 ^ _1291;
  wire _1293 = _1261 ^ _1292;
  wire _1294 = _439 ^ _445;
  wire _1295 = uncoded_block[925] ^ uncoded_block[926];
  wire _1296 = uncoded_block[929] ^ uncoded_block[930];
  wire _1297 = _1295 ^ _1296;
  wire _1298 = _1294 ^ _1297;
  wire _1299 = uncoded_block[933] ^ uncoded_block[936];
  wire _1300 = uncoded_block[940] ^ uncoded_block[944];
  wire _1301 = _1299 ^ _1300;
  wire _1302 = uncoded_block[945] ^ uncoded_block[947];
  wire _1303 = uncoded_block[951] ^ uncoded_block[952];
  wire _1304 = _1302 ^ _1303;
  wire _1305 = _1301 ^ _1304;
  wire _1306 = _1298 ^ _1305;
  wire _1307 = uncoded_block[956] ^ uncoded_block[957];
  wire _1308 = uncoded_block[959] ^ uncoded_block[960];
  wire _1309 = _1307 ^ _1308;
  wire _1310 = uncoded_block[962] ^ uncoded_block[963];
  wire _1311 = uncoded_block[965] ^ uncoded_block[969];
  wire _1312 = _1310 ^ _1311;
  wire _1313 = _1309 ^ _1312;
  wire _1314 = uncoded_block[970] ^ uncoded_block[971];
  wire _1315 = uncoded_block[972] ^ uncoded_block[974];
  wire _1316 = _1314 ^ _1315;
  wire _1317 = uncoded_block[986] ^ uncoded_block[987];
  wire _1318 = uncoded_block[988] ^ uncoded_block[990];
  wire _1319 = _1317 ^ _1318;
  wire _1320 = _1316 ^ _1319;
  wire _1321 = _1313 ^ _1320;
  wire _1322 = _1306 ^ _1321;
  wire _1323 = uncoded_block[991] ^ uncoded_block[992];
  wire _1324 = uncoded_block[993] ^ uncoded_block[1000];
  wire _1325 = _1323 ^ _1324;
  wire _1326 = uncoded_block[1002] ^ uncoded_block[1006];
  wire _1327 = uncoded_block[1007] ^ uncoded_block[1009];
  wire _1328 = _1326 ^ _1327;
  wire _1329 = _1325 ^ _1328;
  wire _1330 = uncoded_block[1010] ^ uncoded_block[1012];
  wire _1331 = uncoded_block[1014] ^ uncoded_block[1015];
  wire _1332 = _1330 ^ _1331;
  wire _1333 = uncoded_block[1017] ^ uncoded_block[1020];
  wire _1334 = uncoded_block[1021] ^ uncoded_block[1022];
  wire _1335 = _1333 ^ _1334;
  wire _1336 = _1332 ^ _1335;
  wire _1337 = _1329 ^ _1336;
  wire _1338 = uncoded_block[1023] ^ uncoded_block[1024];
  wire _1339 = uncoded_block[1027] ^ uncoded_block[1029];
  wire _1340 = _1338 ^ _1339;
  wire _1341 = uncoded_block[1030] ^ uncoded_block[1034];
  wire _1342 = uncoded_block[1035] ^ uncoded_block[1036];
  wire _1343 = _1341 ^ _1342;
  wire _1344 = _1340 ^ _1343;
  wire _1345 = uncoded_block[1038] ^ uncoded_block[1039];
  wire _1346 = uncoded_block[1040] ^ uncoded_block[1041];
  wire _1347 = _1345 ^ _1346;
  wire _1348 = _512 ^ _514;
  wire _1349 = _1347 ^ _1348;
  wire _1350 = _1344 ^ _1349;
  wire _1351 = _1337 ^ _1350;
  wire _1352 = _1322 ^ _1351;
  wire _1353 = _1293 ^ _1352;
  wire _1354 = _1231 ^ _1353;
  wire _1355 = _1106 ^ _1354;
  wire _1356 = uncoded_block[1046] ^ uncoded_block[1047];
  wire _1357 = uncoded_block[1049] ^ uncoded_block[1050];
  wire _1358 = _1356 ^ _1357;
  wire _1359 = uncoded_block[1053] ^ uncoded_block[1054];
  wire _1360 = uncoded_block[1055] ^ uncoded_block[1057];
  wire _1361 = _1359 ^ _1360;
  wire _1362 = _1358 ^ _1361;
  wire _1363 = uncoded_block[1058] ^ uncoded_block[1059];
  wire _1364 = uncoded_block[1061] ^ uncoded_block[1065];
  wire _1365 = _1363 ^ _1364;
  wire _1366 = uncoded_block[1069] ^ uncoded_block[1070];
  wire _1367 = _1366 ^ _529;
  wire _1368 = _1365 ^ _1367;
  wire _1369 = _1362 ^ _1368;
  wire _1370 = uncoded_block[1078] ^ uncoded_block[1081];
  wire _1371 = uncoded_block[1082] ^ uncoded_block[1084];
  wire _1372 = _1370 ^ _1371;
  wire _1373 = uncoded_block[1085] ^ uncoded_block[1087];
  wire _1374 = uncoded_block[1088] ^ uncoded_block[1089];
  wire _1375 = _1373 ^ _1374;
  wire _1376 = _1372 ^ _1375;
  wire _1377 = uncoded_block[1092] ^ uncoded_block[1093];
  wire _1378 = uncoded_block[1094] ^ uncoded_block[1096];
  wire _1379 = _1377 ^ _1378;
  wire _1380 = uncoded_block[1097] ^ uncoded_block[1099];
  wire _1381 = _1380 ^ _546;
  wire _1382 = _1379 ^ _1381;
  wire _1383 = _1376 ^ _1382;
  wire _1384 = _1369 ^ _1383;
  wire _1385 = uncoded_block[1108] ^ uncoded_block[1111];
  wire _1386 = uncoded_block[1112] ^ uncoded_block[1114];
  wire _1387 = _1385 ^ _1386;
  wire _1388 = uncoded_block[1117] ^ uncoded_block[1118];
  wire _1389 = uncoded_block[1120] ^ uncoded_block[1123];
  wire _1390 = _1388 ^ _1389;
  wire _1391 = _1387 ^ _1390;
  wire _1392 = uncoded_block[1124] ^ uncoded_block[1128];
  wire _1393 = uncoded_block[1131] ^ uncoded_block[1132];
  wire _1394 = _1392 ^ _1393;
  wire _1395 = uncoded_block[1133] ^ uncoded_block[1137];
  wire _1396 = uncoded_block[1138] ^ uncoded_block[1141];
  wire _1397 = _1395 ^ _1396;
  wire _1398 = _1394 ^ _1397;
  wire _1399 = _1391 ^ _1398;
  wire _1400 = uncoded_block[1142] ^ uncoded_block[1145];
  wire _1401 = uncoded_block[1147] ^ uncoded_block[1149];
  wire _1402 = _1400 ^ _1401;
  wire _1403 = uncoded_block[1151] ^ uncoded_block[1157];
  wire _1404 = uncoded_block[1159] ^ uncoded_block[1160];
  wire _1405 = _1403 ^ _1404;
  wire _1406 = _1402 ^ _1405;
  wire _1407 = uncoded_block[1163] ^ uncoded_block[1165];
  wire _1408 = uncoded_block[1169] ^ uncoded_block[1170];
  wire _1409 = _1407 ^ _1408;
  wire _1410 = uncoded_block[1172] ^ uncoded_block[1173];
  wire _1411 = uncoded_block[1176] ^ uncoded_block[1179];
  wire _1412 = _1410 ^ _1411;
  wire _1413 = _1409 ^ _1412;
  wire _1414 = _1406 ^ _1413;
  wire _1415 = _1399 ^ _1414;
  wire _1416 = _1384 ^ _1415;
  wire _1417 = uncoded_block[1181] ^ uncoded_block[1183];
  wire _1418 = uncoded_block[1185] ^ uncoded_block[1188];
  wire _1419 = _1417 ^ _1418;
  wire _1420 = uncoded_block[1192] ^ uncoded_block[1193];
  wire _1421 = uncoded_block[1196] ^ uncoded_block[1197];
  wire _1422 = _1420 ^ _1421;
  wire _1423 = _1419 ^ _1422;
  wire _1424 = uncoded_block[1199] ^ uncoded_block[1203];
  wire _1425 = uncoded_block[1204] ^ uncoded_block[1206];
  wire _1426 = _1424 ^ _1425;
  wire _1427 = uncoded_block[1210] ^ uncoded_block[1211];
  wire _1428 = uncoded_block[1212] ^ uncoded_block[1213];
  wire _1429 = _1427 ^ _1428;
  wire _1430 = _1426 ^ _1429;
  wire _1431 = _1423 ^ _1430;
  wire _1432 = uncoded_block[1215] ^ uncoded_block[1218];
  wire _1433 = uncoded_block[1220] ^ uncoded_block[1223];
  wire _1434 = _1432 ^ _1433;
  wire _1435 = uncoded_block[1224] ^ uncoded_block[1225];
  wire _1436 = uncoded_block[1227] ^ uncoded_block[1228];
  wire _1437 = _1435 ^ _1436;
  wire _1438 = _1434 ^ _1437;
  wire _1439 = uncoded_block[1229] ^ uncoded_block[1230];
  wire _1440 = uncoded_block[1231] ^ uncoded_block[1233];
  wire _1441 = _1439 ^ _1440;
  wire _1442 = uncoded_block[1234] ^ uncoded_block[1235];
  wire _1443 = uncoded_block[1236] ^ uncoded_block[1239];
  wire _1444 = _1442 ^ _1443;
  wire _1445 = _1441 ^ _1444;
  wire _1446 = _1438 ^ _1445;
  wire _1447 = _1431 ^ _1446;
  wire _1448 = uncoded_block[1242] ^ uncoded_block[1244];
  wire _1449 = uncoded_block[1246] ^ uncoded_block[1247];
  wire _1450 = _1448 ^ _1449;
  wire _1451 = uncoded_block[1248] ^ uncoded_block[1249];
  wire _1452 = uncoded_block[1251] ^ uncoded_block[1255];
  wire _1453 = _1451 ^ _1452;
  wire _1454 = _1450 ^ _1453;
  wire _1455 = uncoded_block[1256] ^ uncoded_block[1257];
  wire _1456 = uncoded_block[1258] ^ uncoded_block[1261];
  wire _1457 = _1455 ^ _1456;
  wire _1458 = uncoded_block[1264] ^ uncoded_block[1266];
  wire _1459 = uncoded_block[1269] ^ uncoded_block[1270];
  wire _1460 = _1458 ^ _1459;
  wire _1461 = _1457 ^ _1460;
  wire _1462 = _1454 ^ _1461;
  wire _1463 = uncoded_block[1275] ^ uncoded_block[1276];
  wire _1464 = _628 ^ _1463;
  wire _1465 = uncoded_block[1277] ^ uncoded_block[1285];
  wire _1466 = _1465 ^ _639;
  wire _1467 = _1464 ^ _1466;
  wire _1468 = uncoded_block[1290] ^ uncoded_block[1291];
  wire _1469 = uncoded_block[1292] ^ uncoded_block[1293];
  wire _1470 = _1468 ^ _1469;
  wire _1471 = uncoded_block[1296] ^ uncoded_block[1301];
  wire _1472 = uncoded_block[1302] ^ uncoded_block[1304];
  wire _1473 = _1471 ^ _1472;
  wire _1474 = _1470 ^ _1473;
  wire _1475 = _1467 ^ _1474;
  wire _1476 = _1462 ^ _1475;
  wire _1477 = _1447 ^ _1476;
  wire _1478 = _1416 ^ _1477;
  wire _1479 = uncoded_block[1305] ^ uncoded_block[1307];
  wire _1480 = uncoded_block[1309] ^ uncoded_block[1310];
  wire _1481 = _1479 ^ _1480;
  wire _1482 = uncoded_block[1311] ^ uncoded_block[1312];
  wire _1483 = uncoded_block[1313] ^ uncoded_block[1315];
  wire _1484 = _1482 ^ _1483;
  wire _1485 = _1481 ^ _1484;
  wire _1486 = uncoded_block[1317] ^ uncoded_block[1320];
  wire _1487 = uncoded_block[1321] ^ uncoded_block[1323];
  wire _1488 = _1486 ^ _1487;
  wire _1489 = uncoded_block[1326] ^ uncoded_block[1327];
  wire _1490 = uncoded_block[1328] ^ uncoded_block[1329];
  wire _1491 = _1489 ^ _1490;
  wire _1492 = _1488 ^ _1491;
  wire _1493 = _1485 ^ _1492;
  wire _1494 = uncoded_block[1330] ^ uncoded_block[1331];
  wire _1495 = uncoded_block[1334] ^ uncoded_block[1338];
  wire _1496 = _1494 ^ _1495;
  wire _1497 = uncoded_block[1340] ^ uncoded_block[1341];
  wire _1498 = uncoded_block[1344] ^ uncoded_block[1345];
  wire _1499 = _1497 ^ _1498;
  wire _1500 = _1496 ^ _1499;
  wire _1501 = uncoded_block[1346] ^ uncoded_block[1348];
  wire _1502 = uncoded_block[1352] ^ uncoded_block[1355];
  wire _1503 = _1501 ^ _1502;
  wire _1504 = uncoded_block[1362] ^ uncoded_block[1363];
  wire _1505 = _1504 ^ _679;
  wire _1506 = _1503 ^ _1505;
  wire _1507 = _1500 ^ _1506;
  wire _1508 = _1493 ^ _1507;
  wire _1509 = uncoded_block[1369] ^ uncoded_block[1372];
  wire _1510 = uncoded_block[1374] ^ uncoded_block[1382];
  wire _1511 = _1509 ^ _1510;
  wire _1512 = uncoded_block[1385] ^ uncoded_block[1388];
  wire _1513 = uncoded_block[1389] ^ uncoded_block[1390];
  wire _1514 = _1512 ^ _1513;
  wire _1515 = _1511 ^ _1514;
  wire _1516 = uncoded_block[1396] ^ uncoded_block[1398];
  wire _1517 = uncoded_block[1399] ^ uncoded_block[1401];
  wire _1518 = _1516 ^ _1517;
  wire _1519 = uncoded_block[1402] ^ uncoded_block[1404];
  wire _1520 = _1519 ^ _701;
  wire _1521 = _1518 ^ _1520;
  wire _1522 = _1515 ^ _1521;
  wire _1523 = uncoded_block[1409] ^ uncoded_block[1412];
  wire _1524 = uncoded_block[1413] ^ uncoded_block[1417];
  wire _1525 = _1523 ^ _1524;
  wire _1526 = uncoded_block[1420] ^ uncoded_block[1422];
  wire _1527 = uncoded_block[1423] ^ uncoded_block[1425];
  wire _1528 = _1526 ^ _1527;
  wire _1529 = _1525 ^ _1528;
  wire _1530 = uncoded_block[1427] ^ uncoded_block[1429];
  wire _1531 = uncoded_block[1430] ^ uncoded_block[1431];
  wire _1532 = _1530 ^ _1531;
  wire _1533 = uncoded_block[1432] ^ uncoded_block[1433];
  wire _1534 = uncoded_block[1434] ^ uncoded_block[1435];
  wire _1535 = _1533 ^ _1534;
  wire _1536 = _1532 ^ _1535;
  wire _1537 = _1529 ^ _1536;
  wire _1538 = _1522 ^ _1537;
  wire _1539 = _1508 ^ _1538;
  wire _1540 = uncoded_block[1436] ^ uncoded_block[1439];
  wire _1541 = uncoded_block[1442] ^ uncoded_block[1444];
  wire _1542 = _1540 ^ _1541;
  wire _1543 = uncoded_block[1448] ^ uncoded_block[1451];
  wire _1544 = uncoded_block[1452] ^ uncoded_block[1454];
  wire _1545 = _1543 ^ _1544;
  wire _1546 = _1542 ^ _1545;
  wire _1547 = uncoded_block[1456] ^ uncoded_block[1464];
  wire _1548 = uncoded_block[1465] ^ uncoded_block[1466];
  wire _1549 = _1547 ^ _1548;
  wire _1550 = uncoded_block[1467] ^ uncoded_block[1468];
  wire _1551 = uncoded_block[1470] ^ uncoded_block[1472];
  wire _1552 = _1550 ^ _1551;
  wire _1553 = _1549 ^ _1552;
  wire _1554 = _1546 ^ _1553;
  wire _1555 = uncoded_block[1475] ^ uncoded_block[1477];
  wire _1556 = uncoded_block[1478] ^ uncoded_block[1479];
  wire _1557 = _1555 ^ _1556;
  wire _1558 = uncoded_block[1480] ^ uncoded_block[1481];
  wire _1559 = uncoded_block[1482] ^ uncoded_block[1483];
  wire _1560 = _1558 ^ _1559;
  wire _1561 = _1557 ^ _1560;
  wire _1562 = uncoded_block[1485] ^ uncoded_block[1487];
  wire _1563 = uncoded_block[1489] ^ uncoded_block[1490];
  wire _1564 = _1562 ^ _1563;
  wire _1565 = uncoded_block[1492] ^ uncoded_block[1493];
  wire _1566 = uncoded_block[1494] ^ uncoded_block[1498];
  wire _1567 = _1565 ^ _1566;
  wire _1568 = _1564 ^ _1567;
  wire _1569 = _1561 ^ _1568;
  wire _1570 = _1554 ^ _1569;
  wire _1571 = uncoded_block[1500] ^ uncoded_block[1501];
  wire _1572 = uncoded_block[1503] ^ uncoded_block[1504];
  wire _1573 = _1571 ^ _1572;
  wire _1574 = uncoded_block[1506] ^ uncoded_block[1509];
  wire _1575 = uncoded_block[1511] ^ uncoded_block[1513];
  wire _1576 = _1574 ^ _1575;
  wire _1577 = _1573 ^ _1576;
  wire _1578 = uncoded_block[1514] ^ uncoded_block[1518];
  wire _1579 = uncoded_block[1520] ^ uncoded_block[1522];
  wire _1580 = _1578 ^ _1579;
  wire _1581 = uncoded_block[1524] ^ uncoded_block[1526];
  wire _1582 = uncoded_block[1528] ^ uncoded_block[1529];
  wire _1583 = _1581 ^ _1582;
  wire _1584 = _1580 ^ _1583;
  wire _1585 = _1577 ^ _1584;
  wire _1586 = uncoded_block[1534] ^ uncoded_block[1536];
  wire _1587 = uncoded_block[1537] ^ uncoded_block[1539];
  wire _1588 = _1586 ^ _1587;
  wire _1589 = uncoded_block[1541] ^ uncoded_block[1542];
  wire _1590 = uncoded_block[1543] ^ uncoded_block[1544];
  wire _1591 = _1589 ^ _1590;
  wire _1592 = _1588 ^ _1591;
  wire _1593 = uncoded_block[1545] ^ uncoded_block[1547];
  wire _1594 = uncoded_block[1548] ^ uncoded_block[1554];
  wire _1595 = _1593 ^ _1594;
  wire _1596 = uncoded_block[1556] ^ uncoded_block[1557];
  wire _1597 = uncoded_block[1559] ^ uncoded_block[1560];
  wire _1598 = _1596 ^ _1597;
  wire _1599 = _1595 ^ _1598;
  wire _1600 = _1592 ^ _1599;
  wire _1601 = _1585 ^ _1600;
  wire _1602 = _1570 ^ _1601;
  wire _1603 = _1539 ^ _1602;
  wire _1604 = _1478 ^ _1603;
  wire _1605 = uncoded_block[1563] ^ uncoded_block[1566];
  wire _1606 = uncoded_block[1567] ^ uncoded_block[1568];
  wire _1607 = _1605 ^ _1606;
  wire _1608 = uncoded_block[1574] ^ uncoded_block[1576];
  wire _1609 = uncoded_block[1579] ^ uncoded_block[1581];
  wire _1610 = _1608 ^ _1609;
  wire _1611 = _1607 ^ _1610;
  wire _1612 = uncoded_block[1582] ^ uncoded_block[1583];
  wire _1613 = uncoded_block[1584] ^ uncoded_block[1585];
  wire _1614 = _1612 ^ _1613;
  wire _1615 = uncoded_block[1586] ^ uncoded_block[1587];
  wire _1616 = uncoded_block[1588] ^ uncoded_block[1591];
  wire _1617 = _1615 ^ _1616;
  wire _1618 = _1614 ^ _1617;
  wire _1619 = _1611 ^ _1618;
  wire _1620 = uncoded_block[1597] ^ uncoded_block[1598];
  wire _1621 = uncoded_block[1599] ^ uncoded_block[1600];
  wire _1622 = _1620 ^ _1621;
  wire _1623 = _793 ^ _1622;
  wire _1624 = uncoded_block[1601] ^ uncoded_block[1604];
  wire _1625 = uncoded_block[1605] ^ uncoded_block[1606];
  wire _1626 = _1624 ^ _1625;
  wire _1627 = uncoded_block[1607] ^ uncoded_block[1609];
  wire _1628 = _1627 ^ _801;
  wire _1629 = _1626 ^ _1628;
  wire _1630 = _1623 ^ _1629;
  wire _1631 = _1619 ^ _1630;
  wire _1632 = uncoded_block[1613] ^ uncoded_block[1615];
  wire _1633 = uncoded_block[1616] ^ uncoded_block[1619];
  wire _1634 = _1632 ^ _1633;
  wire _1635 = uncoded_block[1620] ^ uncoded_block[1626];
  wire _1636 = uncoded_block[1628] ^ uncoded_block[1629];
  wire _1637 = _1635 ^ _1636;
  wire _1638 = _1634 ^ _1637;
  wire _1639 = uncoded_block[1630] ^ uncoded_block[1631];
  wire _1640 = _1639 ^ _812;
  wire _1641 = uncoded_block[1634] ^ uncoded_block[1635];
  wire _1642 = uncoded_block[1637] ^ uncoded_block[1638];
  wire _1643 = _1641 ^ _1642;
  wire _1644 = _1640 ^ _1643;
  wire _1645 = _1638 ^ _1644;
  wire _1646 = uncoded_block[1640] ^ uncoded_block[1643];
  wire _1647 = uncoded_block[1644] ^ uncoded_block[1646];
  wire _1648 = _1646 ^ _1647;
  wire _1649 = uncoded_block[1648] ^ uncoded_block[1649];
  wire _1650 = uncoded_block[1650] ^ uncoded_block[1654];
  wire _1651 = _1649 ^ _1650;
  wire _1652 = _1648 ^ _1651;
  wire _1653 = uncoded_block[1658] ^ uncoded_block[1659];
  wire _1654 = uncoded_block[1663] ^ uncoded_block[1664];
  wire _1655 = _1653 ^ _1654;
  wire _1656 = uncoded_block[1668] ^ uncoded_block[1673];
  wire _1657 = _1656 ^ _830;
  wire _1658 = _1655 ^ _1657;
  wire _1659 = _1652 ^ _1658;
  wire _1660 = _1645 ^ _1659;
  wire _1661 = _1631 ^ _1660;
  wire _1662 = uncoded_block[1676] ^ uncoded_block[1679];
  wire _1663 = uncoded_block[1680] ^ uncoded_block[1683];
  wire _1664 = _1662 ^ _1663;
  wire _1665 = uncoded_block[1686] ^ uncoded_block[1688];
  wire _1666 = uncoded_block[1690] ^ uncoded_block[1694];
  wire _1667 = _1665 ^ _1666;
  wire _1668 = _1664 ^ _1667;
  wire _1669 = uncoded_block[1696] ^ uncoded_block[1698];
  wire _1670 = uncoded_block[1699] ^ uncoded_block[1704];
  wire _1671 = _1669 ^ _1670;
  wire _1672 = uncoded_block[1705] ^ uncoded_block[1707];
  wire _1673 = uncoded_block[1710] ^ uncoded_block[1715];
  wire _1674 = _1672 ^ _1673;
  wire _1675 = _1671 ^ _1674;
  wire _1676 = _1668 ^ _1675;
  wire _1677 = uncoded_block[1716] ^ uncoded_block[1717];
  wire _1678 = _1677 ^ uncoded_block[1721];
  wire _1679 = _1676 ^ _1678;
  wire _1680 = _1661 ^ _1679;
  wire _1681 = _1604 ^ _1680;
  wire _1682 = _1355 ^ _1681;
  wire _1683 = uncoded_block[2] ^ uncoded_block[4];
  wire _1684 = uncoded_block[7] ^ uncoded_block[10];
  wire _1685 = _1683 ^ _1684;
  wire _1686 = uncoded_block[11] ^ uncoded_block[13];
  wire _1687 = uncoded_block[15] ^ uncoded_block[18];
  wire _1688 = _1686 ^ _1687;
  wire _1689 = _1685 ^ _1688;
  wire _1690 = uncoded_block[20] ^ uncoded_block[21];
  wire _1691 = uncoded_block[22] ^ uncoded_block[26];
  wire _1692 = _1690 ^ _1691;
  wire _1693 = uncoded_block[28] ^ uncoded_block[31];
  wire _1694 = _1693 ^ _15;
  wire _1695 = _1692 ^ _1694;
  wire _1696 = _1689 ^ _1695;
  wire _1697 = uncoded_block[38] ^ uncoded_block[42];
  wire _1698 = _16 ^ _1697;
  wire _1699 = uncoded_block[49] ^ uncoded_block[50];
  wire _1700 = uncoded_block[53] ^ uncoded_block[54];
  wire _1701 = _1699 ^ _1700;
  wire _1702 = _1698 ^ _1701;
  wire _1703 = uncoded_block[56] ^ uncoded_block[57];
  wire _1704 = _1703 ^ _889;
  wire _1705 = uncoded_block[61] ^ uncoded_block[64];
  wire _1706 = uncoded_block[65] ^ uncoded_block[67];
  wire _1707 = _1705 ^ _1706;
  wire _1708 = _1704 ^ _1707;
  wire _1709 = _1702 ^ _1708;
  wire _1710 = _1696 ^ _1709;
  wire _1711 = uncoded_block[71] ^ uncoded_block[72];
  wire _1712 = uncoded_block[75] ^ uncoded_block[76];
  wire _1713 = _1711 ^ _1712;
  wire _1714 = uncoded_block[77] ^ uncoded_block[79];
  wire _1715 = uncoded_block[81] ^ uncoded_block[90];
  wire _1716 = _1714 ^ _1715;
  wire _1717 = _1713 ^ _1716;
  wire _1718 = uncoded_block[91] ^ uncoded_block[93];
  wire _1719 = uncoded_block[95] ^ uncoded_block[99];
  wire _1720 = _1718 ^ _1719;
  wire _1721 = uncoded_block[103] ^ uncoded_block[105];
  wire _1722 = uncoded_block[107] ^ uncoded_block[108];
  wire _1723 = _1721 ^ _1722;
  wire _1724 = _1720 ^ _1723;
  wire _1725 = _1717 ^ _1724;
  wire _1726 = uncoded_block[110] ^ uncoded_block[112];
  wire _1727 = uncoded_block[115] ^ uncoded_block[118];
  wire _1728 = _1726 ^ _1727;
  wire _1729 = uncoded_block[119] ^ uncoded_block[121];
  wire _1730 = uncoded_block[125] ^ uncoded_block[126];
  wire _1731 = _1729 ^ _1730;
  wire _1732 = _1728 ^ _1731;
  wire _1733 = uncoded_block[127] ^ uncoded_block[128];
  wire _1734 = _1733 ^ _923;
  wire _1735 = uncoded_block[131] ^ uncoded_block[132];
  wire _1736 = uncoded_block[136] ^ uncoded_block[137];
  wire _1737 = _1735 ^ _1736;
  wire _1738 = _1734 ^ _1737;
  wire _1739 = _1732 ^ _1738;
  wire _1740 = _1725 ^ _1739;
  wire _1741 = _1710 ^ _1740;
  wire _1742 = uncoded_block[145] ^ uncoded_block[146];
  wire _1743 = _64 ^ _1742;
  wire _1744 = uncoded_block[149] ^ uncoded_block[150];
  wire _1745 = uncoded_block[151] ^ uncoded_block[152];
  wire _1746 = _1744 ^ _1745;
  wire _1747 = _1743 ^ _1746;
  wire _1748 = uncoded_block[156] ^ uncoded_block[157];
  wire _1749 = uncoded_block[163] ^ uncoded_block[164];
  wire _1750 = _1748 ^ _1749;
  wire _1751 = uncoded_block[166] ^ uncoded_block[167];
  wire _1752 = uncoded_block[169] ^ uncoded_block[171];
  wire _1753 = _1751 ^ _1752;
  wire _1754 = _1750 ^ _1753;
  wire _1755 = _1747 ^ _1754;
  wire _1756 = uncoded_block[174] ^ uncoded_block[176];
  wire _1757 = uncoded_block[179] ^ uncoded_block[182];
  wire _1758 = _1756 ^ _1757;
  wire _1759 = uncoded_block[185] ^ uncoded_block[186];
  wire _1760 = uncoded_block[187] ^ uncoded_block[192];
  wire _1761 = _1759 ^ _1760;
  wire _1762 = _1758 ^ _1761;
  wire _1763 = uncoded_block[193] ^ uncoded_block[195];
  wire _1764 = uncoded_block[205] ^ uncoded_block[206];
  wire _1765 = _1763 ^ _1764;
  wire _1766 = uncoded_block[208] ^ uncoded_block[211];
  wire _1767 = uncoded_block[213] ^ uncoded_block[215];
  wire _1768 = _1766 ^ _1767;
  wire _1769 = _1765 ^ _1768;
  wire _1770 = _1762 ^ _1769;
  wire _1771 = _1755 ^ _1770;
  wire _1772 = uncoded_block[217] ^ uncoded_block[219];
  wire _1773 = _1772 ^ _105;
  wire _1774 = uncoded_block[229] ^ uncoded_block[230];
  wire _1775 = uncoded_block[231] ^ uncoded_block[232];
  wire _1776 = _1774 ^ _1775;
  wire _1777 = _1773 ^ _1776;
  wire _1778 = uncoded_block[236] ^ uncoded_block[239];
  wire _1779 = _968 ^ _1778;
  wire _1780 = uncoded_block[240] ^ uncoded_block[242];
  wire _1781 = uncoded_block[245] ^ uncoded_block[247];
  wire _1782 = _1780 ^ _1781;
  wire _1783 = _1779 ^ _1782;
  wire _1784 = _1777 ^ _1783;
  wire _1785 = uncoded_block[251] ^ uncoded_block[254];
  wire _1786 = uncoded_block[256] ^ uncoded_block[257];
  wire _1787 = _1785 ^ _1786;
  wire _1788 = uncoded_block[258] ^ uncoded_block[260];
  wire _1789 = uncoded_block[261] ^ uncoded_block[265];
  wire _1790 = _1788 ^ _1789;
  wire _1791 = _1787 ^ _1790;
  wire _1792 = uncoded_block[266] ^ uncoded_block[269];
  wire _1793 = uncoded_block[270] ^ uncoded_block[273];
  wire _1794 = _1792 ^ _1793;
  wire _1795 = uncoded_block[276] ^ uncoded_block[277];
  wire _1796 = uncoded_block[279] ^ uncoded_block[283];
  wire _1797 = _1795 ^ _1796;
  wire _1798 = _1794 ^ _1797;
  wire _1799 = _1791 ^ _1798;
  wire _1800 = _1784 ^ _1799;
  wire _1801 = _1771 ^ _1800;
  wire _1802 = _1741 ^ _1801;
  wire _1803 = uncoded_block[284] ^ uncoded_block[285];
  wire _1804 = uncoded_block[288] ^ uncoded_block[291];
  wire _1805 = _1803 ^ _1804;
  wire _1806 = uncoded_block[296] ^ uncoded_block[297];
  wire _1807 = uncoded_block[298] ^ uncoded_block[299];
  wire _1808 = _1806 ^ _1807;
  wire _1809 = _1805 ^ _1808;
  wire _1810 = uncoded_block[300] ^ uncoded_block[301];
  wire _1811 = uncoded_block[302] ^ uncoded_block[308];
  wire _1812 = _1810 ^ _1811;
  wire _1813 = uncoded_block[310] ^ uncoded_block[317];
  wire _1814 = uncoded_block[318] ^ uncoded_block[319];
  wire _1815 = _1813 ^ _1814;
  wire _1816 = _1812 ^ _1815;
  wire _1817 = _1809 ^ _1816;
  wire _1818 = uncoded_block[320] ^ uncoded_block[322];
  wire _1819 = uncoded_block[326] ^ uncoded_block[330];
  wire _1820 = _1818 ^ _1819;
  wire _1821 = uncoded_block[332] ^ uncoded_block[333];
  wire _1822 = uncoded_block[334] ^ uncoded_block[337];
  wire _1823 = _1821 ^ _1822;
  wire _1824 = _1820 ^ _1823;
  wire _1825 = uncoded_block[338] ^ uncoded_block[339];
  wire _1826 = uncoded_block[341] ^ uncoded_block[344];
  wire _1827 = _1825 ^ _1826;
  wire _1828 = _159 ^ _161;
  wire _1829 = _1827 ^ _1828;
  wire _1830 = _1824 ^ _1829;
  wire _1831 = _1817 ^ _1830;
  wire _1832 = uncoded_block[350] ^ uncoded_block[355];
  wire _1833 = uncoded_block[356] ^ uncoded_block[360];
  wire _1834 = _1832 ^ _1833;
  wire _1835 = uncoded_block[367] ^ uncoded_block[368];
  wire _1836 = _168 ^ _1835;
  wire _1837 = _1834 ^ _1836;
  wire _1838 = uncoded_block[370] ^ uncoded_block[371];
  wire _1839 = uncoded_block[372] ^ uncoded_block[377];
  wire _1840 = _1838 ^ _1839;
  wire _1841 = uncoded_block[380] ^ uncoded_block[381];
  wire _1842 = uncoded_block[382] ^ uncoded_block[384];
  wire _1843 = _1841 ^ _1842;
  wire _1844 = _1840 ^ _1843;
  wire _1845 = _1837 ^ _1844;
  wire _1846 = uncoded_block[386] ^ uncoded_block[390];
  wire _1847 = uncoded_block[394] ^ uncoded_block[395];
  wire _1848 = _1846 ^ _1847;
  wire _1849 = uncoded_block[397] ^ uncoded_block[399];
  wire _1850 = uncoded_block[401] ^ uncoded_block[407];
  wire _1851 = _1849 ^ _1850;
  wire _1852 = _1848 ^ _1851;
  wire _1853 = uncoded_block[409] ^ uncoded_block[415];
  wire _1854 = uncoded_block[417] ^ uncoded_block[421];
  wire _1855 = _1853 ^ _1854;
  wire _1856 = uncoded_block[423] ^ uncoded_block[430];
  wire _1857 = uncoded_block[432] ^ uncoded_block[433];
  wire _1858 = _1856 ^ _1857;
  wire _1859 = _1855 ^ _1858;
  wire _1860 = _1852 ^ _1859;
  wire _1861 = _1845 ^ _1860;
  wire _1862 = _1831 ^ _1861;
  wire _1863 = uncoded_block[439] ^ uncoded_block[441];
  wire _1864 = uncoded_block[444] ^ uncoded_block[446];
  wire _1865 = _1863 ^ _1864;
  wire _1866 = uncoded_block[448] ^ uncoded_block[451];
  wire _1867 = uncoded_block[453] ^ uncoded_block[455];
  wire _1868 = _1866 ^ _1867;
  wire _1869 = _1865 ^ _1868;
  wire _1870 = uncoded_block[456] ^ uncoded_block[457];
  wire _1871 = uncoded_block[458] ^ uncoded_block[460];
  wire _1872 = _1870 ^ _1871;
  wire _1873 = uncoded_block[461] ^ uncoded_block[464];
  wire _1874 = uncoded_block[465] ^ uncoded_block[467];
  wire _1875 = _1873 ^ _1874;
  wire _1876 = _1872 ^ _1875;
  wire _1877 = _1869 ^ _1876;
  wire _1878 = uncoded_block[468] ^ uncoded_block[469];
  wire _1879 = uncoded_block[471] ^ uncoded_block[473];
  wire _1880 = _1878 ^ _1879;
  wire _1881 = uncoded_block[474] ^ uncoded_block[479];
  wire _1882 = uncoded_block[480] ^ uncoded_block[485];
  wire _1883 = _1881 ^ _1882;
  wire _1884 = _1880 ^ _1883;
  wire _1885 = uncoded_block[491] ^ uncoded_block[496];
  wire _1886 = _224 ^ _1885;
  wire _1887 = uncoded_block[503] ^ uncoded_block[505];
  wire _1888 = _228 ^ _1887;
  wire _1889 = _1886 ^ _1888;
  wire _1890 = _1884 ^ _1889;
  wire _1891 = _1877 ^ _1890;
  wire _1892 = uncoded_block[506] ^ uncoded_block[507];
  wire _1893 = uncoded_block[508] ^ uncoded_block[512];
  wire _1894 = _1892 ^ _1893;
  wire _1895 = uncoded_block[517] ^ uncoded_block[519];
  wire _1896 = _232 ^ _1895;
  wire _1897 = _1894 ^ _1896;
  wire _1898 = uncoded_block[522] ^ uncoded_block[524];
  wire _1899 = _1107 ^ _1898;
  wire _1900 = uncoded_block[526] ^ uncoded_block[527];
  wire _1901 = uncoded_block[529] ^ uncoded_block[531];
  wire _1902 = _1900 ^ _1901;
  wire _1903 = _1899 ^ _1902;
  wire _1904 = _1897 ^ _1903;
  wire _1905 = uncoded_block[534] ^ uncoded_block[535];
  wire _1906 = uncoded_block[536] ^ uncoded_block[542];
  wire _1907 = _1905 ^ _1906;
  wire _1908 = uncoded_block[543] ^ uncoded_block[544];
  wire _1909 = uncoded_block[545] ^ uncoded_block[546];
  wire _1910 = _1908 ^ _1909;
  wire _1911 = _1907 ^ _1910;
  wire _1912 = uncoded_block[548] ^ uncoded_block[549];
  wire _1913 = uncoded_block[550] ^ uncoded_block[552];
  wire _1914 = _1912 ^ _1913;
  wire _1915 = uncoded_block[553] ^ uncoded_block[555];
  wire _1916 = uncoded_block[557] ^ uncoded_block[558];
  wire _1917 = _1915 ^ _1916;
  wire _1918 = _1914 ^ _1917;
  wire _1919 = _1911 ^ _1918;
  wire _1920 = _1904 ^ _1919;
  wire _1921 = _1891 ^ _1920;
  wire _1922 = _1862 ^ _1921;
  wire _1923 = _1802 ^ _1922;
  wire _1924 = uncoded_block[560] ^ uncoded_block[562];
  wire _1925 = uncoded_block[563] ^ uncoded_block[565];
  wire _1926 = _1924 ^ _1925;
  wire _1927 = uncoded_block[566] ^ uncoded_block[569];
  wire _1928 = uncoded_block[571] ^ uncoded_block[574];
  wire _1929 = _1927 ^ _1928;
  wire _1930 = _1926 ^ _1929;
  wire _1931 = uncoded_block[575] ^ uncoded_block[576];
  wire _1932 = _1931 ^ _263;
  wire _1933 = uncoded_block[583] ^ uncoded_block[584];
  wire _1934 = uncoded_block[585] ^ uncoded_block[589];
  wire _1935 = _1933 ^ _1934;
  wire _1936 = _1932 ^ _1935;
  wire _1937 = _1930 ^ _1936;
  wire _1938 = uncoded_block[592] ^ uncoded_block[593];
  wire _1939 = uncoded_block[595] ^ uncoded_block[596];
  wire _1940 = _1938 ^ _1939;
  wire _1941 = uncoded_block[600] ^ uncoded_block[604];
  wire _1942 = uncoded_block[607] ^ uncoded_block[608];
  wire _1943 = _1941 ^ _1942;
  wire _1944 = _1940 ^ _1943;
  wire _1945 = uncoded_block[613] ^ uncoded_block[617];
  wire _1946 = uncoded_block[620] ^ uncoded_block[621];
  wire _1947 = _1945 ^ _1946;
  wire _1948 = uncoded_block[623] ^ uncoded_block[625];
  wire _1949 = _1948 ^ _1154;
  wire _1950 = _1947 ^ _1949;
  wire _1951 = _1944 ^ _1950;
  wire _1952 = _1937 ^ _1951;
  wire _1953 = uncoded_block[629] ^ uncoded_block[631];
  wire _1954 = uncoded_block[634] ^ uncoded_block[639];
  wire _1955 = _1953 ^ _1954;
  wire _1956 = uncoded_block[640] ^ uncoded_block[645];
  wire _1957 = uncoded_block[646] ^ uncoded_block[650];
  wire _1958 = _1956 ^ _1957;
  wire _1959 = _1955 ^ _1958;
  wire _1960 = uncoded_block[651] ^ uncoded_block[652];
  wire _1961 = _1960 ^ _304;
  wire _1962 = uncoded_block[657] ^ uncoded_block[660];
  wire _1963 = uncoded_block[663] ^ uncoded_block[667];
  wire _1964 = _1962 ^ _1963;
  wire _1965 = _1961 ^ _1964;
  wire _1966 = _1959 ^ _1965;
  wire _1967 = _1174 ^ _1178;
  wire _1968 = uncoded_block[678] ^ uncoded_block[679];
  wire _1969 = _1180 ^ _1968;
  wire _1970 = _1967 ^ _1969;
  wire _1971 = uncoded_block[680] ^ uncoded_block[681];
  wire _1972 = uncoded_block[684] ^ uncoded_block[687];
  wire _1973 = _1971 ^ _1972;
  wire _1974 = uncoded_block[688] ^ uncoded_block[690];
  wire _1975 = uncoded_block[697] ^ uncoded_block[702];
  wire _1976 = _1974 ^ _1975;
  wire _1977 = _1973 ^ _1976;
  wire _1978 = _1970 ^ _1977;
  wire _1979 = _1966 ^ _1978;
  wire _1980 = _1952 ^ _1979;
  wire _1981 = uncoded_block[703] ^ uncoded_block[708];
  wire _1982 = _1981 ^ _1192;
  wire _1983 = uncoded_block[714] ^ uncoded_block[717];
  wire _1984 = uncoded_block[718] ^ uncoded_block[720];
  wire _1985 = _1983 ^ _1984;
  wire _1986 = _1982 ^ _1985;
  wire _1987 = uncoded_block[722] ^ uncoded_block[724];
  wire _1988 = uncoded_block[725] ^ uncoded_block[726];
  wire _1989 = _1987 ^ _1988;
  wire _1990 = uncoded_block[727] ^ uncoded_block[730];
  wire _1991 = uncoded_block[731] ^ uncoded_block[732];
  wire _1992 = _1990 ^ _1991;
  wire _1993 = _1989 ^ _1992;
  wire _1994 = _1986 ^ _1993;
  wire _1995 = uncoded_block[735] ^ uncoded_block[736];
  wire _1996 = uncoded_block[738] ^ uncoded_block[739];
  wire _1997 = _1995 ^ _1996;
  wire _1998 = uncoded_block[743] ^ uncoded_block[745];
  wire _1999 = uncoded_block[746] ^ uncoded_block[747];
  wire _2000 = _1998 ^ _1999;
  wire _2001 = _1997 ^ _2000;
  wire _2002 = uncoded_block[750] ^ uncoded_block[751];
  wire _2003 = uncoded_block[754] ^ uncoded_block[755];
  wire _2004 = _2002 ^ _2003;
  wire _2005 = uncoded_block[757] ^ uncoded_block[759];
  wire _2006 = uncoded_block[761] ^ uncoded_block[764];
  wire _2007 = _2005 ^ _2006;
  wire _2008 = _2004 ^ _2007;
  wire _2009 = _2001 ^ _2008;
  wire _2010 = _1994 ^ _2009;
  wire _2011 = uncoded_block[765] ^ uncoded_block[771];
  wire _2012 = uncoded_block[773] ^ uncoded_block[775];
  wire _2013 = _2011 ^ _2012;
  wire _2014 = uncoded_block[776] ^ uncoded_block[777];
  wire _2015 = uncoded_block[782] ^ uncoded_block[783];
  wire _2016 = _2014 ^ _2015;
  wire _2017 = _2013 ^ _2016;
  wire _2018 = uncoded_block[785] ^ uncoded_block[787];
  wire _2019 = uncoded_block[790] ^ uncoded_block[791];
  wire _2020 = _2018 ^ _2019;
  wire _2021 = uncoded_block[794] ^ uncoded_block[797];
  wire _2022 = uncoded_block[798] ^ uncoded_block[801];
  wire _2023 = _2021 ^ _2022;
  wire _2024 = _2020 ^ _2023;
  wire _2025 = _2017 ^ _2024;
  wire _2026 = uncoded_block[812] ^ uncoded_block[813];
  wire _2027 = _1235 ^ _2026;
  wire _2028 = uncoded_block[818] ^ uncoded_block[819];
  wire _2029 = uncoded_block[820] ^ uncoded_block[821];
  wire _2030 = _2028 ^ _2029;
  wire _2031 = _2027 ^ _2030;
  wire _2032 = uncoded_block[826] ^ uncoded_block[827];
  wire _2033 = uncoded_block[831] ^ uncoded_block[833];
  wire _2034 = _2032 ^ _2033;
  wire _2035 = uncoded_block[837] ^ uncoded_block[838];
  wire _2036 = uncoded_block[841] ^ uncoded_block[842];
  wire _2037 = _2035 ^ _2036;
  wire _2038 = _2034 ^ _2037;
  wire _2039 = _2031 ^ _2038;
  wire _2040 = _2025 ^ _2039;
  wire _2041 = _2010 ^ _2040;
  wire _2042 = _1980 ^ _2041;
  wire _2043 = uncoded_block[844] ^ uncoded_block[847];
  wire _2044 = uncoded_block[849] ^ uncoded_block[852];
  wire _2045 = _2043 ^ _2044;
  wire _2046 = uncoded_block[854] ^ uncoded_block[855];
  wire _2047 = uncoded_block[857] ^ uncoded_block[860];
  wire _2048 = _2046 ^ _2047;
  wire _2049 = _2045 ^ _2048;
  wire _2050 = uncoded_block[861] ^ uncoded_block[869];
  wire _2051 = uncoded_block[870] ^ uncoded_block[877];
  wire _2052 = _2050 ^ _2051;
  wire _2053 = uncoded_block[878] ^ uncoded_block[880];
  wire _2054 = uncoded_block[881] ^ uncoded_block[884];
  wire _2055 = _2053 ^ _2054;
  wire _2056 = _2052 ^ _2055;
  wire _2057 = _2049 ^ _2056;
  wire _2058 = uncoded_block[885] ^ uncoded_block[886];
  wire _2059 = uncoded_block[887] ^ uncoded_block[889];
  wire _2060 = _2058 ^ _2059;
  wire _2061 = uncoded_block[890] ^ uncoded_block[891];
  wire _2062 = uncoded_block[893] ^ uncoded_block[896];
  wire _2063 = _2061 ^ _2062;
  wire _2064 = _2060 ^ _2063;
  wire _2065 = uncoded_block[903] ^ uncoded_block[904];
  wire _2066 = _2065 ^ _1281;
  wire _2067 = _430 ^ _2066;
  wire _2068 = _2064 ^ _2067;
  wire _2069 = _2057 ^ _2068;
  wire _2070 = uncoded_block[908] ^ uncoded_block[909];
  wire _2071 = uncoded_block[910] ^ uncoded_block[911];
  wire _2072 = _2070 ^ _2071;
  wire _2073 = uncoded_block[921] ^ uncoded_block[923];
  wire _2074 = _1288 ^ _2073;
  wire _2075 = _2072 ^ _2074;
  wire _2076 = uncoded_block[924] ^ uncoded_block[925];
  wire _2077 = _2076 ^ _1296;
  wire _2078 = uncoded_block[932] ^ uncoded_block[933];
  wire _2079 = uncoded_block[934] ^ uncoded_block[935];
  wire _2080 = _2078 ^ _2079;
  wire _2081 = _2077 ^ _2080;
  wire _2082 = _2075 ^ _2081;
  wire _2083 = uncoded_block[937] ^ uncoded_block[939];
  wire _2084 = uncoded_block[940] ^ uncoded_block[943];
  wire _2085 = _2083 ^ _2084;
  wire _2086 = uncoded_block[945] ^ uncoded_block[946];
  wire _2087 = _2086 ^ _460;
  wire _2088 = _2085 ^ _2087;
  wire _2089 = uncoded_block[953] ^ uncoded_block[955];
  wire _2090 = uncoded_block[957] ^ uncoded_block[958];
  wire _2091 = _2089 ^ _2090;
  wire _2092 = uncoded_block[965] ^ uncoded_block[966];
  wire _2093 = uncoded_block[967] ^ uncoded_block[968];
  wire _2094 = _2092 ^ _2093;
  wire _2095 = _2091 ^ _2094;
  wire _2096 = _2088 ^ _2095;
  wire _2097 = _2082 ^ _2096;
  wire _2098 = _2069 ^ _2097;
  wire _2099 = uncoded_block[972] ^ uncoded_block[978];
  wire _2100 = uncoded_block[979] ^ uncoded_block[980];
  wire _2101 = _2099 ^ _2100;
  wire _2102 = uncoded_block[985] ^ uncoded_block[987];
  wire _2103 = _476 ^ _2102;
  wire _2104 = _2101 ^ _2103;
  wire _2105 = uncoded_block[988] ^ uncoded_block[992];
  wire _2106 = _2105 ^ _479;
  wire _2107 = uncoded_block[999] ^ uncoded_block[1000];
  wire _2108 = _480 ^ _2107;
  wire _2109 = _2106 ^ _2108;
  wire _2110 = _2104 ^ _2109;
  wire _2111 = uncoded_block[1001] ^ uncoded_block[1002];
  wire _2112 = uncoded_block[1003] ^ uncoded_block[1004];
  wire _2113 = _2111 ^ _2112;
  wire _2114 = uncoded_block[1005] ^ uncoded_block[1006];
  wire _2115 = _2114 ^ _487;
  wire _2116 = _2113 ^ _2115;
  wire _2117 = uncoded_block[1013] ^ uncoded_block[1014];
  wire _2118 = uncoded_block[1015] ^ uncoded_block[1018];
  wire _2119 = _2117 ^ _2118;
  wire _2120 = uncoded_block[1020] ^ uncoded_block[1021];
  wire _2121 = uncoded_block[1024] ^ uncoded_block[1027];
  wire _2122 = _2120 ^ _2121;
  wire _2123 = _2119 ^ _2122;
  wire _2124 = _2116 ^ _2123;
  wire _2125 = _2110 ^ _2124;
  wire _2126 = uncoded_block[1028] ^ uncoded_block[1031];
  wire _2127 = uncoded_block[1033] ^ uncoded_block[1034];
  wire _2128 = _2126 ^ _2127;
  wire _2129 = uncoded_block[1037] ^ uncoded_block[1038];
  wire _2130 = uncoded_block[1043] ^ uncoded_block[1044];
  wire _2131 = _2129 ^ _2130;
  wire _2132 = _2128 ^ _2131;
  wire _2133 = uncoded_block[1045] ^ uncoded_block[1046];
  wire _2134 = uncoded_block[1048] ^ uncoded_block[1049];
  wire _2135 = _2133 ^ _2134;
  wire _2136 = uncoded_block[1051] ^ uncoded_block[1052];
  wire _2137 = _2136 ^ _519;
  wire _2138 = _2135 ^ _2137;
  wire _2139 = _2132 ^ _2138;
  wire _2140 = uncoded_block[1061] ^ uncoded_block[1063];
  wire _2141 = _1363 ^ _2140;
  wire _2142 = uncoded_block[1064] ^ uncoded_block[1066];
  wire _2143 = uncoded_block[1070] ^ uncoded_block[1072];
  wire _2144 = _2142 ^ _2143;
  wire _2145 = _2141 ^ _2144;
  wire _2146 = uncoded_block[1074] ^ uncoded_block[1075];
  wire _2147 = uncoded_block[1076] ^ uncoded_block[1078];
  wire _2148 = _2146 ^ _2147;
  wire _2149 = uncoded_block[1087] ^ uncoded_block[1088];
  wire _2150 = _533 ^ _2149;
  wire _2151 = _2148 ^ _2150;
  wire _2152 = _2145 ^ _2151;
  wire _2153 = _2139 ^ _2152;
  wire _2154 = _2125 ^ _2153;
  wire _2155 = _2098 ^ _2154;
  wire _2156 = _2042 ^ _2155;
  wire _2157 = _1923 ^ _2156;
  wire _2158 = uncoded_block[1094] ^ uncoded_block[1102];
  wire _2159 = _536 ^ _2158;
  wire _2160 = uncoded_block[1103] ^ uncoded_block[1104];
  wire _2161 = uncoded_block[1105] ^ uncoded_block[1106];
  wire _2162 = _2160 ^ _2161;
  wire _2163 = _2159 ^ _2162;
  wire _2164 = uncoded_block[1108] ^ uncoded_block[1109];
  wire _2165 = uncoded_block[1110] ^ uncoded_block[1112];
  wire _2166 = _2164 ^ _2165;
  wire _2167 = uncoded_block[1114] ^ uncoded_block[1117];
  wire _2168 = uncoded_block[1118] ^ uncoded_block[1122];
  wire _2169 = _2167 ^ _2168;
  wire _2170 = _2166 ^ _2169;
  wire _2171 = _2163 ^ _2170;
  wire _2172 = uncoded_block[1123] ^ uncoded_block[1125];
  wire _2173 = _2172 ^ _558;
  wire _2174 = uncoded_block[1132] ^ uncoded_block[1135];
  wire _2175 = _560 ^ _2174;
  wire _2176 = _2173 ^ _2175;
  wire _2177 = uncoded_block[1136] ^ uncoded_block[1139];
  wire _2178 = _2177 ^ _567;
  wire _2179 = uncoded_block[1143] ^ uncoded_block[1144];
  wire _2180 = uncoded_block[1145] ^ uncoded_block[1148];
  wire _2181 = _2179 ^ _2180;
  wire _2182 = _2178 ^ _2181;
  wire _2183 = _2176 ^ _2182;
  wire _2184 = _2171 ^ _2183;
  wire _2185 = uncoded_block[1151] ^ uncoded_block[1152];
  wire _2186 = uncoded_block[1153] ^ uncoded_block[1155];
  wire _2187 = _2185 ^ _2186;
  wire _2188 = uncoded_block[1159] ^ uncoded_block[1162];
  wire _2189 = uncoded_block[1167] ^ uncoded_block[1169];
  wire _2190 = _2188 ^ _2189;
  wire _2191 = _2187 ^ _2190;
  wire _2192 = uncoded_block[1172] ^ uncoded_block[1175];
  wire _2193 = uncoded_block[1177] ^ uncoded_block[1180];
  wire _2194 = _2192 ^ _2193;
  wire _2195 = uncoded_block[1181] ^ uncoded_block[1182];
  wire _2196 = uncoded_block[1184] ^ uncoded_block[1186];
  wire _2197 = _2195 ^ _2196;
  wire _2198 = _2194 ^ _2197;
  wire _2199 = _2191 ^ _2198;
  wire _2200 = uncoded_block[1187] ^ uncoded_block[1188];
  wire _2201 = uncoded_block[1189] ^ uncoded_block[1190];
  wire _2202 = _2200 ^ _2201;
  wire _2203 = uncoded_block[1194] ^ uncoded_block[1198];
  wire _2204 = _1420 ^ _2203;
  wire _2205 = _2202 ^ _2204;
  wire _2206 = uncoded_block[1199] ^ uncoded_block[1200];
  wire _2207 = uncoded_block[1201] ^ uncoded_block[1202];
  wire _2208 = _2206 ^ _2207;
  wire _2209 = uncoded_block[1203] ^ uncoded_block[1204];
  wire _2210 = uncoded_block[1205] ^ uncoded_block[1206];
  wire _2211 = _2209 ^ _2210;
  wire _2212 = _2208 ^ _2211;
  wire _2213 = _2205 ^ _2212;
  wire _2214 = _2199 ^ _2213;
  wire _2215 = _2184 ^ _2214;
  wire _2216 = uncoded_block[1207] ^ uncoded_block[1208];
  wire _2217 = uncoded_block[1209] ^ uncoded_block[1210];
  wire _2218 = _2216 ^ _2217;
  wire _2219 = uncoded_block[1215] ^ uncoded_block[1216];
  wire _2220 = uncoded_block[1217] ^ uncoded_block[1219];
  wire _2221 = _2219 ^ _2220;
  wire _2222 = _2218 ^ _2221;
  wire _2223 = uncoded_block[1221] ^ uncoded_block[1226];
  wire _2224 = _2223 ^ _1436;
  wire _2225 = uncoded_block[1231] ^ uncoded_block[1232];
  wire _2226 = uncoded_block[1234] ^ uncoded_block[1236];
  wire _2227 = _2225 ^ _2226;
  wire _2228 = _2224 ^ _2227;
  wire _2229 = _2222 ^ _2228;
  wire _2230 = uncoded_block[1238] ^ uncoded_block[1240];
  wire _2231 = _2230 ^ _1448;
  wire _2232 = uncoded_block[1247] ^ uncoded_block[1248];
  wire _2233 = _2232 ^ _621;
  wire _2234 = _2231 ^ _2233;
  wire _2235 = uncoded_block[1253] ^ uncoded_block[1254];
  wire _2236 = uncoded_block[1256] ^ uncoded_block[1259];
  wire _2237 = _2235 ^ _2236;
  wire _2238 = uncoded_block[1260] ^ uncoded_block[1262];
  wire _2239 = uncoded_block[1266] ^ uncoded_block[1267];
  wire _2240 = _2238 ^ _2239;
  wire _2241 = _2237 ^ _2240;
  wire _2242 = _2234 ^ _2241;
  wire _2243 = _2229 ^ _2242;
  wire _2244 = uncoded_block[1268] ^ uncoded_block[1269];
  wire _2245 = uncoded_block[1270] ^ uncoded_block[1271];
  wire _2246 = _2244 ^ _2245;
  wire _2247 = uncoded_block[1276] ^ uncoded_block[1278];
  wire _2248 = uncoded_block[1280] ^ uncoded_block[1283];
  wire _2249 = _2247 ^ _2248;
  wire _2250 = _2246 ^ _2249;
  wire _2251 = uncoded_block[1286] ^ uncoded_block[1293];
  wire _2252 = uncoded_block[1294] ^ uncoded_block[1299];
  wire _2253 = _2251 ^ _2252;
  wire _2254 = uncoded_block[1302] ^ uncoded_block[1303];
  wire _2255 = uncoded_block[1304] ^ uncoded_block[1305];
  wire _2256 = _2254 ^ _2255;
  wire _2257 = _2253 ^ _2256;
  wire _2258 = _2250 ^ _2257;
  wire _2259 = uncoded_block[1306] ^ uncoded_block[1308];
  wire _2260 = _2259 ^ _1480;
  wire _2261 = uncoded_block[1313] ^ uncoded_block[1314];
  wire _2262 = uncoded_block[1316] ^ uncoded_block[1317];
  wire _2263 = _2261 ^ _2262;
  wire _2264 = _2260 ^ _2263;
  wire _2265 = uncoded_block[1319] ^ uncoded_block[1322];
  wire _2266 = uncoded_block[1325] ^ uncoded_block[1328];
  wire _2267 = _2265 ^ _2266;
  wire _2268 = uncoded_block[1329] ^ uncoded_block[1330];
  wire _2269 = uncoded_block[1331] ^ uncoded_block[1335];
  wire _2270 = _2268 ^ _2269;
  wire _2271 = _2267 ^ _2270;
  wire _2272 = _2264 ^ _2271;
  wire _2273 = _2258 ^ _2272;
  wire _2274 = _2243 ^ _2273;
  wire _2275 = _2215 ^ _2274;
  wire _2276 = uncoded_block[1336] ^ uncoded_block[1338];
  wire _2277 = uncoded_block[1339] ^ uncoded_block[1341];
  wire _2278 = _2276 ^ _2277;
  wire _2279 = uncoded_block[1343] ^ uncoded_block[1352];
  wire _2280 = uncoded_block[1354] ^ uncoded_block[1359];
  wire _2281 = _2279 ^ _2280;
  wire _2282 = _2278 ^ _2281;
  wire _2283 = uncoded_block[1364] ^ uncoded_block[1365];
  wire _2284 = uncoded_block[1366] ^ uncoded_block[1367];
  wire _2285 = _2283 ^ _2284;
  wire _2286 = _680 ^ _684;
  wire _2287 = _2285 ^ _2286;
  wire _2288 = _2282 ^ _2287;
  wire _2289 = uncoded_block[1374] ^ uncoded_block[1375];
  wire _2290 = uncoded_block[1378] ^ uncoded_block[1379];
  wire _2291 = _2289 ^ _2290;
  wire _2292 = uncoded_block[1380] ^ uncoded_block[1387];
  wire _2293 = uncoded_block[1390] ^ uncoded_block[1392];
  wire _2294 = _2292 ^ _2293;
  wire _2295 = _2291 ^ _2294;
  wire _2296 = uncoded_block[1397] ^ uncoded_block[1399];
  wire _2297 = uncoded_block[1400] ^ uncoded_block[1401];
  wire _2298 = _2296 ^ _2297;
  wire _2299 = uncoded_block[1402] ^ uncoded_block[1403];
  wire _2300 = uncoded_block[1406] ^ uncoded_block[1407];
  wire _2301 = _2299 ^ _2300;
  wire _2302 = _2298 ^ _2301;
  wire _2303 = _2295 ^ _2302;
  wire _2304 = _2288 ^ _2303;
  wire _2305 = uncoded_block[1408] ^ uncoded_block[1414];
  wire _2306 = uncoded_block[1416] ^ uncoded_block[1417];
  wire _2307 = _2305 ^ _2306;
  wire _2308 = uncoded_block[1425] ^ uncoded_block[1426];
  wire _2309 = _708 ^ _2308;
  wire _2310 = _2307 ^ _2309;
  wire _2311 = uncoded_block[1427] ^ uncoded_block[1428];
  wire _2312 = _2311 ^ _1531;
  wire _2313 = uncoded_block[1433] ^ uncoded_block[1434];
  wire _2314 = uncoded_block[1435] ^ uncoded_block[1436];
  wire _2315 = _2313 ^ _2314;
  wire _2316 = _2312 ^ _2315;
  wire _2317 = _2310 ^ _2316;
  wire _2318 = uncoded_block[1438] ^ uncoded_block[1439];
  wire _2319 = uncoded_block[1441] ^ uncoded_block[1442];
  wire _2320 = _2318 ^ _2319;
  wire _2321 = uncoded_block[1443] ^ uncoded_block[1444];
  wire _2322 = uncoded_block[1446] ^ uncoded_block[1447];
  wire _2323 = _2321 ^ _2322;
  wire _2324 = _2320 ^ _2323;
  wire _2325 = uncoded_block[1448] ^ uncoded_block[1449];
  wire _2326 = uncoded_block[1451] ^ uncoded_block[1452];
  wire _2327 = _2325 ^ _2326;
  wire _2328 = uncoded_block[1453] ^ uncoded_block[1454];
  wire _2329 = uncoded_block[1456] ^ uncoded_block[1458];
  wire _2330 = _2328 ^ _2329;
  wire _2331 = _2327 ^ _2330;
  wire _2332 = _2324 ^ _2331;
  wire _2333 = _2317 ^ _2332;
  wire _2334 = _2304 ^ _2333;
  wire _2335 = uncoded_block[1459] ^ uncoded_block[1461];
  wire _2336 = uncoded_block[1462] ^ uncoded_block[1463];
  wire _2337 = _2335 ^ _2336;
  wire _2338 = uncoded_block[1468] ^ uncoded_block[1470];
  wire _2339 = _1548 ^ _2338;
  wire _2340 = _2337 ^ _2339;
  wire _2341 = uncoded_block[1471] ^ uncoded_block[1476];
  wire _2342 = uncoded_block[1477] ^ uncoded_block[1478];
  wire _2343 = _2341 ^ _2342;
  wire _2344 = uncoded_block[1479] ^ uncoded_block[1481];
  wire _2345 = uncoded_block[1482] ^ uncoded_block[1484];
  wire _2346 = _2344 ^ _2345;
  wire _2347 = _2343 ^ _2346;
  wire _2348 = _2340 ^ _2347;
  wire _2349 = uncoded_block[1487] ^ uncoded_block[1488];
  wire _2350 = uncoded_block[1493] ^ uncoded_block[1496];
  wire _2351 = _2349 ^ _2350;
  wire _2352 = uncoded_block[1497] ^ uncoded_block[1498];
  wire _2353 = uncoded_block[1502] ^ uncoded_block[1510];
  wire _2354 = _2352 ^ _2353;
  wire _2355 = _2351 ^ _2354;
  wire _2356 = uncoded_block[1512] ^ uncoded_block[1517];
  wire _2357 = uncoded_block[1520] ^ uncoded_block[1521];
  wire _2358 = _2356 ^ _2357;
  wire _2359 = uncoded_block[1523] ^ uncoded_block[1526];
  wire _2360 = uncoded_block[1528] ^ uncoded_block[1530];
  wire _2361 = _2359 ^ _2360;
  wire _2362 = _2358 ^ _2361;
  wire _2363 = _2355 ^ _2362;
  wire _2364 = _2348 ^ _2363;
  wire _2365 = uncoded_block[1537] ^ uncoded_block[1540];
  wire _2366 = _1586 ^ _2365;
  wire _2367 = uncoded_block[1546] ^ uncoded_block[1547];
  wire _2368 = _1590 ^ _2367;
  wire _2369 = _2366 ^ _2368;
  wire _2370 = uncoded_block[1548] ^ uncoded_block[1551];
  wire _2371 = _2370 ^ _769;
  wire _2372 = uncoded_block[1562] ^ uncoded_block[1563];
  wire _2373 = _770 ^ _2372;
  wire _2374 = _2371 ^ _2373;
  wire _2375 = _2369 ^ _2374;
  wire _2376 = uncoded_block[1564] ^ uncoded_block[1565];
  wire _2377 = uncoded_block[1568] ^ uncoded_block[1569];
  wire _2378 = _2376 ^ _2377;
  wire _2379 = uncoded_block[1570] ^ uncoded_block[1574];
  wire _2380 = uncoded_block[1575] ^ uncoded_block[1578];
  wire _2381 = _2379 ^ _2380;
  wire _2382 = _2378 ^ _2381;
  wire _2383 = uncoded_block[1579] ^ uncoded_block[1580];
  wire _2384 = uncoded_block[1582] ^ uncoded_block[1584];
  wire _2385 = _2383 ^ _2384;
  wire _2386 = uncoded_block[1585] ^ uncoded_block[1586];
  wire _2387 = _2386 ^ _1616;
  wire _2388 = _2385 ^ _2387;
  wire _2389 = _2382 ^ _2388;
  wire _2390 = _2375 ^ _2389;
  wire _2391 = _2364 ^ _2390;
  wire _2392 = _2334 ^ _2391;
  wire _2393 = _2275 ^ _2392;
  wire _2394 = uncoded_block[1593] ^ uncoded_block[1595];
  wire _2395 = _2394 ^ _1620;
  wire _2396 = uncoded_block[1607] ^ uncoded_block[1608];
  wire _2397 = _1625 ^ _2396;
  wire _2398 = _2395 ^ _2397;
  wire _2399 = _801 ^ _1632;
  wire _2400 = uncoded_block[1624] ^ uncoded_block[1628];
  wire _2401 = _804 ^ _2400;
  wire _2402 = _2399 ^ _2401;
  wire _2403 = _2398 ^ _2402;
  wire _2404 = uncoded_block[1629] ^ uncoded_block[1631];
  wire _2405 = uncoded_block[1634] ^ uncoded_block[1636];
  wire _2406 = _2404 ^ _2405;
  wire _2407 = uncoded_block[1637] ^ uncoded_block[1640];
  wire _2408 = uncoded_block[1641] ^ uncoded_block[1642];
  wire _2409 = _2407 ^ _2408;
  wire _2410 = _2406 ^ _2409;
  wire _2411 = uncoded_block[1643] ^ uncoded_block[1646];
  wire _2412 = uncoded_block[1647] ^ uncoded_block[1648];
  wire _2413 = _2411 ^ _2412;
  wire _2414 = uncoded_block[1656] ^ uncoded_block[1660];
  wire _2415 = _1650 ^ _2414;
  wire _2416 = _2413 ^ _2415;
  wire _2417 = _2410 ^ _2416;
  wire _2418 = _2403 ^ _2417;
  wire _2419 = uncoded_block[1662] ^ uncoded_block[1663];
  wire _2420 = uncoded_block[1665] ^ uncoded_block[1667];
  wire _2421 = _2419 ^ _2420;
  wire _2422 = uncoded_block[1668] ^ uncoded_block[1669];
  wire _2423 = uncoded_block[1671] ^ uncoded_block[1673];
  wire _2424 = _2422 ^ _2423;
  wire _2425 = _2421 ^ _2424;
  wire _2426 = uncoded_block[1677] ^ uncoded_block[1681];
  wire _2427 = uncoded_block[1682] ^ uncoded_block[1685];
  wire _2428 = _2426 ^ _2427;
  wire _2429 = uncoded_block[1688] ^ uncoded_block[1690];
  wire _2430 = uncoded_block[1694] ^ uncoded_block[1698];
  wire _2431 = _2429 ^ _2430;
  wire _2432 = _2428 ^ _2431;
  wire _2433 = _2425 ^ _2432;
  wire _2434 = uncoded_block[1700] ^ uncoded_block[1705];
  wire _2435 = uncoded_block[1706] ^ uncoded_block[1707];
  wire _2436 = _2434 ^ _2435;
  wire _2437 = uncoded_block[1708] ^ uncoded_block[1709];
  wire _2438 = uncoded_block[1710] ^ uncoded_block[1711];
  wire _2439 = _2437 ^ _2438;
  wire _2440 = _2436 ^ _2439;
  wire _2441 = uncoded_block[1715] ^ uncoded_block[1716];
  wire _2442 = _852 ^ _2441;
  wire _2443 = uncoded_block[1717] ^ uncoded_block[1718];
  wire _2444 = uncoded_block[1719] ^ uncoded_block[1721];
  wire _2445 = _2443 ^ _2444;
  wire _2446 = _2442 ^ _2445;
  wire _2447 = _2440 ^ _2446;
  wire _2448 = _2433 ^ _2447;
  wire _2449 = _2418 ^ _2448;
  wire _2450 = _2449 ^ uncoded_block[1722];
  wire _2451 = _2393 ^ _2450;
  wire _2452 = _2157 ^ _2451;
  wire _2453 = uncoded_block[3] ^ uncoded_block[7];
  wire _2454 = uncoded_block[9] ^ uncoded_block[12];
  wire _2455 = _2453 ^ _2454;
  wire _2456 = _868 ^ _871;
  wire _2457 = _2455 ^ _2456;
  wire _2458 = uncoded_block[19] ^ uncoded_block[21];
  wire _2459 = uncoded_block[23] ^ uncoded_block[28];
  wire _2460 = _2458 ^ _2459;
  wire _2461 = uncoded_block[29] ^ uncoded_block[31];
  wire _2462 = uncoded_block[33] ^ uncoded_block[37];
  wire _2463 = _2461 ^ _2462;
  wire _2464 = _2460 ^ _2463;
  wire _2465 = _2457 ^ _2464;
  wire _2466 = uncoded_block[38] ^ uncoded_block[39];
  wire _2467 = _2466 ^ _882;
  wire _2468 = uncoded_block[45] ^ uncoded_block[49];
  wire _2469 = _22 ^ _2468;
  wire _2470 = _2467 ^ _2469;
  wire _2471 = uncoded_block[56] ^ uncoded_block[58];
  wire _2472 = uncoded_block[60] ^ uncoded_block[61];
  wire _2473 = _2471 ^ _2472;
  wire _2474 = uncoded_block[62] ^ uncoded_block[63];
  wire _2475 = uncoded_block[65] ^ uncoded_block[68];
  wire _2476 = _2474 ^ _2475;
  wire _2477 = _2473 ^ _2476;
  wire _2478 = _2470 ^ _2477;
  wire _2479 = _2465 ^ _2478;
  wire _2480 = uncoded_block[69] ^ uncoded_block[73];
  wire _2481 = uncoded_block[78] ^ uncoded_block[79];
  wire _2482 = _2480 ^ _2481;
  wire _2483 = uncoded_block[82] ^ uncoded_block[85];
  wire _2484 = uncoded_block[86] ^ uncoded_block[87];
  wire _2485 = _2483 ^ _2484;
  wire _2486 = _2482 ^ _2485;
  wire _2487 = uncoded_block[88] ^ uncoded_block[90];
  wire _2488 = uncoded_block[92] ^ uncoded_block[103];
  wire _2489 = _2487 ^ _2488;
  wire _2490 = uncoded_block[104] ^ uncoded_block[106];
  wire _2491 = uncoded_block[108] ^ uncoded_block[109];
  wire _2492 = _2490 ^ _2491;
  wire _2493 = _2489 ^ _2492;
  wire _2494 = _2486 ^ _2493;
  wire _2495 = uncoded_block[115] ^ uncoded_block[116];
  wire _2496 = _1726 ^ _2495;
  wire _2497 = uncoded_block[117] ^ uncoded_block[118];
  wire _2498 = uncoded_block[119] ^ uncoded_block[120];
  wire _2499 = _2497 ^ _2498;
  wire _2500 = _2496 ^ _2499;
  wire _2501 = uncoded_block[121] ^ uncoded_block[122];
  wire _2502 = uncoded_block[124] ^ uncoded_block[125];
  wire _2503 = _2501 ^ _2502;
  wire _2504 = uncoded_block[129] ^ uncoded_block[133];
  wire _2505 = _1733 ^ _2504;
  wire _2506 = _2503 ^ _2505;
  wire _2507 = _2500 ^ _2506;
  wire _2508 = _2494 ^ _2507;
  wire _2509 = _2479 ^ _2508;
  wire _2510 = uncoded_block[136] ^ uncoded_block[138];
  wire _2511 = uncoded_block[143] ^ uncoded_block[145];
  wire _2512 = _2510 ^ _2511;
  wire _2513 = _2512 ^ _1746;
  wire _2514 = uncoded_block[155] ^ uncoded_block[160];
  wire _2515 = _2514 ^ _74;
  wire _2516 = uncoded_block[164] ^ uncoded_block[166];
  wire _2517 = uncoded_block[167] ^ uncoded_block[170];
  wire _2518 = _2516 ^ _2517;
  wire _2519 = _2515 ^ _2518;
  wire _2520 = _2513 ^ _2519;
  wire _2521 = uncoded_block[171] ^ uncoded_block[172];
  wire _2522 = uncoded_block[173] ^ uncoded_block[175];
  wire _2523 = _2521 ^ _2522;
  wire _2524 = uncoded_block[176] ^ uncoded_block[179];
  wire _2525 = uncoded_block[181] ^ uncoded_block[183];
  wire _2526 = _2524 ^ _2525;
  wire _2527 = _2523 ^ _2526;
  wire _2528 = uncoded_block[184] ^ uncoded_block[185];
  wire _2529 = uncoded_block[188] ^ uncoded_block[191];
  wire _2530 = _2528 ^ _2529;
  wire _2531 = uncoded_block[192] ^ uncoded_block[194];
  wire _2532 = uncoded_block[196] ^ uncoded_block[198];
  wire _2533 = _2531 ^ _2532;
  wire _2534 = _2530 ^ _2533;
  wire _2535 = _2527 ^ _2534;
  wire _2536 = _2520 ^ _2535;
  wire _2537 = uncoded_block[199] ^ uncoded_block[203];
  wire _2538 = uncoded_block[205] ^ uncoded_block[211];
  wire _2539 = _2537 ^ _2538;
  wire _2540 = uncoded_block[212] ^ uncoded_block[213];
  wire _2541 = _2540 ^ _101;
  wire _2542 = _2539 ^ _2541;
  wire _2543 = uncoded_block[218] ^ uncoded_block[220];
  wire _2544 = _2543 ^ _104;
  wire _2545 = uncoded_block[224] ^ uncoded_block[225];
  wire _2546 = _2545 ^ _109;
  wire _2547 = _2544 ^ _2546;
  wire _2548 = _2542 ^ _2547;
  wire _2549 = uncoded_block[230] ^ uncoded_block[232];
  wire _2550 = uncoded_block[233] ^ uncoded_block[234];
  wire _2551 = _2549 ^ _2550;
  wire _2552 = uncoded_block[238] ^ uncoded_block[239];
  wire _2553 = uncoded_block[241] ^ uncoded_block[245];
  wire _2554 = _2552 ^ _2553;
  wire _2555 = _2551 ^ _2554;
  wire _2556 = uncoded_block[248] ^ uncoded_block[250];
  wire _2557 = uncoded_block[251] ^ uncoded_block[253];
  wire _2558 = _2556 ^ _2557;
  wire _2559 = uncoded_block[255] ^ uncoded_block[258];
  wire _2560 = _2559 ^ _119;
  wire _2561 = _2558 ^ _2560;
  wire _2562 = _2555 ^ _2561;
  wire _2563 = _2548 ^ _2562;
  wire _2564 = _2536 ^ _2563;
  wire _2565 = _2509 ^ _2564;
  wire _2566 = uncoded_block[270] ^ uncoded_block[271];
  wire _2567 = _1789 ^ _2566;
  wire _2568 = uncoded_block[274] ^ uncoded_block[277];
  wire _2569 = _2568 ^ _988;
  wire _2570 = _2567 ^ _2569;
  wire _2571 = uncoded_block[290] ^ uncoded_block[292];
  wire _2572 = _991 ^ _2571;
  wire _2573 = uncoded_block[293] ^ uncoded_block[295];
  wire _2574 = _2573 ^ _1806;
  wire _2575 = _2572 ^ _2574;
  wire _2576 = _2570 ^ _2575;
  wire _2577 = uncoded_block[298] ^ uncoded_block[300];
  wire _2578 = uncoded_block[306] ^ uncoded_block[312];
  wire _2579 = _2577 ^ _2578;
  wire _2580 = uncoded_block[318] ^ uncoded_block[321];
  wire _2581 = _146 ^ _2580;
  wire _2582 = _2579 ^ _2581;
  wire _2583 = uncoded_block[323] ^ uncoded_block[326];
  wire _2584 = uncoded_block[328] ^ uncoded_block[329];
  wire _2585 = _2583 ^ _2584;
  wire _2586 = uncoded_block[330] ^ uncoded_block[331];
  wire _2587 = uncoded_block[332] ^ uncoded_block[334];
  wire _2588 = _2586 ^ _2587;
  wire _2589 = _2585 ^ _2588;
  wire _2590 = _2582 ^ _2589;
  wire _2591 = _2576 ^ _2590;
  wire _2592 = uncoded_block[336] ^ uncoded_block[337];
  wire _2593 = uncoded_block[338] ^ uncoded_block[340];
  wire _2594 = _2592 ^ _2593;
  wire _2595 = uncoded_block[341] ^ uncoded_block[343];
  wire _2596 = uncoded_block[345] ^ uncoded_block[348];
  wire _2597 = _2595 ^ _2596;
  wire _2598 = _2594 ^ _2597;
  wire _2599 = uncoded_block[349] ^ uncoded_block[351];
  wire _2600 = _2599 ^ _162;
  wire _2601 = uncoded_block[354] ^ uncoded_block[355];
  wire _2602 = uncoded_block[356] ^ uncoded_block[357];
  wire _2603 = _2601 ^ _2602;
  wire _2604 = _2600 ^ _2603;
  wire _2605 = _2598 ^ _2604;
  wire _2606 = uncoded_block[359] ^ uncoded_block[360];
  wire _2607 = _2606 ^ _1031;
  wire _2608 = uncoded_block[364] ^ uncoded_block[371];
  wire _2609 = uncoded_block[378] ^ uncoded_block[380];
  wire _2610 = _2608 ^ _2609;
  wire _2611 = _2607 ^ _2610;
  wire _2612 = uncoded_block[381] ^ uncoded_block[383];
  wire _2613 = uncoded_block[387] ^ uncoded_block[388];
  wire _2614 = _2612 ^ _2613;
  wire _2615 = uncoded_block[390] ^ uncoded_block[391];
  wire _2616 = uncoded_block[392] ^ uncoded_block[396];
  wire _2617 = _2615 ^ _2616;
  wire _2618 = _2614 ^ _2617;
  wire _2619 = _2611 ^ _2618;
  wire _2620 = _2605 ^ _2619;
  wire _2621 = _2591 ^ _2620;
  wire _2622 = uncoded_block[397] ^ uncoded_block[398];
  wire _2623 = uncoded_block[399] ^ uncoded_block[400];
  wire _2624 = _2622 ^ _2623;
  wire _2625 = uncoded_block[402] ^ uncoded_block[403];
  wire _2626 = uncoded_block[404] ^ uncoded_block[408];
  wire _2627 = _2625 ^ _2626;
  wire _2628 = _2624 ^ _2627;
  wire _2629 = uncoded_block[409] ^ uncoded_block[410];
  wire _2630 = uncoded_block[412] ^ uncoded_block[414];
  wire _2631 = _2629 ^ _2630;
  wire _2632 = uncoded_block[418] ^ uncoded_block[423];
  wire _2633 = uncoded_block[424] ^ uncoded_block[425];
  wire _2634 = _2632 ^ _2633;
  wire _2635 = _2631 ^ _2634;
  wire _2636 = _2628 ^ _2635;
  wire _2637 = uncoded_block[426] ^ uncoded_block[428];
  wire _2638 = uncoded_block[431] ^ uncoded_block[432];
  wire _2639 = _2637 ^ _2638;
  wire _2640 = uncoded_block[434] ^ uncoded_block[435];
  wire _2641 = uncoded_block[438] ^ uncoded_block[440];
  wire _2642 = _2640 ^ _2641;
  wire _2643 = _2639 ^ _2642;
  wire _2644 = uncoded_block[445] ^ uncoded_block[450];
  wire _2645 = uncoded_block[452] ^ uncoded_block[453];
  wire _2646 = _2644 ^ _2645;
  wire _2647 = _207 ^ _2646;
  wire _2648 = _2643 ^ _2647;
  wire _2649 = _2636 ^ _2648;
  wire _2650 = uncoded_block[454] ^ uncoded_block[455];
  wire _2651 = uncoded_block[456] ^ uncoded_block[459];
  wire _2652 = _2650 ^ _2651;
  wire _2653 = uncoded_block[460] ^ uncoded_block[461];
  wire _2654 = uncoded_block[464] ^ uncoded_block[467];
  wire _2655 = _2653 ^ _2654;
  wire _2656 = _2652 ^ _2655;
  wire _2657 = uncoded_block[475] ^ uncoded_block[476];
  wire _2658 = _2657 ^ _1085;
  wire _2659 = uncoded_block[481] ^ uncoded_block[484];
  wire _2660 = uncoded_block[485] ^ uncoded_block[487];
  wire _2661 = _2659 ^ _2660;
  wire _2662 = _2658 ^ _2661;
  wire _2663 = _2656 ^ _2662;
  wire _2664 = uncoded_block[491] ^ uncoded_block[492];
  wire _2665 = uncoded_block[493] ^ uncoded_block[496];
  wire _2666 = _2664 ^ _2665;
  wire _2667 = uncoded_block[497] ^ uncoded_block[499];
  wire _2668 = uncoded_block[502] ^ uncoded_block[503];
  wire _2669 = _2667 ^ _2668;
  wire _2670 = _2666 ^ _2669;
  wire _2671 = uncoded_block[504] ^ uncoded_block[505];
  wire _2672 = _2671 ^ _1892;
  wire _2673 = uncoded_block[508] ^ uncoded_block[513];
  wire _2674 = _2673 ^ _232;
  wire _2675 = _2672 ^ _2674;
  wire _2676 = _2670 ^ _2675;
  wire _2677 = _2663 ^ _2676;
  wire _2678 = _2649 ^ _2677;
  wire _2679 = _2621 ^ _2678;
  wire _2680 = _2565 ^ _2679;
  wire _2681 = uncoded_block[518] ^ uncoded_block[523];
  wire _2682 = _2681 ^ _239;
  wire _2683 = uncoded_block[531] ^ uncoded_block[536];
  wire _2684 = uncoded_block[542] ^ uncoded_block[545];
  wire _2685 = _2683 ^ _2684;
  wire _2686 = _2682 ^ _2685;
  wire _2687 = uncoded_block[548] ^ uncoded_block[550];
  wire _2688 = uncoded_block[551] ^ uncoded_block[552];
  wire _2689 = _2687 ^ _2688;
  wire _2690 = uncoded_block[560] ^ uncoded_block[565];
  wire _2691 = _1915 ^ _2690;
  wire _2692 = _2689 ^ _2691;
  wire _2693 = _2686 ^ _2692;
  wire _2694 = _1129 ^ _262;
  wire _2695 = uncoded_block[575] ^ uncoded_block[581];
  wire _2696 = uncoded_block[582] ^ uncoded_block[584];
  wire _2697 = _2695 ^ _2696;
  wire _2698 = _2694 ^ _2697;
  wire _2699 = _1139 ^ _1141;
  wire _2700 = uncoded_block[591] ^ uncoded_block[592];
  wire _2701 = uncoded_block[594] ^ uncoded_block[596];
  wire _2702 = _2700 ^ _2701;
  wire _2703 = _2699 ^ _2702;
  wire _2704 = _2698 ^ _2703;
  wire _2705 = _2693 ^ _2704;
  wire _2706 = uncoded_block[597] ^ uncoded_block[598];
  wire _2707 = uncoded_block[600] ^ uncoded_block[601];
  wire _2708 = _2706 ^ _2707;
  wire _2709 = uncoded_block[602] ^ uncoded_block[603];
  wire _2710 = uncoded_block[604] ^ uncoded_block[605];
  wire _2711 = _2709 ^ _2710;
  wire _2712 = _2708 ^ _2711;
  wire _2713 = uncoded_block[609] ^ uncoded_block[610];
  wire _2714 = _277 ^ _2713;
  wire _2715 = uncoded_block[611] ^ uncoded_block[616];
  wire _2716 = _2715 ^ _281;
  wire _2717 = _2714 ^ _2716;
  wire _2718 = _2712 ^ _2717;
  wire _2719 = uncoded_block[621] ^ uncoded_block[624];
  wire _2720 = uncoded_block[625] ^ uncoded_block[627];
  wire _2721 = _2719 ^ _2720;
  wire _2722 = uncoded_block[628] ^ uncoded_block[631];
  wire _2723 = uncoded_block[632] ^ uncoded_block[636];
  wire _2724 = _2722 ^ _2723;
  wire _2725 = _2721 ^ _2724;
  wire _2726 = uncoded_block[637] ^ uncoded_block[640];
  wire _2727 = uncoded_block[641] ^ uncoded_block[642];
  wire _2728 = _2726 ^ _2727;
  wire _2729 = uncoded_block[644] ^ uncoded_block[645];
  wire _2730 = uncoded_block[647] ^ uncoded_block[648];
  wire _2731 = _2729 ^ _2730;
  wire _2732 = _2728 ^ _2731;
  wire _2733 = _2725 ^ _2732;
  wire _2734 = _2718 ^ _2733;
  wire _2735 = _2705 ^ _2734;
  wire _2736 = uncoded_block[653] ^ uncoded_block[656];
  wire _2737 = _1960 ^ _2736;
  wire _2738 = uncoded_block[657] ^ uncoded_block[658];
  wire _2739 = uncoded_block[660] ^ uncoded_block[661];
  wire _2740 = _2738 ^ _2739;
  wire _2741 = _2737 ^ _2740;
  wire _2742 = uncoded_block[662] ^ uncoded_block[665];
  wire _2743 = _2742 ^ _309;
  wire _2744 = uncoded_block[670] ^ uncoded_block[672];
  wire _2745 = _1174 ^ _2744;
  wire _2746 = _2743 ^ _2745;
  wire _2747 = _2741 ^ _2746;
  wire _2748 = uncoded_block[674] ^ uncoded_block[675];
  wire _2749 = _2748 ^ _1181;
  wire _2750 = uncoded_block[683] ^ uncoded_block[686];
  wire _2751 = uncoded_block[688] ^ uncoded_block[689];
  wire _2752 = _2750 ^ _2751;
  wire _2753 = _2749 ^ _2752;
  wire _2754 = uncoded_block[690] ^ uncoded_block[691];
  wire _2755 = uncoded_block[692] ^ uncoded_block[694];
  wire _2756 = _2754 ^ _2755;
  wire _2757 = uncoded_block[695] ^ uncoded_block[700];
  wire _2758 = _2757 ^ _334;
  wire _2759 = _2756 ^ _2758;
  wire _2760 = _2753 ^ _2759;
  wire _2761 = _2747 ^ _2760;
  wire _2762 = uncoded_block[711] ^ uncoded_block[712];
  wire _2763 = uncoded_block[715] ^ uncoded_block[718];
  wire _2764 = _2762 ^ _2763;
  wire _2765 = uncoded_block[720] ^ uncoded_block[724];
  wire _2766 = _2765 ^ _1988;
  wire _2767 = _2764 ^ _2766;
  wire _2768 = uncoded_block[729] ^ uncoded_block[730];
  wire _2769 = _2768 ^ _1991;
  wire _2770 = uncoded_block[738] ^ uncoded_block[740];
  wire _2771 = _1995 ^ _2770;
  wire _2772 = _2769 ^ _2771;
  wire _2773 = _2767 ^ _2772;
  wire _2774 = uncoded_block[741] ^ uncoded_block[744];
  wire _2775 = uncoded_block[745] ^ uncoded_block[747];
  wire _2776 = _2774 ^ _2775;
  wire _2777 = uncoded_block[749] ^ uncoded_block[751];
  wire _2778 = uncoded_block[755] ^ uncoded_block[756];
  wire _2779 = _2777 ^ _2778;
  wire _2780 = _2776 ^ _2779;
  wire _2781 = uncoded_block[762] ^ uncoded_block[763];
  wire _2782 = _2005 ^ _2781;
  wire _2783 = uncoded_block[764] ^ uncoded_block[765];
  wire _2784 = uncoded_block[766] ^ uncoded_block[769];
  wire _2785 = _2783 ^ _2784;
  wire _2786 = _2782 ^ _2785;
  wire _2787 = _2780 ^ _2786;
  wire _2788 = _2773 ^ _2787;
  wire _2789 = _2761 ^ _2788;
  wire _2790 = _2735 ^ _2789;
  wire _2791 = uncoded_block[770] ^ uncoded_block[773];
  wire _2792 = uncoded_block[774] ^ uncoded_block[776];
  wire _2793 = _2791 ^ _2792;
  wire _2794 = uncoded_block[781] ^ uncoded_block[782];
  wire _2795 = uncoded_block[783] ^ uncoded_block[787];
  wire _2796 = _2794 ^ _2795;
  wire _2797 = _2793 ^ _2796;
  wire _2798 = uncoded_block[788] ^ uncoded_block[791];
  wire _2799 = uncoded_block[793] ^ uncoded_block[794];
  wire _2800 = _2798 ^ _2799;
  wire _2801 = uncoded_block[799] ^ uncoded_block[801];
  wire _2802 = _382 ^ _2801;
  wire _2803 = _2800 ^ _2802;
  wire _2804 = _2797 ^ _2803;
  wire _2805 = uncoded_block[803] ^ uncoded_block[811];
  wire _2806 = uncoded_block[812] ^ uncoded_block[814];
  wire _2807 = _2805 ^ _2806;
  wire _2808 = uncoded_block[815] ^ uncoded_block[816];
  wire _2809 = uncoded_block[819] ^ uncoded_block[823];
  wire _2810 = _2808 ^ _2809;
  wire _2811 = _2807 ^ _2810;
  wire _2812 = uncoded_block[828] ^ uncoded_block[829];
  wire _2813 = _2812 ^ _400;
  wire _2814 = uncoded_block[836] ^ uncoded_block[838];
  wire _2815 = uncoded_block[840] ^ uncoded_block[843];
  wire _2816 = _2814 ^ _2815;
  wire _2817 = _2813 ^ _2816;
  wire _2818 = _2811 ^ _2817;
  wire _2819 = _2804 ^ _2818;
  wire _2820 = uncoded_block[846] ^ uncoded_block[848];
  wire _2821 = uncoded_block[852] ^ uncoded_block[853];
  wire _2822 = _2820 ^ _2821;
  wire _2823 = uncoded_block[854] ^ uncoded_block[859];
  wire _2824 = uncoded_block[861] ^ uncoded_block[863];
  wire _2825 = _2823 ^ _2824;
  wire _2826 = _2822 ^ _2825;
  wire _2827 = uncoded_block[865] ^ uncoded_block[867];
  wire _2828 = uncoded_block[868] ^ uncoded_block[869];
  wire _2829 = _2827 ^ _2828;
  wire _2830 = uncoded_block[870] ^ uncoded_block[873];
  wire _2831 = uncoded_block[874] ^ uncoded_block[876];
  wire _2832 = _2830 ^ _2831;
  wire _2833 = _2829 ^ _2832;
  wire _2834 = _2826 ^ _2833;
  wire _2835 = uncoded_block[878] ^ uncoded_block[879];
  wire _2836 = uncoded_block[881] ^ uncoded_block[882];
  wire _2837 = _2835 ^ _2836;
  wire _2838 = uncoded_block[883] ^ uncoded_block[884];
  wire _2839 = _2838 ^ _2058;
  wire _2840 = _2837 ^ _2839;
  wire _2841 = uncoded_block[893] ^ uncoded_block[898];
  wire _2842 = _1273 ^ _2841;
  wire _2843 = uncoded_block[899] ^ uncoded_block[900];
  wire _2844 = uncoded_block[901] ^ uncoded_block[902];
  wire _2845 = _2843 ^ _2844;
  wire _2846 = _2842 ^ _2845;
  wire _2847 = _2840 ^ _2846;
  wire _2848 = _2834 ^ _2847;
  wire _2849 = _2819 ^ _2848;
  wire _2850 = uncoded_block[904] ^ uncoded_block[907];
  wire _2851 = _2850 ^ _2071;
  wire _2852 = uncoded_block[916] ^ uncoded_block[917];
  wire _2853 = _1287 ^ _2852;
  wire _2854 = _2851 ^ _2853;
  wire _2855 = uncoded_block[924] ^ uncoded_block[926];
  wire _2856 = _445 ^ _2855;
  wire _2857 = uncoded_block[927] ^ uncoded_block[929];
  wire _2858 = uncoded_block[930] ^ uncoded_block[932];
  wire _2859 = _2857 ^ _2858;
  wire _2860 = _2856 ^ _2859;
  wire _2861 = _2854 ^ _2860;
  wire _2862 = uncoded_block[935] ^ uncoded_block[936];
  wire _2863 = uncoded_block[940] ^ uncoded_block[942];
  wire _2864 = _2862 ^ _2863;
  wire _2865 = uncoded_block[943] ^ uncoded_block[944];
  wire _2866 = uncoded_block[946] ^ uncoded_block[952];
  wire _2867 = _2865 ^ _2866;
  wire _2868 = _2864 ^ _2867;
  wire _2869 = uncoded_block[954] ^ uncoded_block[956];
  wire _2870 = _2869 ^ _2090;
  wire _2871 = uncoded_block[959] ^ uncoded_block[961];
  wire _2872 = uncoded_block[962] ^ uncoded_block[964];
  wire _2873 = _2871 ^ _2872;
  wire _2874 = _2870 ^ _2873;
  wire _2875 = _2868 ^ _2874;
  wire _2876 = _2861 ^ _2875;
  wire _2877 = uncoded_block[972] ^ uncoded_block[973];
  wire _2878 = _1311 ^ _2877;
  wire _2879 = uncoded_block[981] ^ uncoded_block[987];
  wire _2880 = _2100 ^ _2879;
  wire _2881 = _2878 ^ _2880;
  wire _2882 = uncoded_block[990] ^ uncoded_block[991];
  wire _2883 = uncoded_block[994] ^ uncoded_block[996];
  wire _2884 = _2882 ^ _2883;
  wire _2885 = uncoded_block[997] ^ uncoded_block[1003];
  wire _2886 = uncoded_block[1006] ^ uncoded_block[1007];
  wire _2887 = _2885 ^ _2886;
  wire _2888 = _2884 ^ _2887;
  wire _2889 = _2881 ^ _2888;
  wire _2890 = uncoded_block[1010] ^ uncoded_block[1013];
  wire _2891 = uncoded_block[1014] ^ uncoded_block[1016];
  wire _2892 = _2890 ^ _2891;
  wire _2893 = uncoded_block[1017] ^ uncoded_block[1018];
  wire _2894 = uncoded_block[1019] ^ uncoded_block[1020];
  wire _2895 = _2893 ^ _2894;
  wire _2896 = _2892 ^ _2895;
  wire _2897 = _1338 ^ _495;
  wire _2898 = uncoded_block[1029] ^ uncoded_block[1030];
  wire _2899 = _498 ^ _2898;
  wire _2900 = _2897 ^ _2899;
  wire _2901 = _2896 ^ _2900;
  wire _2902 = _2889 ^ _2901;
  wire _2903 = _2876 ^ _2902;
  wire _2904 = _2849 ^ _2903;
  wire _2905 = _2790 ^ _2904;
  wire _2906 = _2680 ^ _2905;
  wire _2907 = uncoded_block[1031] ^ uncoded_block[1033];
  wire _2908 = uncoded_block[1035] ^ uncoded_block[1037];
  wire _2909 = _2907 ^ _2908;
  wire _2910 = uncoded_block[1043] ^ uncoded_block[1045];
  wire _2911 = _511 ^ _2910;
  wire _2912 = _2909 ^ _2911;
  wire _2913 = uncoded_block[1046] ^ uncoded_block[1050];
  wire _2914 = uncoded_block[1051] ^ uncoded_block[1054];
  wire _2915 = _2913 ^ _2914;
  wire _2916 = uncoded_block[1058] ^ uncoded_block[1061];
  wire _2917 = uncoded_block[1062] ^ uncoded_block[1064];
  wire _2918 = _2916 ^ _2917;
  wire _2919 = _2915 ^ _2918;
  wire _2920 = _2912 ^ _2919;
  wire _2921 = uncoded_block[1065] ^ uncoded_block[1066];
  wire _2922 = uncoded_block[1068] ^ uncoded_block[1073];
  wire _2923 = _2921 ^ _2922;
  wire _2924 = uncoded_block[1075] ^ uncoded_block[1076];
  wire _2925 = uncoded_block[1077] ^ uncoded_block[1080];
  wire _2926 = _2924 ^ _2925;
  wire _2927 = _2923 ^ _2926;
  wire _2928 = uncoded_block[1084] ^ uncoded_block[1085];
  wire _2929 = _2928 ^ _2149;
  wire _2930 = uncoded_block[1090] ^ uncoded_block[1093];
  wire _2931 = _2930 ^ _542;
  wire _2932 = _2929 ^ _2931;
  wire _2933 = _2927 ^ _2932;
  wire _2934 = _2920 ^ _2933;
  wire _2935 = uncoded_block[1097] ^ uncoded_block[1100];
  wire _2936 = _2935 ^ _2160;
  wire _2937 = uncoded_block[1107] ^ uncoded_block[1112];
  wire _2938 = uncoded_block[1114] ^ uncoded_block[1116];
  wire _2939 = _2937 ^ _2938;
  wire _2940 = _2936 ^ _2939;
  wire _2941 = uncoded_block[1119] ^ uncoded_block[1121];
  wire _2942 = uncoded_block[1122] ^ uncoded_block[1123];
  wire _2943 = _2941 ^ _2942;
  wire _2944 = uncoded_block[1124] ^ uncoded_block[1125];
  wire _2945 = uncoded_block[1127] ^ uncoded_block[1130];
  wire _2946 = _2944 ^ _2945;
  wire _2947 = _2943 ^ _2946;
  wire _2948 = _2940 ^ _2947;
  wire _2949 = uncoded_block[1132] ^ uncoded_block[1134];
  wire _2950 = uncoded_block[1135] ^ uncoded_block[1139];
  wire _2951 = _2949 ^ _2950;
  wire _2952 = uncoded_block[1141] ^ uncoded_block[1143];
  wire _2953 = uncoded_block[1144] ^ uncoded_block[1145];
  wire _2954 = _2952 ^ _2953;
  wire _2955 = _2951 ^ _2954;
  wire _2956 = uncoded_block[1149] ^ uncoded_block[1150];
  wire _2957 = _2956 ^ _577;
  wire _2958 = uncoded_block[1161] ^ uncoded_block[1162];
  wire _2959 = _1404 ^ _2958;
  wire _2960 = _2957 ^ _2959;
  wire _2961 = _2955 ^ _2960;
  wire _2962 = _2948 ^ _2961;
  wire _2963 = _2934 ^ _2962;
  wire _2964 = uncoded_block[1163] ^ uncoded_block[1164];
  wire _2965 = uncoded_block[1168] ^ uncoded_block[1173];
  wire _2966 = _2964 ^ _2965;
  wire _2967 = uncoded_block[1174] ^ uncoded_block[1175];
  wire _2968 = _2967 ^ _589;
  wire _2969 = _2966 ^ _2968;
  wire _2970 = uncoded_block[1180] ^ uncoded_block[1187];
  wire _2971 = uncoded_block[1190] ^ uncoded_block[1191];
  wire _2972 = _2970 ^ _2971;
  wire _2973 = uncoded_block[1196] ^ uncoded_block[1201];
  wire _2974 = uncoded_block[1202] ^ uncoded_block[1203];
  wire _2975 = _2973 ^ _2974;
  wire _2976 = _2972 ^ _2975;
  wire _2977 = _2969 ^ _2976;
  wire _2978 = uncoded_block[1204] ^ uncoded_block[1205];
  wire _2979 = uncoded_block[1206] ^ uncoded_block[1209];
  wire _2980 = _2978 ^ _2979;
  wire _2981 = uncoded_block[1210] ^ uncoded_block[1213];
  wire _2982 = uncoded_block[1214] ^ uncoded_block[1215];
  wire _2983 = _2981 ^ _2982;
  wire _2984 = _2980 ^ _2983;
  wire _2985 = uncoded_block[1219] ^ uncoded_block[1223];
  wire _2986 = uncoded_block[1225] ^ uncoded_block[1227];
  wire _2987 = _2985 ^ _2986;
  wire _2988 = uncoded_block[1232] ^ uncoded_block[1235];
  wire _2989 = uncoded_block[1236] ^ uncoded_block[1237];
  wire _2990 = _2988 ^ _2989;
  wire _2991 = _2987 ^ _2990;
  wire _2992 = _2984 ^ _2991;
  wire _2993 = _2977 ^ _2992;
  wire _2994 = uncoded_block[1239] ^ uncoded_block[1242];
  wire _2995 = uncoded_block[1243] ^ uncoded_block[1244];
  wire _2996 = _2994 ^ _2995;
  wire _2997 = uncoded_block[1246] ^ uncoded_block[1248];
  wire _2998 = uncoded_block[1249] ^ uncoded_block[1252];
  wire _2999 = _2997 ^ _2998;
  wire _3000 = _2996 ^ _2999;
  wire _3001 = uncoded_block[1255] ^ uncoded_block[1256];
  wire _3002 = _3001 ^ _624;
  wire _3003 = uncoded_block[1261] ^ uncoded_block[1262];
  wire _3004 = uncoded_block[1263] ^ uncoded_block[1264];
  wire _3005 = _3003 ^ _3004;
  wire _3006 = _3002 ^ _3005;
  wire _3007 = _3000 ^ _3006;
  wire _3008 = uncoded_block[1267] ^ uncoded_block[1268];
  wire _3009 = _3008 ^ _1459;
  wire _3010 = uncoded_block[1271] ^ uncoded_block[1275];
  wire _3011 = uncoded_block[1279] ^ uncoded_block[1282];
  wire _3012 = _3010 ^ _3011;
  wire _3013 = _3009 ^ _3012;
  wire _3014 = uncoded_block[1283] ^ uncoded_block[1294];
  wire _3015 = uncoded_block[1295] ^ uncoded_block[1296];
  wire _3016 = _3014 ^ _3015;
  wire _3017 = uncoded_block[1297] ^ uncoded_block[1298];
  wire _3018 = uncoded_block[1300] ^ uncoded_block[1303];
  wire _3019 = _3017 ^ _3018;
  wire _3020 = _3016 ^ _3019;
  wire _3021 = _3013 ^ _3020;
  wire _3022 = _3007 ^ _3021;
  wire _3023 = _2993 ^ _3022;
  wire _3024 = _2963 ^ _3023;
  wire _3025 = uncoded_block[1305] ^ uncoded_block[1308];
  wire _3026 = uncoded_block[1313] ^ uncoded_block[1316];
  wire _3027 = _3025 ^ _3026;
  wire _3028 = uncoded_block[1319] ^ uncoded_block[1320];
  wire _3029 = uncoded_block[1321] ^ uncoded_block[1322];
  wire _3030 = _3028 ^ _3029;
  wire _3031 = _3027 ^ _3030;
  wire _3032 = uncoded_block[1324] ^ uncoded_block[1326];
  wire _3033 = _3032 ^ _1490;
  wire _3034 = uncoded_block[1335] ^ uncoded_block[1336];
  wire _3035 = _660 ^ _3034;
  wire _3036 = _3033 ^ _3035;
  wire _3037 = _3031 ^ _3036;
  wire _3038 = uncoded_block[1338] ^ uncoded_block[1344];
  wire _3039 = uncoded_block[1345] ^ uncoded_block[1347];
  wire _3040 = _3038 ^ _3039;
  wire _3041 = uncoded_block[1350] ^ uncoded_block[1351];
  wire _3042 = uncoded_block[1352] ^ uncoded_block[1353];
  wire _3043 = _3041 ^ _3042;
  wire _3044 = _3040 ^ _3043;
  wire _3045 = uncoded_block[1360] ^ uncoded_block[1361];
  wire _3046 = _2280 ^ _3045;
  wire _3047 = uncoded_block[1366] ^ uncoded_block[1368];
  wire _3048 = _2283 ^ _3047;
  wire _3049 = _3046 ^ _3048;
  wire _3050 = _3044 ^ _3049;
  wire _3051 = _3037 ^ _3050;
  wire _3052 = uncoded_block[1369] ^ uncoded_block[1370];
  wire _3053 = _3052 ^ _684;
  wire _3054 = uncoded_block[1374] ^ uncoded_block[1376];
  wire _3055 = uncoded_block[1377] ^ uncoded_block[1378];
  wire _3056 = _3054 ^ _3055;
  wire _3057 = _3053 ^ _3056;
  wire _3058 = uncoded_block[1379] ^ uncoded_block[1380];
  wire _3059 = uncoded_block[1382] ^ uncoded_block[1383];
  wire _3060 = _3058 ^ _3059;
  wire _3061 = uncoded_block[1384] ^ uncoded_block[1385];
  wire _3062 = _3061 ^ _692;
  wire _3063 = _3060 ^ _3062;
  wire _3064 = _3057 ^ _3063;
  wire _3065 = uncoded_block[1395] ^ uncoded_block[1397];
  wire _3066 = uncoded_block[1399] ^ uncoded_block[1400];
  wire _3067 = _3065 ^ _3066;
  wire _3068 = uncoded_block[1403] ^ uncoded_block[1406];
  wire _3069 = uncoded_block[1411] ^ uncoded_block[1415];
  wire _3070 = _3068 ^ _3069;
  wire _3071 = _3067 ^ _3070;
  wire _3072 = uncoded_block[1418] ^ uncoded_block[1422];
  wire _3073 = _2306 ^ _3072;
  wire _3074 = uncoded_block[1423] ^ uncoded_block[1424];
  wire _3075 = uncoded_block[1426] ^ uncoded_block[1429];
  wire _3076 = _3074 ^ _3075;
  wire _3077 = _3073 ^ _3076;
  wire _3078 = _3071 ^ _3077;
  wire _3079 = _3064 ^ _3078;
  wire _3080 = _3051 ^ _3079;
  wire _3081 = uncoded_block[1431] ^ uncoded_block[1433];
  wire _3082 = _3081 ^ _1534;
  wire _3083 = uncoded_block[1438] ^ uncoded_block[1441];
  wire _3084 = uncoded_block[1445] ^ uncoded_block[1446];
  wire _3085 = _3083 ^ _3084;
  wire _3086 = _3082 ^ _3085;
  wire _3087 = _2325 ^ _719;
  wire _3088 = uncoded_block[1456] ^ uncoded_block[1457];
  wire _3089 = uncoded_block[1458] ^ uncoded_block[1459];
  wire _3090 = _3088 ^ _3089;
  wire _3091 = _3087 ^ _3090;
  wire _3092 = _3086 ^ _3091;
  wire _3093 = uncoded_block[1460] ^ uncoded_block[1462];
  wire _3094 = uncoded_block[1464] ^ uncoded_block[1465];
  wire _3095 = _3093 ^ _3094;
  wire _3096 = uncoded_block[1466] ^ uncoded_block[1468];
  wire _3097 = uncoded_block[1472] ^ uncoded_block[1473];
  wire _3098 = _3096 ^ _3097;
  wire _3099 = _3095 ^ _3098;
  wire _3100 = uncoded_block[1477] ^ uncoded_block[1481];
  wire _3101 = uncoded_block[1483] ^ uncoded_block[1485];
  wire _3102 = _3100 ^ _3101;
  wire _3103 = uncoded_block[1490] ^ uncoded_block[1491];
  wire _3104 = _2349 ^ _3103;
  wire _3105 = _3102 ^ _3104;
  wire _3106 = _3099 ^ _3105;
  wire _3107 = _3092 ^ _3106;
  wire _3108 = uncoded_block[1492] ^ uncoded_block[1496];
  wire _3109 = uncoded_block[1498] ^ uncoded_block[1500];
  wire _3110 = _3108 ^ _3109;
  wire _3111 = uncoded_block[1501] ^ uncoded_block[1503];
  wire _3112 = uncoded_block[1506] ^ uncoded_block[1507];
  wire _3113 = _3111 ^ _3112;
  wire _3114 = _3110 ^ _3113;
  wire _3115 = uncoded_block[1513] ^ uncoded_block[1514];
  wire _3116 = _750 ^ _3115;
  wire _3117 = uncoded_block[1515] ^ uncoded_block[1519];
  wire _3118 = uncoded_block[1523] ^ uncoded_block[1524];
  wire _3119 = _3117 ^ _3118;
  wire _3120 = _3116 ^ _3119;
  wire _3121 = _3114 ^ _3120;
  wire _3122 = uncoded_block[1525] ^ uncoded_block[1526];
  wire _3123 = uncoded_block[1527] ^ uncoded_block[1529];
  wire _3124 = _3122 ^ _3123;
  wire _3125 = uncoded_block[1531] ^ uncoded_block[1534];
  wire _3126 = _3125 ^ _1587;
  wire _3127 = _3124 ^ _3126;
  wire _3128 = uncoded_block[1540] ^ uncoded_block[1542];
  wire _3129 = uncoded_block[1543] ^ uncoded_block[1545];
  wire _3130 = _3128 ^ _3129;
  wire _3131 = uncoded_block[1554] ^ uncoded_block[1556];
  wire _3132 = _2367 ^ _3131;
  wire _3133 = _3130 ^ _3132;
  wire _3134 = _3127 ^ _3133;
  wire _3135 = _3121 ^ _3134;
  wire _3136 = _3107 ^ _3135;
  wire _3137 = _3080 ^ _3136;
  wire _3138 = _3024 ^ _3137;
  wire _3139 = uncoded_block[1560] ^ uncoded_block[1563];
  wire _3140 = _3139 ^ _2376;
  wire _3141 = uncoded_block[1567] ^ uncoded_block[1572];
  wire _3142 = _3141 ^ _781;
  wire _3143 = _3140 ^ _3142;
  wire _3144 = _1613 ^ _1615;
  wire _3145 = uncoded_block[1588] ^ uncoded_block[1590];
  wire _3146 = uncoded_block[1591] ^ uncoded_block[1592];
  wire _3147 = _3145 ^ _3146;
  wire _3148 = _3144 ^ _3147;
  wire _3149 = _3143 ^ _3148;
  wire _3150 = uncoded_block[1595] ^ uncoded_block[1600];
  wire _3151 = uncoded_block[1601] ^ uncoded_block[1602];
  wire _3152 = _3150 ^ _3151;
  wire _3153 = uncoded_block[1604] ^ uncoded_block[1605];
  wire _3154 = uncoded_block[1608] ^ uncoded_block[1610];
  wire _3155 = _3153 ^ _3154;
  wire _3156 = _3152 ^ _3155;
  wire _3157 = uncoded_block[1611] ^ uncoded_block[1613];
  wire _3158 = uncoded_block[1614] ^ uncoded_block[1619];
  wire _3159 = _3157 ^ _3158;
  wire _3160 = uncoded_block[1620] ^ uncoded_block[1622];
  wire _3161 = uncoded_block[1627] ^ uncoded_block[1629];
  wire _3162 = _3160 ^ _3161;
  wire _3163 = _3159 ^ _3162;
  wire _3164 = _3156 ^ _3163;
  wire _3165 = _3149 ^ _3164;
  wire _3166 = uncoded_block[1630] ^ uncoded_block[1632];
  wire _3167 = uncoded_block[1635] ^ uncoded_block[1640];
  wire _3168 = _3166 ^ _3167;
  wire _3169 = uncoded_block[1643] ^ uncoded_block[1644];
  wire _3170 = _2408 ^ _3169;
  wire _3171 = _3168 ^ _3170;
  wire _3172 = uncoded_block[1650] ^ uncoded_block[1651];
  wire _3173 = _816 ^ _3172;
  wire _3174 = uncoded_block[1657] ^ uncoded_block[1658];
  wire _3175 = uncoded_block[1661] ^ uncoded_block[1663];
  wire _3176 = _3174 ^ _3175;
  wire _3177 = _3173 ^ _3176;
  wire _3178 = _3171 ^ _3177;
  wire _3179 = uncoded_block[1664] ^ uncoded_block[1665];
  wire _3180 = uncoded_block[1666] ^ uncoded_block[1669];
  wire _3181 = _3179 ^ _3180;
  wire _3182 = uncoded_block[1670] ^ uncoded_block[1671];
  wire _3183 = uncoded_block[1675] ^ uncoded_block[1676];
  wire _3184 = _3182 ^ _3183;
  wire _3185 = _3181 ^ _3184;
  wire _3186 = uncoded_block[1678] ^ uncoded_block[1680];
  wire _3187 = uncoded_block[1684] ^ uncoded_block[1685];
  wire _3188 = _3186 ^ _3187;
  wire _3189 = uncoded_block[1687] ^ uncoded_block[1688];
  wire _3190 = uncoded_block[1689] ^ uncoded_block[1692];
  wire _3191 = _3189 ^ _3190;
  wire _3192 = _3188 ^ _3191;
  wire _3193 = _3185 ^ _3192;
  wire _3194 = _3178 ^ _3193;
  wire _3195 = _3165 ^ _3194;
  wire _3196 = uncoded_block[1702] ^ uncoded_block[1706];
  wire _3197 = _840 ^ _3196;
  wire _3198 = _848 ^ _2438;
  wire _3199 = _3197 ^ _3198;
  wire _3200 = uncoded_block[1713] ^ uncoded_block[1714];
  wire _3201 = _3200 ^ _2441;
  wire _3202 = _2443 ^ _860;
  wire _3203 = _3201 ^ _3202;
  wire _3204 = _3199 ^ _3203;
  wire _3205 = _3204 ^ uncoded_block[1722];
  wire _3206 = _3195 ^ _3205;
  wire _3207 = _3138 ^ _3206;
  wire _3208 = _2906 ^ _3207;
  wire _3209 = uncoded_block[0] ^ uncoded_block[1];
  wire _3210 = uncoded_block[2] ^ uncoded_block[3];
  wire _3211 = _3209 ^ _3210;
  wire _3212 = uncoded_block[5] ^ uncoded_block[8];
  wire _3213 = uncoded_block[9] ^ uncoded_block[11];
  wire _3214 = _3212 ^ _3213;
  wire _3215 = _3211 ^ _3214;
  wire _3216 = uncoded_block[12] ^ uncoded_block[15];
  wire _3217 = uncoded_block[19] ^ uncoded_block[20];
  wire _3218 = _3216 ^ _3217;
  wire _3219 = uncoded_block[21] ^ uncoded_block[22];
  wire _3220 = uncoded_block[23] ^ uncoded_block[24];
  wire _3221 = _3219 ^ _3220;
  wire _3222 = _3218 ^ _3221;
  wire _3223 = _3215 ^ _3222;
  wire _3224 = uncoded_block[25] ^ uncoded_block[28];
  wire _3225 = uncoded_block[31] ^ uncoded_block[33];
  wire _3226 = _3224 ^ _3225;
  wire _3227 = uncoded_block[34] ^ uncoded_block[36];
  wire _3228 = _3227 ^ _18;
  wire _3229 = _3226 ^ _3228;
  wire _3230 = uncoded_block[40] ^ uncoded_block[41];
  wire _3231 = _3230 ^ _22;
  wire _3232 = uncoded_block[48] ^ uncoded_block[49];
  wire _3233 = uncoded_block[50] ^ uncoded_block[51];
  wire _3234 = _3232 ^ _3233;
  wire _3235 = _3231 ^ _3234;
  wire _3236 = _3229 ^ _3235;
  wire _3237 = _3223 ^ _3236;
  wire _3238 = _1700 ^ _1703;
  wire _3239 = _889 ^ _1706;
  wire _3240 = _3238 ^ _3239;
  wire _3241 = uncoded_block[70] ^ uncoded_block[72];
  wire _3242 = _35 ^ _3241;
  wire _3243 = uncoded_block[76] ^ uncoded_block[79];
  wire _3244 = _3243 ^ _2483;
  wire _3245 = _3242 ^ _3244;
  wire _3246 = _3240 ^ _3245;
  wire _3247 = uncoded_block[88] ^ uncoded_block[93];
  wire _3248 = _2484 ^ _3247;
  wire _3249 = uncoded_block[97] ^ uncoded_block[99];
  wire _3250 = uncoded_block[102] ^ uncoded_block[106];
  wire _3251 = _3249 ^ _3250;
  wire _3252 = _3248 ^ _3251;
  wire _3253 = uncoded_block[113] ^ uncoded_block[115];
  wire _3254 = _1722 ^ _3253;
  wire _3255 = uncoded_block[122] ^ uncoded_block[123];
  wire _3256 = uncoded_block[124] ^ uncoded_block[127];
  wire _3257 = _3255 ^ _3256;
  wire _3258 = _3254 ^ _3257;
  wire _3259 = _3252 ^ _3258;
  wire _3260 = _3246 ^ _3259;
  wire _3261 = _3237 ^ _3260;
  wire _3262 = uncoded_block[128] ^ uncoded_block[129];
  wire _3263 = uncoded_block[134] ^ uncoded_block[136];
  wire _3264 = _3262 ^ _3263;
  wire _3265 = uncoded_block[139] ^ uncoded_block[140];
  wire _3266 = _3265 ^ _2511;
  wire _3267 = _3264 ^ _3266;
  wire _3268 = uncoded_block[149] ^ uncoded_block[151];
  wire _3269 = uncoded_block[152] ^ uncoded_block[153];
  wire _3270 = _3268 ^ _3269;
  wire _3271 = uncoded_block[155] ^ uncoded_block[156];
  wire _3272 = uncoded_block[157] ^ uncoded_block[162];
  wire _3273 = _3271 ^ _3272;
  wire _3274 = _3270 ^ _3273;
  wire _3275 = _3267 ^ _3274;
  wire _3276 = uncoded_block[163] ^ uncoded_block[168];
  wire _3277 = _3276 ^ _81;
  wire _3278 = uncoded_block[174] ^ uncoded_block[175];
  wire _3279 = _3278 ^ _82;
  wire _3280 = _3277 ^ _3279;
  wire _3281 = uncoded_block[179] ^ uncoded_block[184];
  wire _3282 = _3281 ^ _1759;
  wire _3283 = uncoded_block[191] ^ uncoded_block[193];
  wire _3284 = uncoded_block[194] ^ uncoded_block[195];
  wire _3285 = _3283 ^ _3284;
  wire _3286 = _3282 ^ _3285;
  wire _3287 = _3280 ^ _3286;
  wire _3288 = _3275 ^ _3287;
  wire _3289 = uncoded_block[202] ^ uncoded_block[203];
  wire _3290 = _952 ^ _3289;
  wire _3291 = uncoded_block[204] ^ uncoded_block[206];
  wire _3292 = uncoded_block[210] ^ uncoded_block[211];
  wire _3293 = _3291 ^ _3292;
  wire _3294 = _3290 ^ _3293;
  wire _3295 = uncoded_block[212] ^ uncoded_block[214];
  wire _3296 = uncoded_block[215] ^ uncoded_block[216];
  wire _3297 = _3295 ^ _3296;
  wire _3298 = uncoded_block[219] ^ uncoded_block[222];
  wire _3299 = uncoded_block[225] ^ uncoded_block[226];
  wire _3300 = _3298 ^ _3299;
  wire _3301 = _3297 ^ _3300;
  wire _3302 = _3294 ^ _3301;
  wire _3303 = uncoded_block[227] ^ uncoded_block[232];
  wire _3304 = _3303 ^ _2550;
  wire _3305 = uncoded_block[236] ^ uncoded_block[238];
  wire _3306 = _3305 ^ _112;
  wire _3307 = _3304 ^ _3306;
  wire _3308 = uncoded_block[244] ^ uncoded_block[249];
  wire _3309 = uncoded_block[252] ^ uncoded_block[254];
  wire _3310 = _3308 ^ _3309;
  wire _3311 = uncoded_block[255] ^ uncoded_block[256];
  wire _3312 = uncoded_block[257] ^ uncoded_block[260];
  wire _3313 = _3311 ^ _3312;
  wire _3314 = _3310 ^ _3313;
  wire _3315 = _3307 ^ _3314;
  wire _3316 = _3302 ^ _3315;
  wire _3317 = _3288 ^ _3316;
  wire _3318 = _3261 ^ _3317;
  wire _3319 = _120 ^ _127;
  wire _3320 = uncoded_block[271] ^ uncoded_block[272];
  wire _3321 = uncoded_block[273] ^ uncoded_block[274];
  wire _3322 = _3320 ^ _3321;
  wire _3323 = _3319 ^ _3322;
  wire _3324 = uncoded_block[275] ^ uncoded_block[278];
  wire _3325 = uncoded_block[279] ^ uncoded_block[285];
  wire _3326 = _3324 ^ _3325;
  wire _3327 = uncoded_block[286] ^ uncoded_block[288];
  wire _3328 = uncoded_block[291] ^ uncoded_block[293];
  wire _3329 = _3327 ^ _3328;
  wire _3330 = _3326 ^ _3329;
  wire _3331 = _3323 ^ _3330;
  wire _3332 = uncoded_block[296] ^ uncoded_block[299];
  wire _3333 = _3332 ^ _999;
  wire _3334 = uncoded_block[307] ^ uncoded_block[308];
  wire _3335 = _1000 ^ _3334;
  wire _3336 = _3333 ^ _3335;
  wire _3337 = uncoded_block[309] ^ uncoded_block[310];
  wire _3338 = uncoded_block[311] ^ uncoded_block[313];
  wire _3339 = _3337 ^ _3338;
  wire _3340 = uncoded_block[314] ^ uncoded_block[315];
  wire _3341 = uncoded_block[316] ^ uncoded_block[318];
  wire _3342 = _3340 ^ _3341;
  wire _3343 = _3339 ^ _3342;
  wire _3344 = _3336 ^ _3343;
  wire _3345 = _3331 ^ _3344;
  wire _3346 = uncoded_block[321] ^ uncoded_block[322];
  wire _3347 = uncoded_block[323] ^ uncoded_block[324];
  wire _3348 = _3346 ^ _3347;
  wire _3349 = uncoded_block[328] ^ uncoded_block[332];
  wire _3350 = _152 ^ _3349;
  wire _3351 = _3348 ^ _3350;
  wire _3352 = uncoded_block[333] ^ uncoded_block[334];
  wire _3353 = uncoded_block[337] ^ uncoded_block[341];
  wire _3354 = _3352 ^ _3353;
  wire _3355 = uncoded_block[342] ^ uncoded_block[344];
  wire _3356 = _3355 ^ _159;
  wire _3357 = _3354 ^ _3356;
  wire _3358 = _3351 ^ _3357;
  wire _3359 = uncoded_block[348] ^ uncoded_block[349];
  wire _3360 = _3359 ^ _1024;
  wire _3361 = uncoded_block[355] ^ uncoded_block[356];
  wire _3362 = uncoded_block[357] ^ uncoded_block[358];
  wire _3363 = _3361 ^ _3362;
  wire _3364 = _3360 ^ _3363;
  wire _3365 = uncoded_block[359] ^ uncoded_block[361];
  wire _3366 = uncoded_block[362] ^ uncoded_block[364];
  wire _3367 = _3365 ^ _3366;
  wire _3368 = uncoded_block[365] ^ uncoded_block[367];
  wire _3369 = uncoded_block[368] ^ uncoded_block[369];
  wire _3370 = _3368 ^ _3369;
  wire _3371 = _3367 ^ _3370;
  wire _3372 = _3364 ^ _3371;
  wire _3373 = _3358 ^ _3372;
  wire _3374 = _3345 ^ _3373;
  wire _3375 = uncoded_block[373] ^ uncoded_block[379];
  wire _3376 = _1838 ^ _3375;
  wire _3377 = uncoded_block[383] ^ uncoded_block[384];
  wire _3378 = _1841 ^ _3377;
  wire _3379 = _3376 ^ _3378;
  wire _3380 = uncoded_block[385] ^ uncoded_block[386];
  wire _3381 = uncoded_block[388] ^ uncoded_block[389];
  wire _3382 = _3380 ^ _3381;
  wire _3383 = uncoded_block[392] ^ uncoded_block[393];
  wire _3384 = uncoded_block[395] ^ uncoded_block[396];
  wire _3385 = _3383 ^ _3384;
  wire _3386 = _3382 ^ _3385;
  wire _3387 = _3379 ^ _3386;
  wire _3388 = uncoded_block[397] ^ uncoded_block[400];
  wire _3389 = uncoded_block[402] ^ uncoded_block[406];
  wire _3390 = _3388 ^ _3389;
  wire _3391 = uncoded_block[407] ^ uncoded_block[408];
  wire _3392 = _3391 ^ _2629;
  wire _3393 = _3390 ^ _3392;
  wire _3394 = uncoded_block[411] ^ uncoded_block[412];
  wire _3395 = _3394 ^ _1055;
  wire _3396 = uncoded_block[416] ^ uncoded_block[417];
  wire _3397 = uncoded_block[419] ^ uncoded_block[421];
  wire _3398 = _3396 ^ _3397;
  wire _3399 = _3395 ^ _3398;
  wire _3400 = _3393 ^ _3399;
  wire _3401 = _3387 ^ _3400;
  wire _3402 = uncoded_block[429] ^ uncoded_block[434];
  wire _3403 = _1062 ^ _3402;
  wire _3404 = uncoded_block[436] ^ uncoded_block[438];
  wire _3405 = uncoded_block[439] ^ uncoded_block[440];
  wire _3406 = _3404 ^ _3405;
  wire _3407 = _3403 ^ _3406;
  wire _3408 = uncoded_block[441] ^ uncoded_block[443];
  wire _3409 = uncoded_block[446] ^ uncoded_block[448];
  wire _3410 = _3408 ^ _3409;
  wire _3411 = uncoded_block[449] ^ uncoded_block[450];
  wire _3412 = _3411 ^ _2650;
  wire _3413 = _3410 ^ _3412;
  wire _3414 = _3407 ^ _3413;
  wire _3415 = uncoded_block[458] ^ uncoded_block[459];
  wire _3416 = uncoded_block[466] ^ uncoded_block[468];
  wire _3417 = _3415 ^ _3416;
  wire _3418 = uncoded_block[470] ^ uncoded_block[471];
  wire _3419 = _3418 ^ _221;
  wire _3420 = _3417 ^ _3419;
  wire _3421 = uncoded_block[477] ^ uncoded_block[478];
  wire _3422 = _3421 ^ _1085;
  wire _3423 = uncoded_block[481] ^ uncoded_block[485];
  wire _3424 = uncoded_block[490] ^ uncoded_block[492];
  wire _3425 = _3423 ^ _3424;
  wire _3426 = _3422 ^ _3425;
  wire _3427 = _3420 ^ _3426;
  wire _3428 = _3414 ^ _3427;
  wire _3429 = _3401 ^ _3428;
  wire _3430 = _3374 ^ _3429;
  wire _3431 = _3318 ^ _3430;
  wire _3432 = uncoded_block[493] ^ uncoded_block[494];
  wire _3433 = _3432 ^ _1094;
  wire _3434 = uncoded_block[500] ^ uncoded_block[501];
  wire _3435 = _3434 ^ _2668;
  wire _3436 = _3433 ^ _3435;
  wire _3437 = uncoded_block[509] ^ uncoded_block[510];
  wire _3438 = _2671 ^ _3437;
  wire _3439 = uncoded_block[512] ^ uncoded_block[513];
  wire _3440 = uncoded_block[514] ^ uncoded_block[518];
  wire _3441 = _3439 ^ _3440;
  wire _3442 = _3438 ^ _3441;
  wire _3443 = _3436 ^ _3442;
  wire _3444 = uncoded_block[519] ^ uncoded_block[520];
  wire _3445 = uncoded_block[521] ^ uncoded_block[522];
  wire _3446 = _3444 ^ _3445;
  wire _3447 = uncoded_block[528] ^ uncoded_block[530];
  wire _3448 = _1900 ^ _3447;
  wire _3449 = _3446 ^ _3448;
  wire _3450 = uncoded_block[531] ^ uncoded_block[535];
  wire _3451 = uncoded_block[536] ^ uncoded_block[537];
  wire _3452 = _3450 ^ _3451;
  wire _3453 = uncoded_block[542] ^ uncoded_block[546];
  wire _3454 = uncoded_block[547] ^ uncoded_block[551];
  wire _3455 = _3453 ^ _3454;
  wire _3456 = _3452 ^ _3455;
  wire _3457 = _3449 ^ _3456;
  wire _3458 = _3443 ^ _3457;
  wire _3459 = uncoded_block[552] ^ uncoded_block[553];
  wire _3460 = _3459 ^ _1122;
  wire _3461 = uncoded_block[559] ^ uncoded_block[561];
  wire _3462 = _1123 ^ _3461;
  wire _3463 = _3460 ^ _3462;
  wire _3464 = uncoded_block[562] ^ uncoded_block[563];
  wire _3465 = uncoded_block[564] ^ uncoded_block[565];
  wire _3466 = _3464 ^ _3465;
  wire _3467 = uncoded_block[566] ^ uncoded_block[567];
  wire _3468 = uncoded_block[569] ^ uncoded_block[570];
  wire _3469 = _3467 ^ _3468;
  wire _3470 = _3466 ^ _3469;
  wire _3471 = _3463 ^ _3470;
  wire _3472 = uncoded_block[572] ^ uncoded_block[574];
  wire _3473 = _3472 ^ _1931;
  wire _3474 = uncoded_block[577] ^ uncoded_block[580];
  wire _3475 = uncoded_block[581] ^ uncoded_block[583];
  wire _3476 = _3474 ^ _3475;
  wire _3477 = _3473 ^ _3476;
  wire _3478 = uncoded_block[587] ^ uncoded_block[588];
  wire _3479 = _3478 ^ _1141;
  wire _3480 = uncoded_block[592] ^ uncoded_block[594];
  wire _3481 = _3480 ^ _1939;
  wire _3482 = _3479 ^ _3481;
  wire _3483 = _3477 ^ _3482;
  wire _3484 = _3471 ^ _3483;
  wire _3485 = _3458 ^ _3484;
  wire _3486 = uncoded_block[598] ^ uncoded_block[599];
  wire _3487 = uncoded_block[601] ^ uncoded_block[602];
  wire _3488 = _3486 ^ _3487;
  wire _3489 = uncoded_block[603] ^ uncoded_block[604];
  wire _3490 = _3489 ^ _1146;
  wire _3491 = _3488 ^ _3490;
  wire _3492 = uncoded_block[611] ^ uncoded_block[615];
  wire _3493 = _2713 ^ _3492;
  wire _3494 = uncoded_block[617] ^ uncoded_block[620];
  wire _3495 = uncoded_block[621] ^ uncoded_block[622];
  wire _3496 = _3494 ^ _3495;
  wire _3497 = _3493 ^ _3496;
  wire _3498 = _3491 ^ _3497;
  wire _3499 = uncoded_block[624] ^ uncoded_block[628];
  wire _3500 = _3499 ^ _289;
  wire _3501 = uncoded_block[633] ^ uncoded_block[634];
  wire _3502 = uncoded_block[636] ^ uncoded_block[640];
  wire _3503 = _3501 ^ _3502;
  wire _3504 = _3500 ^ _3503;
  wire _3505 = uncoded_block[644] ^ uncoded_block[646];
  wire _3506 = _294 ^ _3505;
  wire _3507 = uncoded_block[650] ^ uncoded_block[653];
  wire _3508 = uncoded_block[656] ^ uncoded_block[657];
  wire _3509 = _3507 ^ _3508;
  wire _3510 = _3506 ^ _3509;
  wire _3511 = _3504 ^ _3510;
  wire _3512 = _3498 ^ _3511;
  wire _3513 = uncoded_block[658] ^ uncoded_block[659];
  wire _3514 = uncoded_block[660] ^ uncoded_block[662];
  wire _3515 = _3513 ^ _3514;
  wire _3516 = uncoded_block[666] ^ uncoded_block[669];
  wire _3517 = _308 ^ _3516;
  wire _3518 = _3515 ^ _3517;
  wire _3519 = uncoded_block[673] ^ uncoded_block[676];
  wire _3520 = _1177 ^ _3519;
  wire _3521 = uncoded_block[677] ^ uncoded_block[679];
  wire _3522 = uncoded_block[681] ^ uncoded_block[682];
  wire _3523 = _3521 ^ _3522;
  wire _3524 = _3520 ^ _3523;
  wire _3525 = _3518 ^ _3524;
  wire _3526 = uncoded_block[683] ^ uncoded_block[684];
  wire _3527 = uncoded_block[685] ^ uncoded_block[689];
  wire _3528 = _3526 ^ _3527;
  wire _3529 = uncoded_block[696] ^ uncoded_block[697];
  wire _3530 = _1186 ^ _3529;
  wire _3531 = _3528 ^ _3530;
  wire _3532 = uncoded_block[699] ^ uncoded_block[701];
  wire _3533 = uncoded_block[705] ^ uncoded_block[706];
  wire _3534 = _3532 ^ _3533;
  wire _3535 = uncoded_block[709] ^ uncoded_block[711];
  wire _3536 = uncoded_block[712] ^ uncoded_block[713];
  wire _3537 = _3535 ^ _3536;
  wire _3538 = _3534 ^ _3537;
  wire _3539 = _3531 ^ _3538;
  wire _3540 = _3525 ^ _3539;
  wire _3541 = _3512 ^ _3540;
  wire _3542 = _3485 ^ _3541;
  wire _3543 = _1194 ^ _341;
  wire _3544 = uncoded_block[724] ^ uncoded_block[725];
  wire _3545 = _3544 ^ _344;
  wire _3546 = _3543 ^ _3545;
  wire _3547 = uncoded_block[733] ^ uncoded_block[734];
  wire _3548 = _2768 ^ _3547;
  wire _3549 = uncoded_block[737] ^ uncoded_block[740];
  wire _3550 = uncoded_block[742] ^ uncoded_block[744];
  wire _3551 = _3549 ^ _3550;
  wire _3552 = _3548 ^ _3551;
  wire _3553 = _3546 ^ _3552;
  wire _3554 = uncoded_block[746] ^ uncoded_block[748];
  wire _3555 = _3554 ^ _1210;
  wire _3556 = uncoded_block[756] ^ uncoded_block[758];
  wire _3557 = _1214 ^ _3556;
  wire _3558 = _3555 ^ _3557;
  wire _3559 = uncoded_block[759] ^ uncoded_block[760];
  wire _3560 = _3559 ^ _1217;
  wire _3561 = uncoded_block[765] ^ uncoded_block[769];
  wire _3562 = uncoded_block[775] ^ uncoded_block[776];
  wire _3563 = _3561 ^ _3562;
  wire _3564 = _3560 ^ _3563;
  wire _3565 = _3558 ^ _3564;
  wire _3566 = _3553 ^ _3565;
  wire _3567 = uncoded_block[777] ^ uncoded_block[779];
  wire _3568 = uncoded_block[780] ^ uncoded_block[782];
  wire _3569 = _3567 ^ _3568;
  wire _3570 = uncoded_block[784] ^ uncoded_block[785];
  wire _3571 = uncoded_block[786] ^ uncoded_block[790];
  wire _3572 = _3570 ^ _3571;
  wire _3573 = _3569 ^ _3572;
  wire _3574 = uncoded_block[792] ^ uncoded_block[793];
  wire _3575 = _3574 ^ _375;
  wire _3576 = uncoded_block[797] ^ uncoded_block[800];
  wire _3577 = uncoded_block[803] ^ uncoded_block[804];
  wire _3578 = _3576 ^ _3577;
  wire _3579 = _3575 ^ _3578;
  wire _3580 = _3573 ^ _3579;
  wire _3581 = uncoded_block[805] ^ uncoded_block[807];
  wire _3582 = uncoded_block[809] ^ uncoded_block[812];
  wire _3583 = _3581 ^ _3582;
  wire _3584 = uncoded_block[818] ^ uncoded_block[822];
  wire _3585 = _1239 ^ _3584;
  wire _3586 = _3583 ^ _3585;
  wire _3587 = uncoded_block[823] ^ uncoded_block[824];
  wire _3588 = uncoded_block[825] ^ uncoded_block[827];
  wire _3589 = _3587 ^ _3588;
  wire _3590 = uncoded_block[830] ^ uncoded_block[831];
  wire _3591 = _2812 ^ _3590;
  wire _3592 = _3589 ^ _3591;
  wire _3593 = _3586 ^ _3592;
  wire _3594 = _3580 ^ _3593;
  wire _3595 = _3566 ^ _3594;
  wire _3596 = uncoded_block[835] ^ uncoded_block[839];
  wire _3597 = uncoded_block[844] ^ uncoded_block[845];
  wire _3598 = _3596 ^ _3597;
  wire _3599 = uncoded_block[847] ^ uncoded_block[848];
  wire _3600 = uncoded_block[855] ^ uncoded_block[856];
  wire _3601 = _3599 ^ _3600;
  wire _3602 = _3598 ^ _3601;
  wire _3603 = uncoded_block[860] ^ uncoded_block[861];
  wire _3604 = uncoded_block[863] ^ uncoded_block[869];
  wire _3605 = _3603 ^ _3604;
  wire _3606 = _3605 ^ _418;
  wire _3607 = _3602 ^ _3606;
  wire _3608 = uncoded_block[876] ^ uncoded_block[877];
  wire _3609 = _3608 ^ _2835;
  wire _3610 = uncoded_block[880] ^ uncoded_block[883];
  wire _3611 = _3610 ^ _423;
  wire _3612 = _3609 ^ _3611;
  wire _3613 = uncoded_block[886] ^ uncoded_block[890];
  wire _3614 = uncoded_block[892] ^ uncoded_block[894];
  wire _3615 = _3613 ^ _3614;
  wire _3616 = uncoded_block[895] ^ uncoded_block[897];
  wire _3617 = uncoded_block[898] ^ uncoded_block[900];
  wire _3618 = _3616 ^ _3617;
  wire _3619 = _3615 ^ _3618;
  wire _3620 = _3612 ^ _3619;
  wire _3621 = _3607 ^ _3620;
  wire _3622 = uncoded_block[902] ^ uncoded_block[905];
  wire _3623 = uncoded_block[906] ^ uncoded_block[907];
  wire _3624 = _3622 ^ _3623;
  wire _3625 = uncoded_block[911] ^ uncoded_block[914];
  wire _3626 = _432 ^ _3625;
  wire _3627 = _3624 ^ _3626;
  wire _3628 = uncoded_block[915] ^ uncoded_block[916];
  wire _3629 = uncoded_block[917] ^ uncoded_block[918];
  wire _3630 = _3628 ^ _3629;
  wire _3631 = uncoded_block[919] ^ uncoded_block[920];
  wire _3632 = uncoded_block[921] ^ uncoded_block[922];
  wire _3633 = _3631 ^ _3632;
  wire _3634 = _3630 ^ _3633;
  wire _3635 = _3627 ^ _3634;
  wire _3636 = _2855 ^ _2857;
  wire _3637 = uncoded_block[931] ^ uncoded_block[933];
  wire _3638 = uncoded_block[935] ^ uncoded_block[940];
  wire _3639 = _3637 ^ _3638;
  wire _3640 = _3636 ^ _3639;
  wire _3641 = uncoded_block[942] ^ uncoded_block[945];
  wire _3642 = _3641 ^ _456;
  wire _3643 = uncoded_block[948] ^ uncoded_block[952];
  wire _3644 = _3643 ^ _2089;
  wire _3645 = _3642 ^ _3644;
  wire _3646 = _3640 ^ _3645;
  wire _3647 = _3635 ^ _3646;
  wire _3648 = _3621 ^ _3647;
  wire _3649 = _3595 ^ _3648;
  wire _3650 = _3542 ^ _3649;
  wire _3651 = _3431 ^ _3650;
  wire _3652 = _1307 ^ _2871;
  wire _3653 = uncoded_block[962] ^ uncoded_block[966];
  wire _3654 = _3653 ^ _2093;
  wire _3655 = _3652 ^ _3654;
  wire _3656 = uncoded_block[969] ^ uncoded_block[972];
  wire _3657 = uncoded_block[975] ^ uncoded_block[976];
  wire _3658 = _3656 ^ _3657;
  wire _3659 = uncoded_block[983] ^ uncoded_block[984];
  wire _3660 = _3659 ^ _2102;
  wire _3661 = _3658 ^ _3660;
  wire _3662 = _3655 ^ _3661;
  wire _3663 = uncoded_block[991] ^ uncoded_block[993];
  wire _3664 = uncoded_block[994] ^ uncoded_block[1000];
  wire _3665 = _3663 ^ _3664;
  wire _3666 = uncoded_block[1005] ^ uncoded_block[1009];
  wire _3667 = _2112 ^ _3666;
  wire _3668 = _3665 ^ _3667;
  wire _3669 = _2890 ^ _1331;
  wire _3670 = uncoded_block[1019] ^ uncoded_block[1025];
  wire _3671 = _2893 ^ _3670;
  wire _3672 = _3669 ^ _3671;
  wire _3673 = _3668 ^ _3672;
  wire _3674 = _3662 ^ _3673;
  wire _3675 = uncoded_block[1029] ^ uncoded_block[1031];
  wire _3676 = uncoded_block[1032] ^ uncoded_block[1036];
  wire _3677 = _3675 ^ _3676;
  wire _3678 = uncoded_block[1037] ^ uncoded_block[1041];
  wire _3679 = _3678 ^ _2130;
  wire _3680 = _3677 ^ _3679;
  wire _3681 = uncoded_block[1046] ^ uncoded_block[1048];
  wire _3682 = uncoded_block[1052] ^ uncoded_block[1055];
  wire _3683 = _3681 ^ _3682;
  wire _3684 = uncoded_block[1060] ^ uncoded_block[1062];
  wire _3685 = uncoded_block[1063] ^ uncoded_block[1064];
  wire _3686 = _3684 ^ _3685;
  wire _3687 = _3683 ^ _3686;
  wire _3688 = _3680 ^ _3687;
  wire _3689 = uncoded_block[1067] ^ uncoded_block[1068];
  wire _3690 = _2921 ^ _3689;
  wire _3691 = uncoded_block[1069] ^ uncoded_block[1072];
  wire _3692 = uncoded_block[1073] ^ uncoded_block[1076];
  wire _3693 = _3691 ^ _3692;
  wire _3694 = _3690 ^ _3693;
  wire _3695 = uncoded_block[1077] ^ uncoded_block[1079];
  wire _3696 = uncoded_block[1086] ^ uncoded_block[1087];
  wire _3697 = _3695 ^ _3696;
  wire _3698 = uncoded_block[1094] ^ uncoded_block[1095];
  wire _3699 = _2930 ^ _3698;
  wire _3700 = _3697 ^ _3699;
  wire _3701 = _3694 ^ _3700;
  wire _3702 = _3688 ^ _3701;
  wire _3703 = _3674 ^ _3702;
  wire _3704 = uncoded_block[1096] ^ uncoded_block[1098];
  wire _3705 = uncoded_block[1099] ^ uncoded_block[1103];
  wire _3706 = _3704 ^ _3705;
  wire _3707 = uncoded_block[1104] ^ uncoded_block[1105];
  wire _3708 = uncoded_block[1106] ^ uncoded_block[1107];
  wire _3709 = _3707 ^ _3708;
  wire _3710 = _3706 ^ _3709;
  wire _3711 = uncoded_block[1108] ^ uncoded_block[1110];
  wire _3712 = _3711 ^ _1386;
  wire _3713 = uncoded_block[1115] ^ uncoded_block[1116];
  wire _3714 = uncoded_block[1119] ^ uncoded_block[1120];
  wire _3715 = _3713 ^ _3714;
  wire _3716 = _3712 ^ _3715;
  wire _3717 = _3710 ^ _3716;
  wire _3718 = uncoded_block[1122] ^ uncoded_block[1124];
  wire _3719 = _3718 ^ _558;
  wire _3720 = uncoded_block[1130] ^ uncoded_block[1137];
  wire _3721 = uncoded_block[1139] ^ uncoded_block[1140];
  wire _3722 = _3720 ^ _3721;
  wire _3723 = _3719 ^ _3722;
  wire _3724 = uncoded_block[1145] ^ uncoded_block[1147];
  wire _3725 = uncoded_block[1148] ^ uncoded_block[1150];
  wire _3726 = _3724 ^ _3725;
  wire _3727 = uncoded_block[1154] ^ uncoded_block[1155];
  wire _3728 = uncoded_block[1156] ^ uncoded_block[1157];
  wire _3729 = _3727 ^ _3728;
  wire _3730 = _3726 ^ _3729;
  wire _3731 = _3723 ^ _3730;
  wire _3732 = _3717 ^ _3731;
  wire _3733 = uncoded_block[1159] ^ uncoded_block[1161];
  wire _3734 = uncoded_block[1162] ^ uncoded_block[1164];
  wire _3735 = _3733 ^ _3734;
  wire _3736 = uncoded_block[1165] ^ uncoded_block[1166];
  wire _3737 = _3736 ^ _2189;
  wire _3738 = _3735 ^ _3737;
  wire _3739 = uncoded_block[1173] ^ uncoded_block[1174];
  wire _3740 = uncoded_block[1176] ^ uncoded_block[1178];
  wire _3741 = _3739 ^ _3740;
  wire _3742 = uncoded_block[1179] ^ uncoded_block[1180];
  wire _3743 = _3742 ^ _1417;
  wire _3744 = _3741 ^ _3743;
  wire _3745 = _3738 ^ _3744;
  wire _3746 = uncoded_block[1185] ^ uncoded_block[1186];
  wire _3747 = uncoded_block[1188] ^ uncoded_block[1190];
  wire _3748 = _3746 ^ _3747;
  wire _3749 = uncoded_block[1191] ^ uncoded_block[1192];
  wire _3750 = uncoded_block[1193] ^ uncoded_block[1198];
  wire _3751 = _3749 ^ _3750;
  wire _3752 = _3748 ^ _3751;
  wire _3753 = uncoded_block[1201] ^ uncoded_block[1204];
  wire _3754 = _2206 ^ _3753;
  wire _3755 = uncoded_block[1205] ^ uncoded_block[1208];
  wire _3756 = _3755 ^ _2217;
  wire _3757 = _3754 ^ _3756;
  wire _3758 = _3752 ^ _3757;
  wire _3759 = _3745 ^ _3758;
  wire _3760 = _3732 ^ _3759;
  wire _3761 = _3703 ^ _3760;
  wire _3762 = uncoded_block[1213] ^ uncoded_block[1214];
  wire _3763 = uncoded_block[1217] ^ uncoded_block[1218];
  wire _3764 = _3762 ^ _3763;
  wire _3765 = uncoded_block[1219] ^ uncoded_block[1220];
  wire _3766 = uncoded_block[1221] ^ uncoded_block[1223];
  wire _3767 = _3765 ^ _3766;
  wire _3768 = _3764 ^ _3767;
  wire _3769 = uncoded_block[1229] ^ uncoded_block[1232];
  wire _3770 = _612 ^ _3769;
  wire _3771 = uncoded_block[1235] ^ uncoded_block[1236];
  wire _3772 = uncoded_block[1237] ^ uncoded_block[1238];
  wire _3773 = _3771 ^ _3772;
  wire _3774 = _3770 ^ _3773;
  wire _3775 = _3768 ^ _3774;
  wire _3776 = uncoded_block[1240] ^ uncoded_block[1244];
  wire _3777 = uncoded_block[1245] ^ uncoded_block[1247];
  wire _3778 = _3776 ^ _3777;
  wire _3779 = uncoded_block[1248] ^ uncoded_block[1251];
  wire _3780 = uncoded_block[1253] ^ uncoded_block[1255];
  wire _3781 = _3779 ^ _3780;
  wire _3782 = _3778 ^ _3781;
  wire _3783 = uncoded_block[1256] ^ uncoded_block[1258];
  wire _3784 = uncoded_block[1260] ^ uncoded_block[1261];
  wire _3785 = _3783 ^ _3784;
  wire _3786 = uncoded_block[1265] ^ uncoded_block[1267];
  wire _3787 = _3004 ^ _3786;
  wire _3788 = _3785 ^ _3787;
  wire _3789 = _3782 ^ _3788;
  wire _3790 = _3775 ^ _3789;
  wire _3791 = uncoded_block[1273] ^ uncoded_block[1277];
  wire _3792 = _2245 ^ _3791;
  wire _3793 = uncoded_block[1278] ^ uncoded_block[1279];
  wire _3794 = uncoded_block[1280] ^ uncoded_block[1281];
  wire _3795 = _3793 ^ _3794;
  wire _3796 = _3792 ^ _3795;
  wire _3797 = uncoded_block[1283] ^ uncoded_block[1285];
  wire _3798 = uncoded_block[1286] ^ uncoded_block[1290];
  wire _3799 = _3797 ^ _3798;
  wire _3800 = uncoded_block[1291] ^ uncoded_block[1292];
  wire _3801 = uncoded_block[1294] ^ uncoded_block[1295];
  wire _3802 = _3800 ^ _3801;
  wire _3803 = _3799 ^ _3802;
  wire _3804 = _3796 ^ _3803;
  wire _3805 = uncoded_block[1303] ^ uncoded_block[1304];
  wire _3806 = _3017 ^ _3805;
  wire _3807 = uncoded_block[1307] ^ uncoded_block[1308];
  wire _3808 = uncoded_block[1310] ^ uncoded_block[1311];
  wire _3809 = _3807 ^ _3808;
  wire _3810 = _3806 ^ _3809;
  wire _3811 = uncoded_block[1314] ^ uncoded_block[1316];
  wire _3812 = uncoded_block[1317] ^ uncoded_block[1321];
  wire _3813 = _3811 ^ _3812;
  wire _3814 = uncoded_block[1322] ^ uncoded_block[1323];
  wire _3815 = _3814 ^ _1490;
  wire _3816 = _3813 ^ _3815;
  wire _3817 = _3810 ^ _3816;
  wire _3818 = _3804 ^ _3817;
  wire _3819 = _3790 ^ _3818;
  wire _3820 = uncoded_block[1332] ^ uncoded_block[1334];
  wire _3821 = _1494 ^ _3820;
  wire _3822 = uncoded_block[1337] ^ uncoded_block[1339];
  wire _3823 = uncoded_block[1341] ^ uncoded_block[1344];
  wire _3824 = _3822 ^ _3823;
  wire _3825 = _3821 ^ _3824;
  wire _3826 = uncoded_block[1348] ^ uncoded_block[1355];
  wire _3827 = _3039 ^ _3826;
  wire _3828 = uncoded_block[1364] ^ uncoded_block[1369];
  wire _3829 = _3045 ^ _3828;
  wire _3830 = _3827 ^ _3829;
  wire _3831 = _3825 ^ _3830;
  wire _3832 = uncoded_block[1370] ^ uncoded_block[1372];
  wire _3833 = _3832 ^ _2290;
  wire _3834 = uncoded_block[1381] ^ uncoded_block[1382];
  wire _3835 = uncoded_block[1383] ^ uncoded_block[1385];
  wire _3836 = _3834 ^ _3835;
  wire _3837 = _3833 ^ _3836;
  wire _3838 = uncoded_block[1387] ^ uncoded_block[1389];
  wire _3839 = _3838 ^ _692;
  wire _3840 = uncoded_block[1394] ^ uncoded_block[1396];
  wire _3841 = uncoded_block[1400] ^ uncoded_block[1402];
  wire _3842 = _3840 ^ _3841;
  wire _3843 = _3839 ^ _3842;
  wire _3844 = _3837 ^ _3843;
  wire _3845 = _3831 ^ _3844;
  wire _3846 = uncoded_block[1403] ^ uncoded_block[1404];
  wire _3847 = uncoded_block[1405] ^ uncoded_block[1406];
  wire _3848 = _3846 ^ _3847;
  wire _3849 = uncoded_block[1408] ^ uncoded_block[1410];
  wire _3850 = uncoded_block[1417] ^ uncoded_block[1420];
  wire _3851 = _3849 ^ _3850;
  wire _3852 = _3848 ^ _3851;
  wire _3853 = uncoded_block[1421] ^ uncoded_block[1423];
  wire _3854 = uncoded_block[1424] ^ uncoded_block[1430];
  wire _3855 = _3853 ^ _3854;
  wire _3856 = uncoded_block[1431] ^ uncoded_block[1434];
  wire _3857 = uncoded_block[1436] ^ uncoded_block[1437];
  wire _3858 = _3856 ^ _3857;
  wire _3859 = _3855 ^ _3858;
  wire _3860 = _3852 ^ _3859;
  wire _3861 = uncoded_block[1439] ^ uncoded_block[1440];
  wire _3862 = uncoded_block[1443] ^ uncoded_block[1446];
  wire _3863 = _3861 ^ _3862;
  wire _3864 = uncoded_block[1447] ^ uncoded_block[1448];
  wire _3865 = uncoded_block[1449] ^ uncoded_block[1450];
  wire _3866 = _3864 ^ _3865;
  wire _3867 = _3863 ^ _3866;
  wire _3868 = uncoded_block[1455] ^ uncoded_block[1457];
  wire _3869 = _2328 ^ _3868;
  wire _3870 = uncoded_block[1460] ^ uncoded_block[1461];
  wire _3871 = uncoded_block[1462] ^ uncoded_block[1464];
  wire _3872 = _3870 ^ _3871;
  wire _3873 = _3869 ^ _3872;
  wire _3874 = _3867 ^ _3873;
  wire _3875 = _3860 ^ _3874;
  wire _3876 = _3845 ^ _3875;
  wire _3877 = _3819 ^ _3876;
  wire _3878 = _3761 ^ _3877;
  wire _3879 = uncoded_block[1467] ^ uncoded_block[1469];
  wire _3880 = _1548 ^ _3879;
  wire _3881 = uncoded_block[1475] ^ uncoded_block[1476];
  wire _3882 = _1551 ^ _3881;
  wire _3883 = _3880 ^ _3882;
  wire _3884 = uncoded_block[1479] ^ uncoded_block[1480];
  wire _3885 = uncoded_block[1482] ^ uncoded_block[1485];
  wire _3886 = _3884 ^ _3885;
  wire _3887 = _740 ^ _3103;
  wire _3888 = _3886 ^ _3887;
  wire _3889 = _3883 ^ _3888;
  wire _3890 = uncoded_block[1495] ^ uncoded_block[1496];
  wire _3891 = uncoded_block[1499] ^ uncoded_block[1501];
  wire _3892 = _3890 ^ _3891;
  wire _3893 = uncoded_block[1502] ^ uncoded_block[1504];
  wire _3894 = uncoded_block[1505] ^ uncoded_block[1506];
  wire _3895 = _3893 ^ _3894;
  wire _3896 = _3892 ^ _3895;
  wire _3897 = uncoded_block[1508] ^ uncoded_block[1517];
  wire _3898 = uncoded_block[1518] ^ uncoded_block[1521];
  wire _3899 = _3897 ^ _3898;
  wire _3900 = uncoded_block[1522] ^ uncoded_block[1524];
  wire _3901 = _3900 ^ _3122;
  wire _3902 = _3899 ^ _3901;
  wire _3903 = _3896 ^ _3902;
  wire _3904 = _3889 ^ _3903;
  wire _3905 = uncoded_block[1532] ^ uncoded_block[1534];
  wire _3906 = uncoded_block[1536] ^ uncoded_block[1537];
  wire _3907 = _3905 ^ _3906;
  wire _3908 = uncoded_block[1538] ^ uncoded_block[1539];
  wire _3909 = uncoded_block[1540] ^ uncoded_block[1543];
  wire _3910 = _3908 ^ _3909;
  wire _3911 = _3907 ^ _3910;
  wire _3912 = uncoded_block[1546] ^ uncoded_block[1550];
  wire _3913 = _3912 ^ _769;
  wire _3914 = uncoded_block[1556] ^ uncoded_block[1558];
  wire _3915 = _3914 ^ _1597;
  wire _3916 = _3913 ^ _3915;
  wire _3917 = _3911 ^ _3916;
  wire _3918 = uncoded_block[1564] ^ uncoded_block[1572];
  wire _3919 = _774 ^ _3918;
  wire _3920 = uncoded_block[1575] ^ uncoded_block[1577];
  wire _3921 = uncoded_block[1578] ^ uncoded_block[1579];
  wire _3922 = _3920 ^ _3921;
  wire _3923 = _3919 ^ _3922;
  wire _3924 = uncoded_block[1580] ^ uncoded_block[1583];
  wire _3925 = uncoded_block[1584] ^ uncoded_block[1586];
  wire _3926 = _3924 ^ _3925;
  wire _3927 = uncoded_block[1587] ^ uncoded_block[1589];
  wire _3928 = _3927 ^ _791;
  wire _3929 = _3926 ^ _3928;
  wire _3930 = _3923 ^ _3929;
  wire _3931 = _3917 ^ _3930;
  wire _3932 = _3904 ^ _3931;
  wire _3933 = uncoded_block[1594] ^ uncoded_block[1596];
  wire _3934 = uncoded_block[1597] ^ uncoded_block[1600];
  wire _3935 = _3933 ^ _3934;
  wire _3936 = uncoded_block[1601] ^ uncoded_block[1603];
  wire _3937 = uncoded_block[1610] ^ uncoded_block[1612];
  wire _3938 = _3936 ^ _3937;
  wire _3939 = _3935 ^ _3938;
  wire _3940 = _1633 ^ _3160;
  wire _3941 = uncoded_block[1623] ^ uncoded_block[1624];
  wire _3942 = uncoded_block[1626] ^ uncoded_block[1628];
  wire _3943 = _3941 ^ _3942;
  wire _3944 = _3940 ^ _3943;
  wire _3945 = _3939 ^ _3944;
  wire _3946 = uncoded_block[1633] ^ uncoded_block[1635];
  wire _3947 = _1639 ^ _3946;
  wire _3948 = uncoded_block[1639] ^ uncoded_block[1640];
  wire _3949 = _1642 ^ _3948;
  wire _3950 = _3947 ^ _3949;
  wire _3951 = uncoded_block[1641] ^ uncoded_block[1644];
  wire _3952 = _3951 ^ _2412;
  wire _3953 = uncoded_block[1649] ^ uncoded_block[1653];
  wire _3954 = _3953 ^ _3174;
  wire _3955 = _3952 ^ _3954;
  wire _3956 = _3950 ^ _3955;
  wire _3957 = _3945 ^ _3956;
  wire _3958 = uncoded_block[1659] ^ uncoded_block[1662];
  wire _3959 = uncoded_block[1663] ^ uncoded_block[1671];
  wire _3960 = _3958 ^ _3959;
  wire _3961 = uncoded_block[1672] ^ uncoded_block[1676];
  wire _3962 = uncoded_block[1677] ^ uncoded_block[1678];
  wire _3963 = _3961 ^ _3962;
  wire _3964 = _3960 ^ _3963;
  wire _3965 = uncoded_block[1684] ^ uncoded_block[1686];
  wire _3966 = _1663 ^ _3965;
  wire _3967 = uncoded_block[1689] ^ uncoded_block[1690];
  wire _3968 = uncoded_block[1692] ^ uncoded_block[1694];
  wire _3969 = _3967 ^ _3968;
  wire _3970 = _3966 ^ _3969;
  wire _3971 = _3964 ^ _3970;
  wire _3972 = uncoded_block[1695] ^ uncoded_block[1696];
  wire _3973 = uncoded_block[1699] ^ uncoded_block[1700];
  wire _3974 = _3972 ^ _3973;
  wire _3975 = uncoded_block[1701] ^ uncoded_block[1703];
  wire _3976 = uncoded_block[1704] ^ uncoded_block[1705];
  wire _3977 = _3975 ^ _3976;
  wire _3978 = _3974 ^ _3977;
  wire _3979 = uncoded_block[1706] ^ uncoded_block[1709];
  wire _3980 = uncoded_block[1710] ^ uncoded_block[1712];
  wire _3981 = _3979 ^ _3980;
  wire _3982 = _3200 ^ _1677;
  wire _3983 = _3981 ^ _3982;
  wire _3984 = _3978 ^ _3983;
  wire _3985 = _3971 ^ _3984;
  wire _3986 = _3957 ^ _3985;
  wire _3987 = _3932 ^ _3986;
  wire _3988 = uncoded_block[1718] ^ uncoded_block[1719];
  wire _3989 = _3988 ^ uncoded_block[1722];
  wire _3990 = _3987 ^ _3989;
  wire _3991 = _3878 ^ _3990;
  wire _3992 = _3651 ^ _3991;
  wire _3993 = uncoded_block[6] ^ uncoded_block[7];
  wire _3994 = _1683 ^ _3993;
  wire _3995 = uncoded_block[8] ^ uncoded_block[9];
  wire _3996 = _3995 ^ _1686;
  wire _3997 = _3994 ^ _3996;
  wire _3998 = uncoded_block[14] ^ uncoded_block[16];
  wire _3999 = _3998 ^ _3217;
  wire _4000 = uncoded_block[22] ^ uncoded_block[23];
  wire _4001 = uncoded_block[24] ^ uncoded_block[25];
  wire _4002 = _4000 ^ _4001;
  wire _4003 = _3999 ^ _4002;
  wire _4004 = _3997 ^ _4003;
  wire _4005 = uncoded_block[26] ^ uncoded_block[33];
  wire _4006 = _4005 ^ _3227;
  wire _4007 = _4006 ^ _20;
  wire _4008 = uncoded_block[41] ^ uncoded_block[42];
  wire _4009 = uncoded_block[43] ^ uncoded_block[46];
  wire _4010 = _4008 ^ _4009;
  wire _4011 = _4010 ^ _3234;
  wire _4012 = _4007 ^ _4011;
  wire _4013 = _4004 ^ _4012;
  wire _4014 = uncoded_block[52] ^ uncoded_block[53];
  wire _4015 = uncoded_block[54] ^ uncoded_block[63];
  wire _4016 = _4014 ^ _4015;
  wire _4017 = uncoded_block[68] ^ uncoded_block[71];
  wire _4018 = _1706 ^ _4017;
  wire _4019 = _4016 ^ _4018;
  wire _4020 = uncoded_block[74] ^ uncoded_block[75];
  wire _4021 = _897 ^ _4020;
  wire _4022 = _1714 ^ _41;
  wire _4023 = _4021 ^ _4022;
  wire _4024 = _4019 ^ _4023;
  wire _4025 = uncoded_block[84] ^ uncoded_block[87];
  wire _4026 = uncoded_block[94] ^ uncoded_block[95];
  wire _4027 = _4025 ^ _4026;
  wire _4028 = uncoded_block[101] ^ uncoded_block[102];
  wire _4029 = _3249 ^ _4028;
  wire _4030 = _4027 ^ _4029;
  wire _4031 = uncoded_block[103] ^ uncoded_block[106];
  wire _4032 = uncoded_block[107] ^ uncoded_block[110];
  wire _4033 = _4031 ^ _4032;
  wire _4034 = uncoded_block[111] ^ uncoded_block[112];
  wire _4035 = _4034 ^ _3253;
  wire _4036 = _4033 ^ _4035;
  wire _4037 = _4030 ^ _4036;
  wire _4038 = _4024 ^ _4037;
  wire _4039 = _4013 ^ _4038;
  wire _4040 = uncoded_block[117] ^ uncoded_block[124];
  wire _4041 = _4040 ^ _57;
  wire _4042 = uncoded_block[130] ^ uncoded_block[132];
  wire _4043 = uncoded_block[140] ^ uncoded_block[143];
  wire _4044 = _4042 ^ _4043;
  wire _4045 = _4041 ^ _4044;
  wire _4046 = uncoded_block[146] ^ uncoded_block[147];
  wire _4047 = _4046 ^ _1745;
  wire _4048 = uncoded_block[154] ^ uncoded_block[156];
  wire _4049 = uncoded_block[158] ^ uncoded_block[159];
  wire _4050 = _4048 ^ _4049;
  wire _4051 = _4047 ^ _4050;
  wire _4052 = _4045 ^ _4051;
  wire _4053 = uncoded_block[162] ^ uncoded_block[163];
  wire _4054 = uncoded_block[164] ^ uncoded_block[165];
  wire _4055 = _4053 ^ _4054;
  wire _4056 = uncoded_block[166] ^ uncoded_block[169];
  wire _4057 = uncoded_block[173] ^ uncoded_block[177];
  wire _4058 = _4056 ^ _4057;
  wire _4059 = _4055 ^ _4058;
  wire _4060 = uncoded_block[178] ^ uncoded_block[182];
  wire _4061 = _4060 ^ _2528;
  wire _4062 = uncoded_block[186] ^ uncoded_block[187];
  wire _4063 = _4062 ^ _947;
  wire _4064 = _4061 ^ _4063;
  wire _4065 = _4059 ^ _4064;
  wire _4066 = _4052 ^ _4065;
  wire _4067 = uncoded_block[192] ^ uncoded_block[196];
  wire _4068 = uncoded_block[197] ^ uncoded_block[201];
  wire _4069 = _4067 ^ _4068;
  wire _4070 = uncoded_block[204] ^ uncoded_block[205];
  wire _4071 = uncoded_block[209] ^ uncoded_block[212];
  wire _4072 = _4070 ^ _4071;
  wire _4073 = _4069 ^ _4072;
  wire _4074 = uncoded_block[216] ^ uncoded_block[217];
  wire _4075 = _1767 ^ _4074;
  wire _4076 = uncoded_block[223] ^ uncoded_block[224];
  wire _4077 = _2543 ^ _4076;
  wire _4078 = _4075 ^ _4077;
  wire _4079 = _4073 ^ _4078;
  wire _4080 = uncoded_block[227] ^ uncoded_block[229];
  wire _4081 = uncoded_block[230] ^ uncoded_block[231];
  wire _4082 = _4080 ^ _4081;
  wire _4083 = _4082 ^ _969;
  wire _4084 = uncoded_block[236] ^ uncoded_block[241];
  wire _4085 = uncoded_block[243] ^ uncoded_block[245];
  wire _4086 = _4084 ^ _4085;
  wire _4087 = uncoded_block[247] ^ uncoded_block[251];
  wire _4088 = uncoded_block[254] ^ uncoded_block[258];
  wire _4089 = _4087 ^ _4088;
  wire _4090 = _4086 ^ _4089;
  wire _4091 = _4083 ^ _4090;
  wire _4092 = _4079 ^ _4091;
  wire _4093 = _4066 ^ _4092;
  wire _4094 = _4039 ^ _4093;
  wire _4095 = uncoded_block[259] ^ uncoded_block[261];
  wire _4096 = uncoded_block[262] ^ uncoded_block[263];
  wire _4097 = _4095 ^ _4096;
  wire _4098 = uncoded_block[264] ^ uncoded_block[266];
  wire _4099 = uncoded_block[267] ^ uncoded_block[270];
  wire _4100 = _4098 ^ _4099;
  wire _4101 = _4097 ^ _4100;
  wire _4102 = uncoded_block[271] ^ uncoded_block[273];
  wire _4103 = uncoded_block[276] ^ uncoded_block[279];
  wire _4104 = _4102 ^ _4103;
  wire _4105 = uncoded_block[283] ^ uncoded_block[284];
  wire _4106 = _4105 ^ _991;
  wire _4107 = _4104 ^ _4106;
  wire _4108 = _4101 ^ _4107;
  wire _4109 = _992 ^ _2573;
  wire _4110 = uncoded_block[296] ^ uncoded_block[298];
  wire _4111 = uncoded_block[302] ^ uncoded_block[303];
  wire _4112 = _4110 ^ _4111;
  wire _4113 = _4109 ^ _4112;
  wire _4114 = uncoded_block[305] ^ uncoded_block[307];
  wire _4115 = uncoded_block[308] ^ uncoded_block[310];
  wire _4116 = _4114 ^ _4115;
  wire _4117 = uncoded_block[312] ^ uncoded_block[313];
  wire _4118 = uncoded_block[317] ^ uncoded_block[320];
  wire _4119 = _4117 ^ _4118;
  wire _4120 = _4116 ^ _4119;
  wire _4121 = _4113 ^ _4120;
  wire _4122 = _4108 ^ _4121;
  wire _4123 = uncoded_block[324] ^ uncoded_block[325];
  wire _4124 = _4123 ^ _2584;
  wire _4125 = uncoded_block[330] ^ uncoded_block[332];
  wire _4126 = uncoded_block[333] ^ uncoded_block[335];
  wire _4127 = _4125 ^ _4126;
  wire _4128 = _4124 ^ _4127;
  wire _4129 = uncoded_block[340] ^ uncoded_block[342];
  wire _4130 = _1825 ^ _4129;
  wire _4131 = uncoded_block[344] ^ uncoded_block[346];
  wire _4132 = uncoded_block[350] ^ uncoded_block[351];
  wire _4133 = _4131 ^ _4132;
  wire _4134 = _4130 ^ _4133;
  wire _4135 = _4128 ^ _4134;
  wire _4136 = _162 ^ _2602;
  wire _4137 = uncoded_block[358] ^ uncoded_block[363];
  wire _4138 = _4137 ^ _168;
  wire _4139 = _4136 ^ _4138;
  wire _4140 = uncoded_block[371] ^ uncoded_block[373];
  wire _4141 = uncoded_block[374] ^ uncoded_block[376];
  wire _4142 = _4140 ^ _4141;
  wire _4143 = uncoded_block[377] ^ uncoded_block[380];
  wire _4144 = _4143 ^ _2612;
  wire _4145 = _4142 ^ _4144;
  wire _4146 = _4139 ^ _4145;
  wire _4147 = _4135 ^ _4146;
  wire _4148 = _4122 ^ _4147;
  wire _4149 = uncoded_block[386] ^ uncoded_block[387];
  wire _4150 = _1039 ^ _4149;
  wire _4151 = uncoded_block[389] ^ uncoded_block[392];
  wire _4152 = uncoded_block[393] ^ uncoded_block[394];
  wire _4153 = _4151 ^ _4152;
  wire _4154 = _4150 ^ _4153;
  wire _4155 = uncoded_block[399] ^ uncoded_block[401];
  wire _4156 = uncoded_block[402] ^ uncoded_block[405];
  wire _4157 = _4155 ^ _4156;
  wire _4158 = _184 ^ _190;
  wire _4159 = _4157 ^ _4158;
  wire _4160 = _4154 ^ _4159;
  wire _4161 = uncoded_block[417] ^ uncoded_block[419];
  wire _4162 = _2630 ^ _4161;
  wire _4163 = uncoded_block[420] ^ uncoded_block[421];
  wire _4164 = uncoded_block[422] ^ uncoded_block[423];
  wire _4165 = _4163 ^ _4164;
  wire _4166 = _4162 ^ _4165;
  wire _4167 = uncoded_block[429] ^ uncoded_block[430];
  wire _4168 = _2633 ^ _4167;
  wire _4169 = uncoded_block[436] ^ uncoded_block[437];
  wire _4170 = _200 ^ _4169;
  wire _4171 = _4168 ^ _4170;
  wire _4172 = _4166 ^ _4171;
  wire _4173 = _4160 ^ _4172;
  wire _4174 = uncoded_block[442] ^ uncoded_block[446];
  wire _4175 = _3405 ^ _4174;
  wire _4176 = uncoded_block[448] ^ uncoded_block[449];
  wire _4177 = uncoded_block[451] ^ uncoded_block[452];
  wire _4178 = _4176 ^ _4177;
  wire _4179 = _4175 ^ _4178;
  wire _4180 = _1075 ^ _212;
  wire _4181 = uncoded_block[461] ^ uncoded_block[462];
  wire _4182 = _213 ^ _4181;
  wire _4183 = _4180 ^ _4182;
  wire _4184 = _4179 ^ _4183;
  wire _4185 = uncoded_block[463] ^ uncoded_block[464];
  wire _4186 = uncoded_block[469] ^ uncoded_block[470];
  wire _4187 = _4185 ^ _4186;
  wire _4188 = uncoded_block[472] ^ uncoded_block[473];
  wire _4189 = uncoded_block[474] ^ uncoded_block[476];
  wire _4190 = _4188 ^ _4189;
  wire _4191 = _4187 ^ _4190;
  wire _4192 = uncoded_block[477] ^ uncoded_block[481];
  wire _4193 = _4192 ^ _1090;
  wire _4194 = uncoded_block[487] ^ uncoded_block[489];
  wire _4195 = uncoded_block[494] ^ uncoded_block[499];
  wire _4196 = _4194 ^ _4195;
  wire _4197 = _4193 ^ _4196;
  wire _4198 = _4191 ^ _4197;
  wire _4199 = _4184 ^ _4198;
  wire _4200 = _4173 ^ _4199;
  wire _4201 = _4148 ^ _4200;
  wire _4202 = _4094 ^ _4201;
  wire _4203 = uncoded_block[500] ^ uncoded_block[505];
  wire _4204 = _4203 ^ _1892;
  wire _4205 = uncoded_block[508] ^ uncoded_block[511];
  wire _4206 = _4205 ^ _3439;
  wire _4207 = _4204 ^ _4206;
  wire _4208 = uncoded_block[516] ^ uncoded_block[518];
  wire _4209 = _232 ^ _4208;
  wire _4210 = uncoded_block[521] ^ uncoded_block[525];
  wire _4211 = _4210 ^ _1900;
  wire _4212 = _4209 ^ _4211;
  wire _4213 = _4207 ^ _4212;
  wire _4214 = uncoded_block[529] ^ uncoded_block[532];
  wire _4215 = uncoded_block[533] ^ uncoded_block[537];
  wire _4216 = _4214 ^ _4215;
  wire _4217 = uncoded_block[539] ^ uncoded_block[540];
  wire _4218 = uncoded_block[541] ^ uncoded_block[548];
  wire _4219 = _4217 ^ _4218;
  wire _4220 = _4216 ^ _4219;
  wire _4221 = uncoded_block[561] ^ uncoded_block[565];
  wire _4222 = _247 ^ _4221;
  wire _4223 = uncoded_block[569] ^ uncoded_block[571];
  wire _4224 = uncoded_block[572] ^ uncoded_block[573];
  wire _4225 = _4223 ^ _4224;
  wire _4226 = _4222 ^ _4225;
  wire _4227 = _4220 ^ _4226;
  wire _4228 = _4213 ^ _4227;
  wire _4229 = uncoded_block[578] ^ uncoded_block[581];
  wire _4230 = _1132 ^ _4229;
  wire _4231 = _1933 ^ _1139;
  wire _4232 = _4230 ^ _4231;
  wire _4233 = uncoded_block[587] ^ uncoded_block[589];
  wire _4234 = uncoded_block[590] ^ uncoded_block[591];
  wire _4235 = _4233 ^ _4234;
  wire _4236 = uncoded_block[593] ^ uncoded_block[595];
  wire _4237 = _4236 ^ _1142;
  wire _4238 = _4235 ^ _4237;
  wire _4239 = _4232 ^ _4238;
  wire _4240 = uncoded_block[606] ^ uncoded_block[608];
  wire _4241 = _1145 ^ _4240;
  wire _4242 = uncoded_block[611] ^ uncoded_block[613];
  wire _4243 = uncoded_block[618] ^ uncoded_block[619];
  wire _4244 = _4242 ^ _4243;
  wire _4245 = _4241 ^ _4244;
  wire _4246 = uncoded_block[621] ^ uncoded_block[623];
  wire _4247 = uncoded_block[625] ^ uncoded_block[629];
  wire _4248 = _4246 ^ _4247;
  wire _4249 = uncoded_block[636] ^ uncoded_block[638];
  wire _4250 = _1157 ^ _4249;
  wire _4251 = _4248 ^ _4250;
  wire _4252 = _4245 ^ _4251;
  wire _4253 = _4239 ^ _4252;
  wire _4254 = _4228 ^ _4253;
  wire _4255 = uncoded_block[639] ^ uncoded_block[640];
  wire _4256 = uncoded_block[643] ^ uncoded_block[645];
  wire _4257 = _4255 ^ _4256;
  wire _4258 = uncoded_block[652] ^ uncoded_block[656];
  wire _4259 = _297 ^ _4258;
  wire _4260 = _4257 ^ _4259;
  wire _4261 = uncoded_block[659] ^ uncoded_block[660];
  wire _4262 = uncoded_block[662] ^ uncoded_block[664];
  wire _4263 = _4261 ^ _4262;
  wire _4264 = uncoded_block[666] ^ uncoded_block[668];
  wire _4265 = uncoded_block[669] ^ uncoded_block[672];
  wire _4266 = _4264 ^ _4265;
  wire _4267 = _4263 ^ _4266;
  wire _4268 = _4260 ^ _4267;
  wire _4269 = uncoded_block[673] ^ uncoded_block[682];
  wire _4270 = _4269 ^ _321;
  wire _4271 = uncoded_block[687] ^ uncoded_block[688];
  wire _4272 = uncoded_block[692] ^ uncoded_block[693];
  wire _4273 = _4271 ^ _4272;
  wire _4274 = _4270 ^ _4273;
  wire _4275 = uncoded_block[697] ^ uncoded_block[700];
  wire _4276 = _328 ^ _4275;
  wire _4277 = _3533 ^ _3535;
  wire _4278 = _4276 ^ _4277;
  wire _4279 = _4274 ^ _4278;
  wire _4280 = _4268 ^ _4279;
  wire _4281 = uncoded_block[716] ^ uncoded_block[720];
  wire _4282 = _1194 ^ _4281;
  wire _4283 = uncoded_block[724] ^ uncoded_block[726];
  wire _4284 = _343 ^ _4283;
  wire _4285 = _4282 ^ _4284;
  wire _4286 = uncoded_block[727] ^ uncoded_block[729];
  wire _4287 = uncoded_block[731] ^ uncoded_block[733];
  wire _4288 = _4286 ^ _4287;
  wire _4289 = uncoded_block[739] ^ uncoded_block[741];
  wire _4290 = _1206 ^ _4289;
  wire _4291 = _4288 ^ _4290;
  wire _4292 = _4285 ^ _4291;
  wire _4293 = uncoded_block[748] ^ uncoded_block[750];
  wire _4294 = _1209 ^ _4293;
  wire _4295 = uncoded_block[751] ^ uncoded_block[752];
  wire _4296 = _4295 ^ _2778;
  wire _4297 = _4294 ^ _4296;
  wire _4298 = uncoded_block[757] ^ uncoded_block[758];
  wire _4299 = uncoded_block[759] ^ uncoded_block[761];
  wire _4300 = _4298 ^ _4299;
  wire _4301 = uncoded_block[765] ^ uncoded_block[766];
  wire _4302 = _1217 ^ _4301;
  wire _4303 = _4300 ^ _4302;
  wire _4304 = _4297 ^ _4303;
  wire _4305 = _4292 ^ _4304;
  wire _4306 = _4280 ^ _4305;
  wire _4307 = _4254 ^ _4306;
  wire _4308 = uncoded_block[770] ^ uncoded_block[780];
  wire _4309 = uncoded_block[783] ^ uncoded_block[784];
  wire _4310 = _4308 ^ _4309;
  wire _4311 = uncoded_block[788] ^ uncoded_block[789];
  wire _4312 = _371 ^ _4311;
  wire _4313 = _4310 ^ _4312;
  wire _4314 = uncoded_block[791] ^ uncoded_block[793];
  wire _4315 = _4314 ^ _1233;
  wire _4316 = uncoded_block[798] ^ uncoded_block[800];
  wire _4317 = uncoded_block[801] ^ uncoded_block[802];
  wire _4318 = _4316 ^ _4317;
  wire _4319 = _4315 ^ _4318;
  wire _4320 = _4313 ^ _4319;
  wire _4321 = uncoded_block[803] ^ uncoded_block[807];
  wire _4322 = uncoded_block[808] ^ uncoded_block[811];
  wire _4323 = _4321 ^ _4322;
  wire _4324 = uncoded_block[814] ^ uncoded_block[815];
  wire _4325 = uncoded_block[816] ^ uncoded_block[818];
  wire _4326 = _4324 ^ _4325;
  wire _4327 = _4323 ^ _4326;
  wire _4328 = uncoded_block[825] ^ uncoded_block[826];
  wire _4329 = _1242 ^ _4328;
  wire _4330 = uncoded_block[827] ^ uncoded_block[831];
  wire _4331 = uncoded_block[832] ^ uncoded_block[833];
  wire _4332 = _4330 ^ _4331;
  wire _4333 = _4329 ^ _4332;
  wire _4334 = _4327 ^ _4333;
  wire _4335 = _4320 ^ _4334;
  wire _4336 = uncoded_block[834] ^ uncoded_block[836];
  wire _4337 = uncoded_block[838] ^ uncoded_block[839];
  wire _4338 = _4336 ^ _4337;
  wire _4339 = uncoded_block[842] ^ uncoded_block[844];
  wire _4340 = uncoded_block[848] ^ uncoded_block[849];
  wire _4341 = _4339 ^ _4340;
  wire _4342 = _4338 ^ _4341;
  wire _4343 = uncoded_block[853] ^ uncoded_block[857];
  wire _4344 = uncoded_block[860] ^ uncoded_block[865];
  wire _4345 = _4343 ^ _4344;
  wire _4346 = uncoded_block[869] ^ uncoded_block[872];
  wire _4347 = uncoded_block[873] ^ uncoded_block[876];
  wire _4348 = _4346 ^ _4347;
  wire _4349 = _4345 ^ _4348;
  wire _4350 = _4342 ^ _4349;
  wire _4351 = uncoded_block[879] ^ uncoded_block[882];
  wire _4352 = uncoded_block[885] ^ uncoded_block[888];
  wire _4353 = _4351 ^ _4352;
  wire _4354 = uncoded_block[889] ^ uncoded_block[890];
  wire _4355 = uncoded_block[894] ^ uncoded_block[895];
  wire _4356 = _4354 ^ _4355;
  wire _4357 = _4353 ^ _4356;
  wire _4358 = uncoded_block[896] ^ uncoded_block[899];
  wire _4359 = _4358 ^ _429;
  wire _4360 = uncoded_block[903] ^ uncoded_block[907];
  wire _4361 = uncoded_block[908] ^ uncoded_block[912];
  wire _4362 = _4360 ^ _4361;
  wire _4363 = _4359 ^ _4362;
  wire _4364 = _4357 ^ _4363;
  wire _4365 = _4350 ^ _4364;
  wire _4366 = _4335 ^ _4365;
  wire _4367 = uncoded_block[917] ^ uncoded_block[920];
  wire _4368 = uncoded_block[922] ^ uncoded_block[924];
  wire _4369 = _4367 ^ _4368;
  wire _4370 = uncoded_block[925] ^ uncoded_block[927];
  wire _4371 = uncoded_block[928] ^ uncoded_block[929];
  wire _4372 = _4370 ^ _4371;
  wire _4373 = _4369 ^ _4372;
  wire _4374 = uncoded_block[930] ^ uncoded_block[937];
  wire _4375 = uncoded_block[939] ^ uncoded_block[940];
  wire _4376 = _4374 ^ _4375;
  wire _4377 = uncoded_block[941] ^ uncoded_block[943];
  wire _4378 = _4377 ^ _456;
  wire _4379 = _4376 ^ _4378;
  wire _4380 = _4373 ^ _4379;
  wire _4381 = uncoded_block[950] ^ uncoded_block[951];
  wire _4382 = uncoded_block[952] ^ uncoded_block[954];
  wire _4383 = _4381 ^ _4382;
  wire _4384 = uncoded_block[955] ^ uncoded_block[956];
  wire _4385 = uncoded_block[960] ^ uncoded_block[961];
  wire _4386 = _4384 ^ _4385;
  wire _4387 = _4383 ^ _4386;
  wire _4388 = uncoded_block[966] ^ uncoded_block[969];
  wire _4389 = _4388 ^ _468;
  wire _4390 = uncoded_block[973] ^ uncoded_block[975];
  wire _4391 = uncoded_block[976] ^ uncoded_block[978];
  wire _4392 = _4390 ^ _4391;
  wire _4393 = _4389 ^ _4392;
  wire _4394 = _4387 ^ _4393;
  wire _4395 = _4380 ^ _4394;
  wire _4396 = _2100 ^ _476;
  wire _4397 = uncoded_block[983] ^ uncoded_block[986];
  wire _4398 = uncoded_block[987] ^ uncoded_block[991];
  wire _4399 = _4397 ^ _4398;
  wire _4400 = _4396 ^ _4399;
  wire _4401 = uncoded_block[992] ^ uncoded_block[993];
  wire _4402 = uncoded_block[995] ^ uncoded_block[997];
  wire _4403 = _4401 ^ _4402;
  wire _4404 = uncoded_block[1002] ^ uncoded_block[1003];
  wire _4405 = uncoded_block[1007] ^ uncoded_block[1008];
  wire _4406 = _4404 ^ _4405;
  wire _4407 = _4403 ^ _4406;
  wire _4408 = _4400 ^ _4407;
  wire _4409 = uncoded_block[1009] ^ uncoded_block[1010];
  wire _4410 = uncoded_block[1011] ^ uncoded_block[1012];
  wire _4411 = _4409 ^ _4410;
  wire _4412 = uncoded_block[1013] ^ uncoded_block[1016];
  wire _4413 = _4412 ^ _1333;
  wire _4414 = _4411 ^ _4413;
  wire _4415 = uncoded_block[1022] ^ uncoded_block[1026];
  wire _4416 = _4415 ^ _498;
  wire _4417 = uncoded_block[1030] ^ uncoded_block[1031];
  wire _4418 = uncoded_block[1032] ^ uncoded_block[1033];
  wire _4419 = _4417 ^ _4418;
  wire _4420 = _4416 ^ _4419;
  wire _4421 = _4414 ^ _4420;
  wire _4422 = _4408 ^ _4421;
  wire _4423 = _4395 ^ _4422;
  wire _4424 = _4366 ^ _4423;
  wire _4425 = _4307 ^ _4424;
  wire _4426 = _4202 ^ _4425;
  wire _4427 = _2129 ^ _511;
  wire _4428 = _2910 ^ _1356;
  wire _4429 = _4427 ^ _4428;
  wire _4430 = uncoded_block[1054] ^ uncoded_block[1055];
  wire _4431 = uncoded_block[1057] ^ uncoded_block[1059];
  wire _4432 = _4430 ^ _4431;
  wire _4433 = uncoded_block[1060] ^ uncoded_block[1061];
  wire _4434 = uncoded_block[1064] ^ uncoded_block[1075];
  wire _4435 = _4433 ^ _4434;
  wire _4436 = _4432 ^ _4435;
  wire _4437 = _4429 ^ _4436;
  wire _4438 = uncoded_block[1084] ^ uncoded_block[1086];
  wire _4439 = _530 ^ _4438;
  wire _4440 = uncoded_block[1089] ^ uncoded_block[1090];
  wire _4441 = _2149 ^ _4440;
  wire _4442 = _4439 ^ _4441;
  wire _4443 = _1377 ^ _3698;
  wire _4444 = uncoded_block[1100] ^ uncoded_block[1102];
  wire _4445 = _4444 ^ _2160;
  wire _4446 = _4443 ^ _4445;
  wire _4447 = _4442 ^ _4446;
  wire _4448 = _4437 ^ _4447;
  wire _4449 = _2161 ^ _549;
  wire _4450 = uncoded_block[1109] ^ uncoded_block[1110];
  wire _4451 = uncoded_block[1111] ^ uncoded_block[1112];
  wire _4452 = _4450 ^ _4451;
  wire _4453 = _4449 ^ _4452;
  wire _4454 = _2938 ^ _3714;
  wire _4455 = uncoded_block[1121] ^ uncoded_block[1122];
  wire _4456 = _4455 ^ _2172;
  wire _4457 = _4454 ^ _4456;
  wire _4458 = _4453 ^ _4457;
  wire _4459 = uncoded_block[1126] ^ uncoded_block[1127];
  wire _4460 = uncoded_block[1129] ^ uncoded_block[1131];
  wire _4461 = _4459 ^ _4460;
  wire _4462 = uncoded_block[1138] ^ uncoded_block[1140];
  wire _4463 = _2174 ^ _4462;
  wire _4464 = _4461 ^ _4463;
  wire _4465 = uncoded_block[1147] ^ uncoded_block[1148];
  wire _4466 = uncoded_block[1150] ^ uncoded_block[1151];
  wire _4467 = _4465 ^ _4466;
  wire _4468 = uncoded_block[1152] ^ uncoded_block[1153];
  wire _4469 = uncoded_block[1154] ^ uncoded_block[1158];
  wire _4470 = _4468 ^ _4469;
  wire _4471 = _4467 ^ _4470;
  wire _4472 = _4464 ^ _4471;
  wire _4473 = _4458 ^ _4472;
  wire _4474 = _4448 ^ _4473;
  wire _4475 = _3733 ^ _2964;
  wire _4476 = uncoded_block[1167] ^ uncoded_block[1168];
  wire _4477 = _3736 ^ _4476;
  wire _4478 = _4475 ^ _4477;
  wire _4479 = uncoded_block[1171] ^ uncoded_block[1175];
  wire _4480 = _1408 ^ _4479;
  wire _4481 = uncoded_block[1177] ^ uncoded_block[1179];
  wire _4482 = uncoded_block[1180] ^ uncoded_block[1182];
  wire _4483 = _4481 ^ _4482;
  wire _4484 = _4480 ^ _4483;
  wire _4485 = _4478 ^ _4484;
  wire _4486 = uncoded_block[1184] ^ uncoded_block[1185];
  wire _4487 = _4486 ^ _2200;
  wire _4488 = uncoded_block[1192] ^ uncoded_block[1194];
  wire _4489 = _4488 ^ _597;
  wire _4490 = _4487 ^ _4489;
  wire _4491 = uncoded_block[1206] ^ uncoded_block[1208];
  wire _4492 = _2209 ^ _4491;
  wire _4493 = _2208 ^ _4492;
  wire _4494 = _4490 ^ _4493;
  wire _4495 = _4485 ^ _4494;
  wire _4496 = uncoded_block[1212] ^ uncoded_block[1214];
  wire _4497 = _2217 ^ _4496;
  wire _4498 = uncoded_block[1215] ^ uncoded_block[1217];
  wire _4499 = uncoded_block[1218] ^ uncoded_block[1220];
  wire _4500 = _4498 ^ _4499;
  wire _4501 = _4497 ^ _4500;
  wire _4502 = uncoded_block[1221] ^ uncoded_block[1222];
  wire _4503 = _4502 ^ _1435;
  wire _4504 = uncoded_block[1226] ^ uncoded_block[1229];
  wire _4505 = uncoded_block[1230] ^ uncoded_block[1239];
  wire _4506 = _4504 ^ _4505;
  wire _4507 = _4503 ^ _4506;
  wire _4508 = _4501 ^ _4507;
  wire _4509 = uncoded_block[1242] ^ uncoded_block[1243];
  wire _4510 = _4509 ^ _3777;
  wire _4511 = uncoded_block[1248] ^ uncoded_block[1250];
  wire _4512 = _4511 ^ _2235;
  wire _4513 = _4510 ^ _4512;
  wire _4514 = uncoded_block[1259] ^ uncoded_block[1261];
  wire _4515 = _3001 ^ _4514;
  wire _4516 = uncoded_block[1263] ^ uncoded_block[1265];
  wire _4517 = _4516 ^ _2244;
  wire _4518 = _4515 ^ _4517;
  wire _4519 = _4513 ^ _4518;
  wire _4520 = _4508 ^ _4519;
  wire _4521 = _4495 ^ _4520;
  wire _4522 = _4474 ^ _4521;
  wire _4523 = uncoded_block[1273] ^ uncoded_block[1274];
  wire _4524 = _628 ^ _4523;
  wire _4525 = uncoded_block[1281] ^ uncoded_block[1282];
  wire _4526 = uncoded_block[1283] ^ uncoded_block[1287];
  wire _4527 = _4525 ^ _4526;
  wire _4528 = _4524 ^ _4527;
  wire _4529 = uncoded_block[1289] ^ uncoded_block[1290];
  wire _4530 = _4529 ^ _3801;
  wire _4531 = uncoded_block[1296] ^ uncoded_block[1297];
  wire _4532 = uncoded_block[1298] ^ uncoded_block[1299];
  wire _4533 = _4531 ^ _4532;
  wire _4534 = _4530 ^ _4533;
  wire _4535 = _4528 ^ _4534;
  wire _4536 = uncoded_block[1301] ^ uncoded_block[1303];
  wire _4537 = uncoded_block[1305] ^ uncoded_block[1309];
  wire _4538 = _4536 ^ _4537;
  wire _4539 = uncoded_block[1311] ^ uncoded_block[1314];
  wire _4540 = uncoded_block[1318] ^ uncoded_block[1319];
  wire _4541 = _4539 ^ _4540;
  wire _4542 = _4538 ^ _4541;
  wire _4543 = uncoded_block[1323] ^ uncoded_block[1324];
  wire _4544 = _3029 ^ _4543;
  wire _4545 = uncoded_block[1327] ^ uncoded_block[1328];
  wire _4546 = _4545 ^ _1494;
  wire _4547 = _4544 ^ _4546;
  wire _4548 = _4542 ^ _4547;
  wire _4549 = _4535 ^ _4548;
  wire _4550 = uncoded_block[1332] ^ uncoded_block[1333];
  wire _4551 = uncoded_block[1334] ^ uncoded_block[1335];
  wire _4552 = _4550 ^ _4551;
  wire _4553 = uncoded_block[1339] ^ uncoded_block[1340];
  wire _4554 = _2276 ^ _4553;
  wire _4555 = _4552 ^ _4554;
  wire _4556 = uncoded_block[1345] ^ uncoded_block[1346];
  wire _4557 = _4556 ^ _670;
  wire _4558 = uncoded_block[1353] ^ uncoded_block[1356];
  wire _4559 = uncoded_block[1358] ^ uncoded_block[1360];
  wire _4560 = _4558 ^ _4559;
  wire _4561 = _4557 ^ _4560;
  wire _4562 = _4555 ^ _4561;
  wire _4563 = uncoded_block[1369] ^ uncoded_block[1373];
  wire _4564 = uncoded_block[1378] ^ uncoded_block[1381];
  wire _4565 = _4563 ^ _4564;
  wire _4566 = _688 ^ _1513;
  wire _4567 = _4565 ^ _4566;
  wire _4568 = uncoded_block[1391] ^ uncoded_block[1392];
  wire _4569 = uncoded_block[1393] ^ uncoded_block[1394];
  wire _4570 = _4568 ^ _4569;
  wire _4571 = uncoded_block[1395] ^ uncoded_block[1396];
  wire _4572 = uncoded_block[1398] ^ uncoded_block[1399];
  wire _4573 = _4571 ^ _4572;
  wire _4574 = _4570 ^ _4573;
  wire _4575 = _4567 ^ _4574;
  wire _4576 = _4562 ^ _4575;
  wire _4577 = _4549 ^ _4576;
  wire _4578 = uncoded_block[1404] ^ uncoded_block[1405];
  wire _4579 = _3841 ^ _4578;
  wire _4580 = uncoded_block[1411] ^ uncoded_block[1412];
  wire _4581 = _2300 ^ _4580;
  wire _4582 = _4579 ^ _4581;
  wire _4583 = uncoded_block[1414] ^ uncoded_block[1418];
  wire _4584 = uncoded_block[1421] ^ uncoded_block[1424];
  wire _4585 = _4583 ^ _4584;
  wire _4586 = uncoded_block[1432] ^ uncoded_block[1434];
  wire _4587 = _1531 ^ _4586;
  wire _4588 = _4585 ^ _4587;
  wire _4589 = _4582 ^ _4588;
  wire _4590 = uncoded_block[1440] ^ uncoded_block[1441];
  wire _4591 = _3857 ^ _4590;
  wire _4592 = _2321 ^ _3084;
  wire _4593 = _4591 ^ _4592;
  wire _4594 = uncoded_block[1447] ^ uncoded_block[1451];
  wire _4595 = _4594 ^ _719;
  wire _4596 = uncoded_block[1458] ^ uncoded_block[1461];
  wire _4597 = _720 ^ _4596;
  wire _4598 = _4595 ^ _4597;
  wire _4599 = _4593 ^ _4598;
  wire _4600 = _4589 ^ _4599;
  wire _4601 = uncoded_block[1464] ^ uncoded_block[1470];
  wire _4602 = _2336 ^ _4601;
  wire _4603 = uncoded_block[1473] ^ uncoded_block[1474];
  wire _4604 = uncoded_block[1476] ^ uncoded_block[1478];
  wire _4605 = _4603 ^ _4604;
  wire _4606 = _4602 ^ _4605;
  wire _4607 = uncoded_block[1479] ^ uncoded_block[1483];
  wire _4608 = uncoded_block[1484] ^ uncoded_block[1490];
  wire _4609 = _4607 ^ _4608;
  wire _4610 = uncoded_block[1491] ^ uncoded_block[1492];
  wire _4611 = _4610 ^ _2350;
  wire _4612 = _4609 ^ _4611;
  wire _4613 = _4606 ^ _4612;
  wire _4614 = uncoded_block[1502] ^ uncoded_block[1503];
  wire _4615 = _4614 ^ _3894;
  wire _4616 = uncoded_block[1507] ^ uncoded_block[1508];
  wire _4617 = uncoded_block[1509] ^ uncoded_block[1512];
  wire _4618 = _4616 ^ _4617;
  wire _4619 = _4615 ^ _4618;
  wire _4620 = uncoded_block[1517] ^ uncoded_block[1521];
  wire _4621 = uncoded_block[1522] ^ uncoded_block[1525];
  wire _4622 = _4620 ^ _4621;
  wire _4623 = uncoded_block[1526] ^ uncoded_block[1527];
  wire _4624 = uncoded_block[1529] ^ uncoded_block[1532];
  wire _4625 = _4623 ^ _4624;
  wire _4626 = _4622 ^ _4625;
  wire _4627 = _4619 ^ _4626;
  wire _4628 = _4613 ^ _4627;
  wire _4629 = _4600 ^ _4628;
  wire _4630 = _4577 ^ _4629;
  wire _4631 = _4522 ^ _4630;
  wire _4632 = uncoded_block[1535] ^ uncoded_block[1539];
  wire _4633 = _4632 ^ _3909;
  wire _4634 = uncoded_block[1544] ^ uncoded_block[1545];
  wire _4635 = _4634 ^ _2367;
  wire _4636 = _4633 ^ _4635;
  wire _4637 = uncoded_block[1549] ^ uncoded_block[1556];
  wire _4638 = uncoded_block[1558] ^ uncoded_block[1559];
  wire _4639 = _4637 ^ _4638;
  wire _4640 = uncoded_block[1560] ^ uncoded_block[1561];
  wire _4641 = _4640 ^ _2376;
  wire _4642 = _4639 ^ _4641;
  wire _4643 = _4636 ^ _4642;
  wire _4644 = uncoded_block[1566] ^ uncoded_block[1568];
  wire _4645 = uncoded_block[1570] ^ uncoded_block[1572];
  wire _4646 = _4644 ^ _4645;
  wire _4647 = uncoded_block[1573] ^ uncoded_block[1574];
  wire _4648 = uncoded_block[1575] ^ uncoded_block[1576];
  wire _4649 = _4647 ^ _4648;
  wire _4650 = _4646 ^ _4649;
  wire _4651 = uncoded_block[1577] ^ uncoded_block[1579];
  wire _4652 = _4651 ^ _1615;
  wire _4653 = uncoded_block[1590] ^ uncoded_block[1591];
  wire _4654 = uncoded_block[1594] ^ uncoded_block[1595];
  wire _4655 = _4653 ^ _4654;
  wire _4656 = _4652 ^ _4655;
  wire _4657 = _4650 ^ _4656;
  wire _4658 = _4643 ^ _4657;
  wire _4659 = uncoded_block[1598] ^ uncoded_block[1601];
  wire _4660 = uncoded_block[1604] ^ uncoded_block[1607];
  wire _4661 = _4659 ^ _4660;
  wire _4662 = uncoded_block[1610] ^ uncoded_block[1611];
  wire _4663 = _4662 ^ _804;
  wire _4664 = _4661 ^ _4663;
  wire _4665 = uncoded_block[1625] ^ uncoded_block[1627];
  wire _4666 = _3941 ^ _4665;
  wire _4667 = uncoded_block[1629] ^ uncoded_block[1630];
  wire _4668 = uncoded_block[1634] ^ uncoded_block[1637];
  wire _4669 = _4667 ^ _4668;
  wire _4670 = _4666 ^ _4669;
  wire _4671 = _4664 ^ _4670;
  wire _4672 = _3948 ^ _2408;
  wire _4673 = uncoded_block[1643] ^ uncoded_block[1645];
  wire _4674 = uncoded_block[1647] ^ uncoded_block[1650];
  wire _4675 = _4673 ^ _4674;
  wire _4676 = _4672 ^ _4675;
  wire _4677 = uncoded_block[1651] ^ uncoded_block[1652];
  wire _4678 = uncoded_block[1653] ^ uncoded_block[1654];
  wire _4679 = _4677 ^ _4678;
  wire _4680 = uncoded_block[1659] ^ uncoded_block[1660];
  wire _4681 = _3174 ^ _4680;
  wire _4682 = _4679 ^ _4681;
  wire _4683 = _4676 ^ _4682;
  wire _4684 = _4671 ^ _4683;
  wire _4685 = _4658 ^ _4684;
  wire _4686 = _2419 ^ _3179;
  wire _4687 = uncoded_block[1667] ^ uncoded_block[1668];
  wire _4688 = _4687 ^ _3182;
  wire _4689 = _4686 ^ _4688;
  wire _4690 = uncoded_block[1673] ^ uncoded_block[1678];
  wire _4691 = uncoded_block[1681] ^ uncoded_block[1682];
  wire _4692 = _4690 ^ _4691;
  wire _4693 = uncoded_block[1683] ^ uncoded_block[1684];
  wire _4694 = uncoded_block[1685] ^ uncoded_block[1689];
  wire _4695 = _4693 ^ _4694;
  wire _4696 = _4692 ^ _4695;
  wire _4697 = _4689 ^ _4696;
  wire _4698 = uncoded_block[1694] ^ uncoded_block[1701];
  wire _4699 = _839 ^ _4698;
  wire _4700 = uncoded_block[1702] ^ uncoded_block[1703];
  wire _4701 = _4700 ^ _3976;
  wire _4702 = _4699 ^ _4701;
  wire _4703 = uncoded_block[1714] ^ uncoded_block[1720];
  wire _4704 = _4703 ^ uncoded_block[1722];
  wire _4705 = _4702 ^ _4704;
  wire _4706 = _4697 ^ _4705;
  wire _4707 = _4685 ^ _4706;
  wire _4708 = _4631 ^ _4707;
  wire _4709 = _4426 ^ _4708;
  wire _4710 = uncoded_block[0] ^ uncoded_block[2];
  wire _4711 = _4710 ^ _1;
  wire _4712 = uncoded_block[5] ^ uncoded_block[6];
  wire _4713 = uncoded_block[12] ^ uncoded_block[13];
  wire _4714 = _4712 ^ _4713;
  wire _4715 = _4711 ^ _4714;
  wire _4716 = uncoded_block[17] ^ uncoded_block[19];
  wire _4717 = _4716 ^ _3219;
  wire _4718 = uncoded_block[29] ^ uncoded_block[36];
  wire _4719 = _4001 ^ _4718;
  wire _4720 = _4717 ^ _4719;
  wire _4721 = _4715 ^ _4720;
  wire _4722 = _18 ^ _3230;
  wire _4723 = uncoded_block[42] ^ uncoded_block[44];
  wire _4724 = _4723 ^ _885;
  wire _4725 = _4722 ^ _4724;
  wire _4726 = uncoded_block[50] ^ uncoded_block[53];
  wire _4727 = _4726 ^ _2474;
  wire _4728 = uncoded_block[65] ^ uncoded_block[69];
  wire _4729 = _4728 ^ _1711;
  wire _4730 = _4727 ^ _4729;
  wire _4731 = _4725 ^ _4730;
  wire _4732 = _4721 ^ _4731;
  wire _4733 = uncoded_block[73] ^ uncoded_block[74];
  wire _4734 = _4733 ^ _1714;
  wire _4735 = uncoded_block[80] ^ uncoded_block[81];
  wire _4736 = _4735 ^ _41;
  wire _4737 = _4734 ^ _4736;
  wire _4738 = uncoded_block[85] ^ uncoded_block[89];
  wire _4739 = uncoded_block[91] ^ uncoded_block[92];
  wire _4740 = _4738 ^ _4739;
  wire _4741 = uncoded_block[93] ^ uncoded_block[96];
  wire _4742 = _4741 ^ _47;
  wire _4743 = _4740 ^ _4742;
  wire _4744 = _4737 ^ _4743;
  wire _4745 = uncoded_block[99] ^ uncoded_block[100];
  wire _4746 = _4745 ^ _4028;
  wire _4747 = uncoded_block[108] ^ uncoded_block[116];
  wire _4748 = _2490 ^ _4747;
  wire _4749 = _4746 ^ _4748;
  wire _4750 = uncoded_block[118] ^ uncoded_block[119];
  wire _4751 = uncoded_block[122] ^ uncoded_block[124];
  wire _4752 = _4750 ^ _4751;
  wire _4753 = uncoded_block[126] ^ uncoded_block[127];
  wire _4754 = uncoded_block[130] ^ uncoded_block[131];
  wire _4755 = _4753 ^ _4754;
  wire _4756 = _4752 ^ _4755;
  wire _4757 = _4749 ^ _4756;
  wire _4758 = _4744 ^ _4757;
  wire _4759 = _4732 ^ _4758;
  wire _4760 = uncoded_block[137] ^ uncoded_block[138];
  wire _4761 = uncoded_block[142] ^ uncoded_block[147];
  wire _4762 = _4760 ^ _4761;
  wire _4763 = _4762 ^ _1746;
  wire _4764 = uncoded_block[157] ^ uncoded_block[161];
  wire _4765 = _3271 ^ _4764;
  wire _4766 = uncoded_block[173] ^ uncoded_block[178];
  wire _4767 = _1749 ^ _4766;
  wire _4768 = _4765 ^ _4767;
  wire _4769 = _4763 ^ _4768;
  wire _4770 = uncoded_block[179] ^ uncoded_block[181];
  wire _4771 = _4770 ^ _2528;
  wire _4772 = uncoded_block[186] ^ uncoded_block[188];
  wire _4773 = uncoded_block[189] ^ uncoded_block[190];
  wire _4774 = _4772 ^ _4773;
  wire _4775 = _4771 ^ _4774;
  wire _4776 = uncoded_block[192] ^ uncoded_block[193];
  wire _4777 = uncoded_block[195] ^ uncoded_block[200];
  wire _4778 = _4776 ^ _4777;
  wire _4779 = uncoded_block[202] ^ uncoded_block[205];
  wire _4780 = uncoded_block[206] ^ uncoded_block[208];
  wire _4781 = _4779 ^ _4780;
  wire _4782 = _4778 ^ _4781;
  wire _4783 = _4775 ^ _4782;
  wire _4784 = _4769 ^ _4783;
  wire _4785 = uncoded_block[213] ^ uncoded_block[216];
  wire _4786 = _3292 ^ _4785;
  wire _4787 = uncoded_block[218] ^ uncoded_block[219];
  wire _4788 = uncoded_block[221] ^ uncoded_block[222];
  wire _4789 = _4787 ^ _4788;
  wire _4790 = _4786 ^ _4789;
  wire _4791 = uncoded_block[228] ^ uncoded_block[229];
  wire _4792 = _2545 ^ _4791;
  wire _4793 = uncoded_block[234] ^ uncoded_block[238];
  wire _4794 = _2549 ^ _4793;
  wire _4795 = _4792 ^ _4794;
  wire _4796 = _4790 ^ _4795;
  wire _4797 = uncoded_block[243] ^ uncoded_block[244];
  wire _4798 = _112 ^ _4797;
  wire _4799 = uncoded_block[245] ^ uncoded_block[249];
  wire _4800 = uncoded_block[250] ^ uncoded_block[251];
  wire _4801 = _4799 ^ _4800;
  wire _4802 = _4798 ^ _4801;
  wire _4803 = uncoded_block[252] ^ uncoded_block[253];
  wire _4804 = _4803 ^ _119;
  wire _4805 = _4096 ^ _977;
  wire _4806 = _4804 ^ _4805;
  wire _4807 = _4802 ^ _4806;
  wire _4808 = _4796 ^ _4807;
  wire _4809 = _4784 ^ _4808;
  wire _4810 = _4759 ^ _4809;
  wire _4811 = uncoded_block[268] ^ uncoded_block[272];
  wire _4812 = _984 ^ _4811;
  wire _4813 = uncoded_block[273] ^ uncoded_block[276];
  wire _4814 = uncoded_block[277] ^ uncoded_block[279];
  wire _4815 = _4813 ^ _4814;
  wire _4816 = _4812 ^ _4815;
  wire _4817 = uncoded_block[281] ^ uncoded_block[284];
  wire _4818 = _4817 ^ _3327;
  wire _4819 = uncoded_block[292] ^ uncoded_block[293];
  wire _4820 = uncoded_block[294] ^ uncoded_block[295];
  wire _4821 = _4819 ^ _4820;
  wire _4822 = _4818 ^ _4821;
  wire _4823 = _4816 ^ _4822;
  wire _4824 = uncoded_block[300] ^ uncoded_block[302];
  wire _4825 = _1806 ^ _4824;
  wire _4826 = uncoded_block[303] ^ uncoded_block[304];
  wire _4827 = uncoded_block[305] ^ uncoded_block[312];
  wire _4828 = _4826 ^ _4827;
  wire _4829 = _4825 ^ _4828;
  wire _4830 = uncoded_block[317] ^ uncoded_block[318];
  wire _4831 = _146 ^ _4830;
  wire _4832 = uncoded_block[319] ^ uncoded_block[321];
  wire _4833 = _4832 ^ _4123;
  wire _4834 = _4831 ^ _4833;
  wire _4835 = _4829 ^ _4834;
  wire _4836 = _4823 ^ _4835;
  wire _4837 = uncoded_block[328] ^ uncoded_block[331];
  wire _4838 = uncoded_block[332] ^ uncoded_block[335];
  wire _4839 = _4837 ^ _4838;
  wire _4840 = uncoded_block[339] ^ uncoded_block[341];
  wire _4841 = uncoded_block[343] ^ uncoded_block[344];
  wire _4842 = _4840 ^ _4841;
  wire _4843 = _4839 ^ _4842;
  wire _4844 = uncoded_block[346] ^ uncoded_block[347];
  wire _4845 = uncoded_block[348] ^ uncoded_block[351];
  wire _4846 = _4844 ^ _4845;
  wire _4847 = uncoded_block[354] ^ uncoded_block[359];
  wire _4848 = _162 ^ _4847;
  wire _4849 = _4846 ^ _4848;
  wire _4850 = _4843 ^ _4849;
  wire _4851 = uncoded_block[363] ^ uncoded_block[365];
  wire _4852 = _166 ^ _4851;
  wire _4853 = uncoded_block[373] ^ uncoded_block[375];
  wire _4854 = uncoded_block[377] ^ uncoded_block[378];
  wire _4855 = _4853 ^ _4854;
  wire _4856 = _4852 ^ _4855;
  wire _4857 = uncoded_block[380] ^ uncoded_block[382];
  wire _4858 = uncoded_block[383] ^ uncoded_block[385];
  wire _4859 = _4857 ^ _4858;
  wire _4860 = _4149 ^ _2615;
  wire _4861 = _4859 ^ _4860;
  wire _4862 = _4856 ^ _4861;
  wire _4863 = _4850 ^ _4862;
  wire _4864 = _4836 ^ _4863;
  wire _4865 = uncoded_block[400] ^ uncoded_block[403];
  wire _4866 = _180 ^ _4865;
  wire _4867 = uncoded_block[407] ^ uncoded_block[409];
  wire _4868 = uncoded_block[411] ^ uncoded_block[413];
  wire _4869 = _4867 ^ _4868;
  wire _4870 = _4866 ^ _4869;
  wire _4871 = uncoded_block[415] ^ uncoded_block[417];
  wire _4872 = uncoded_block[419] ^ uncoded_block[420];
  wire _4873 = _4871 ^ _4872;
  wire _4874 = uncoded_block[422] ^ uncoded_block[424];
  wire _4875 = _4874 ^ _197;
  wire _4876 = _4873 ^ _4875;
  wire _4877 = _4870 ^ _4876;
  wire _4878 = uncoded_block[428] ^ uncoded_block[435];
  wire _4879 = _4878 ^ _3404;
  wire _4880 = _3405 ^ _205;
  wire _4881 = _4879 ^ _4880;
  wire _4882 = uncoded_block[443] ^ uncoded_block[449];
  wire _4883 = uncoded_block[450] ^ uncoded_block[451];
  wire _4884 = _4882 ^ _4883;
  wire _4885 = uncoded_block[457] ^ uncoded_block[460];
  wire _4886 = _212 ^ _4885;
  wire _4887 = _4884 ^ _4886;
  wire _4888 = _4881 ^ _4887;
  wire _4889 = _4877 ^ _4888;
  wire _4890 = uncoded_block[464] ^ uncoded_block[465];
  wire _4891 = _4181 ^ _4890;
  wire _4892 = _4186 ^ _1082;
  wire _4893 = _4891 ^ _4892;
  wire _4894 = uncoded_block[473] ^ uncoded_block[480];
  wire _4895 = uncoded_block[481] ^ uncoded_block[482];
  wire _4896 = _4894 ^ _4895;
  wire _4897 = uncoded_block[484] ^ uncoded_block[485];
  wire _4898 = uncoded_block[487] ^ uncoded_block[490];
  wire _4899 = _4897 ^ _4898;
  wire _4900 = _4896 ^ _4899;
  wire _4901 = _4893 ^ _4900;
  wire _4902 = uncoded_block[491] ^ uncoded_block[493];
  wire _4903 = uncoded_block[494] ^ uncoded_block[497];
  wire _4904 = _4902 ^ _4903;
  wire _4905 = uncoded_block[498] ^ uncoded_block[499];
  wire _4906 = _4905 ^ _2668;
  wire _4907 = _4904 ^ _4906;
  wire _4908 = uncoded_block[510] ^ uncoded_block[511];
  wire _4909 = _4908 ^ _3439;
  wire _4910 = uncoded_block[516] ^ uncoded_block[517];
  wire _4911 = _232 ^ _4910;
  wire _4912 = _4909 ^ _4911;
  wire _4913 = _4907 ^ _4912;
  wire _4914 = _4901 ^ _4913;
  wire _4915 = _4889 ^ _4914;
  wire _4916 = _4864 ^ _4915;
  wire _4917 = _4810 ^ _4916;
  wire _4918 = uncoded_block[518] ^ uncoded_block[520];
  wire _4919 = uncoded_block[521] ^ uncoded_block[524];
  wire _4920 = _4918 ^ _4919;
  wire _4921 = uncoded_block[525] ^ uncoded_block[526];
  wire _4922 = uncoded_block[527] ^ uncoded_block[528];
  wire _4923 = _4921 ^ _4922;
  wire _4924 = _4920 ^ _4923;
  wire _4925 = uncoded_block[529] ^ uncoded_block[530];
  wire _4926 = uncoded_block[532] ^ uncoded_block[535];
  wire _4927 = _4925 ^ _4926;
  wire _4928 = _3451 ^ _4217;
  wire _4929 = _4927 ^ _4928;
  wire _4930 = _4924 ^ _4929;
  wire _4931 = uncoded_block[546] ^ uncoded_block[548];
  wire _4932 = _244 ^ _4931;
  wire _4933 = uncoded_block[549] ^ uncoded_block[550];
  wire _4934 = uncoded_block[553] ^ uncoded_block[557];
  wire _4935 = _4933 ^ _4934;
  wire _4936 = _4932 ^ _4935;
  wire _4937 = uncoded_block[558] ^ uncoded_block[559];
  wire _4938 = uncoded_block[560] ^ uncoded_block[561];
  wire _4939 = _4937 ^ _4938;
  wire _4940 = uncoded_block[563] ^ uncoded_block[569];
  wire _4941 = uncoded_block[574] ^ uncoded_block[575];
  wire _4942 = _4940 ^ _4941;
  wire _4943 = _4939 ^ _4942;
  wire _4944 = _4936 ^ _4943;
  wire _4945 = _4930 ^ _4944;
  wire _4946 = uncoded_block[581] ^ uncoded_block[582];
  wire _4947 = uncoded_block[585] ^ uncoded_block[587];
  wire _4948 = _4946 ^ _4947;
  wire _4949 = _1134 ^ _4948;
  wire _4950 = uncoded_block[588] ^ uncoded_block[589];
  wire _4951 = _4950 ^ _4234;
  wire _4952 = uncoded_block[596] ^ uncoded_block[598];
  wire _4953 = uncoded_block[599] ^ uncoded_block[600];
  wire _4954 = _4952 ^ _4953;
  wire _4955 = _4951 ^ _4954;
  wire _4956 = _4949 ^ _4955;
  wire _4957 = uncoded_block[604] ^ uncoded_block[607];
  wire _4958 = _3487 ^ _4957;
  wire _4959 = uncoded_block[610] ^ uncoded_block[615];
  wire _4960 = uncoded_block[618] ^ uncoded_block[620];
  wire _4961 = _4959 ^ _4960;
  wire _4962 = _4958 ^ _4961;
  wire _4963 = uncoded_block[622] ^ uncoded_block[623];
  wire _4964 = uncoded_block[625] ^ uncoded_block[626];
  wire _4965 = _4963 ^ _4964;
  wire _4966 = _289 ^ _3501;
  wire _4967 = _4965 ^ _4966;
  wire _4968 = _4962 ^ _4967;
  wire _4969 = _4956 ^ _4968;
  wire _4970 = _4945 ^ _4969;
  wire _4971 = _293 ^ _2727;
  wire _4972 = uncoded_block[643] ^ uncoded_block[644];
  wire _4973 = _4972 ^ _1957;
  wire _4974 = _4971 ^ _4973;
  wire _4975 = uncoded_block[653] ^ uncoded_block[654];
  wire _4976 = _1960 ^ _4975;
  wire _4977 = uncoded_block[657] ^ uncoded_block[661];
  wire _4978 = uncoded_block[664] ^ uncoded_block[665];
  wire _4979 = _4977 ^ _4978;
  wire _4980 = _4976 ^ _4979;
  wire _4981 = _4974 ^ _4980;
  wire _4982 = uncoded_block[668] ^ uncoded_block[673];
  wire _4983 = _4982 ^ _1180;
  wire _4984 = uncoded_block[683] ^ uncoded_block[689];
  wire _4985 = _1971 ^ _4984;
  wire _4986 = _4983 ^ _4985;
  wire _4987 = uncoded_block[694] ^ uncoded_block[696];
  wire _4988 = _1186 ^ _4987;
  wire _4989 = uncoded_block[698] ^ uncoded_block[700];
  wire _4990 = uncoded_block[701] ^ uncoded_block[703];
  wire _4991 = _4989 ^ _4990;
  wire _4992 = _4988 ^ _4991;
  wire _4993 = _4986 ^ _4992;
  wire _4994 = _4981 ^ _4993;
  wire _4995 = uncoded_block[706] ^ uncoded_block[707];
  wire _4996 = uncoded_block[709] ^ uncoded_block[710];
  wire _4997 = _4995 ^ _4996;
  wire _4998 = uncoded_block[711] ^ uncoded_block[714];
  wire _4999 = uncoded_block[715] ^ uncoded_block[716];
  wire _5000 = _4998 ^ _4999;
  wire _5001 = _4997 ^ _5000;
  wire _5002 = uncoded_block[717] ^ uncoded_block[718];
  wire _5003 = uncoded_block[724] ^ uncoded_block[728];
  wire _5004 = _5002 ^ _5003;
  wire _5005 = uncoded_block[730] ^ uncoded_block[732];
  wire _5006 = uncoded_block[733] ^ uncoded_block[735];
  wire _5007 = _5005 ^ _5006;
  wire _5008 = _5004 ^ _5007;
  wire _5009 = _5001 ^ _5008;
  wire _5010 = uncoded_block[741] ^ uncoded_block[742];
  wire _5011 = _350 ^ _5010;
  wire _5012 = uncoded_block[745] ^ uncoded_block[746];
  wire _5013 = uncoded_block[747] ^ uncoded_block[748];
  wire _5014 = _5012 ^ _5013;
  wire _5015 = _5011 ^ _5014;
  wire _5016 = uncoded_block[751] ^ uncoded_block[753];
  wire _5017 = uncoded_block[754] ^ uncoded_block[757];
  wire _5018 = _5016 ^ _5017;
  wire _5019 = uncoded_block[759] ^ uncoded_block[762];
  wire _5020 = uncoded_block[763] ^ uncoded_block[766];
  wire _5021 = _5019 ^ _5020;
  wire _5022 = _5018 ^ _5021;
  wire _5023 = _5015 ^ _5022;
  wire _5024 = _5009 ^ _5023;
  wire _5025 = _4994 ^ _5024;
  wire _5026 = _4970 ^ _5025;
  wire _5027 = uncoded_block[768] ^ uncoded_block[769];
  wire _5028 = _5027 ^ _2791;
  wire _5029 = uncoded_block[780] ^ uncoded_block[784];
  wire _5030 = _2014 ^ _5029;
  wire _5031 = _5028 ^ _5030;
  wire _5032 = uncoded_block[787] ^ uncoded_block[788];
  wire _5033 = uncoded_block[789] ^ uncoded_block[790];
  wire _5034 = _5032 ^ _5033;
  wire _5035 = uncoded_block[795] ^ uncoded_block[798];
  wire _5036 = _1232 ^ _5035;
  wire _5037 = _5034 ^ _5036;
  wire _5038 = _5031 ^ _5037;
  wire _5039 = uncoded_block[800] ^ uncoded_block[802];
  wire _5040 = _5039 ^ _1235;
  wire _5041 = uncoded_block[808] ^ uncoded_block[809];
  wire _5042 = uncoded_block[810] ^ uncoded_block[811];
  wire _5043 = _5041 ^ _5042;
  wire _5044 = _5040 ^ _5043;
  wire _5045 = uncoded_block[813] ^ uncoded_block[815];
  wire _5046 = uncoded_block[816] ^ uncoded_block[817];
  wire _5047 = _5045 ^ _5046;
  wire _5048 = _5047 ^ _2030;
  wire _5049 = _5044 ^ _5048;
  wire _5050 = _5038 ^ _5049;
  wire _5051 = uncoded_block[822] ^ uncoded_block[824];
  wire _5052 = uncoded_block[827] ^ uncoded_block[830];
  wire _5053 = _5051 ^ _5052;
  wire _5054 = uncoded_block[835] ^ uncoded_block[838];
  wire _5055 = _2033 ^ _5054;
  wire _5056 = _5053 ^ _5055;
  wire _5057 = uncoded_block[840] ^ uncoded_block[841];
  wire _5058 = uncoded_block[842] ^ uncoded_block[843];
  wire _5059 = _5057 ^ _5058;
  wire _5060 = uncoded_block[844] ^ uncoded_block[846];
  wire _5061 = _5060 ^ _3599;
  wire _5062 = _5059 ^ _5061;
  wire _5063 = _5056 ^ _5062;
  wire _5064 = uncoded_block[849] ^ uncoded_block[853];
  wire _5065 = _5064 ^ _3600;
  wire _5066 = uncoded_block[858] ^ uncoded_block[859];
  wire _5067 = _5066 ^ _3603;
  wire _5068 = _5065 ^ _5067;
  wire _5069 = uncoded_block[864] ^ uncoded_block[865];
  wire _5070 = _413 ^ _5069;
  wire _5071 = uncoded_block[866] ^ uncoded_block[867];
  wire _5072 = uncoded_block[869] ^ uncoded_block[870];
  wire _5073 = _5071 ^ _5072;
  wire _5074 = _5070 ^ _5073;
  wire _5075 = _5068 ^ _5074;
  wire _5076 = _5063 ^ _5075;
  wire _5077 = _5050 ^ _5076;
  wire _5078 = uncoded_block[876] ^ uncoded_block[878];
  wire _5079 = uncoded_block[880] ^ uncoded_block[881];
  wire _5080 = _5078 ^ _5079;
  wire _5081 = _418 ^ _5080;
  wire _5082 = uncoded_block[886] ^ uncoded_block[888];
  wire _5083 = uncoded_block[893] ^ uncoded_block[894];
  wire _5084 = _5082 ^ _5083;
  wire _5085 = uncoded_block[895] ^ uncoded_block[896];
  wire _5086 = _5085 ^ _428;
  wire _5087 = _5084 ^ _5086;
  wire _5088 = _5081 ^ _5087;
  wire _5089 = uncoded_block[899] ^ uncoded_block[902];
  wire _5090 = uncoded_block[903] ^ uncoded_block[909];
  wire _5091 = _5089 ^ _5090;
  wire _5092 = uncoded_block[914] ^ uncoded_block[917];
  wire _5093 = _435 ^ _5092;
  wire _5094 = _5091 ^ _5093;
  wire _5095 = _445 ^ _2857;
  wire _5096 = uncoded_block[931] ^ uncoded_block[932];
  wire _5097 = _5096 ^ _2079;
  wire _5098 = _5095 ^ _5097;
  wire _5099 = _5094 ^ _5098;
  wire _5100 = _5088 ^ _5099;
  wire _5101 = uncoded_block[936] ^ uncoded_block[937];
  wire _5102 = _5101 ^ _4375;
  wire _5103 = _5102 ^ _457;
  wire _5104 = uncoded_block[948] ^ uncoded_block[953];
  wire _5105 = uncoded_block[955] ^ uncoded_block[959];
  wire _5106 = _5104 ^ _5105;
  wire _5107 = uncoded_block[960] ^ uncoded_block[962];
  wire _5108 = uncoded_block[964] ^ uncoded_block[969];
  wire _5109 = _5107 ^ _5108;
  wire _5110 = _5106 ^ _5109;
  wire _5111 = _5103 ^ _5110;
  wire _5112 = uncoded_block[973] ^ uncoded_block[974];
  wire _5113 = _1314 ^ _5112;
  wire _5114 = uncoded_block[976] ^ uncoded_block[977];
  wire _5115 = uncoded_block[978] ^ uncoded_block[984];
  wire _5116 = _5114 ^ _5115;
  wire _5117 = _5113 ^ _5116;
  wire _5118 = uncoded_block[985] ^ uncoded_block[988];
  wire _5119 = uncoded_block[989] ^ uncoded_block[995];
  wire _5120 = _5118 ^ _5119;
  wire _5121 = _480 ^ _4404;
  wire _5122 = _5120 ^ _5121;
  wire _5123 = _5117 ^ _5122;
  wire _5124 = _5111 ^ _5123;
  wire _5125 = _5100 ^ _5124;
  wire _5126 = _5077 ^ _5125;
  wire _5127 = _5026 ^ _5126;
  wire _5128 = _4917 ^ _5127;
  wire _5129 = uncoded_block[1008] ^ uncoded_block[1009];
  wire _5130 = _2114 ^ _5129;
  wire _5131 = uncoded_block[1013] ^ uncoded_block[1015];
  wire _5132 = _4410 ^ _5131;
  wire _5133 = _5130 ^ _5132;
  wire _5134 = uncoded_block[1016] ^ uncoded_block[1017];
  wire _5135 = uncoded_block[1019] ^ uncoded_block[1021];
  wire _5136 = _5134 ^ _5135;
  wire _5137 = uncoded_block[1022] ^ uncoded_block[1023];
  wire _5138 = uncoded_block[1024] ^ uncoded_block[1028];
  wire _5139 = _5137 ^ _5138;
  wire _5140 = _5136 ^ _5139;
  wire _5141 = _5133 ^ _5140;
  wire _5142 = _2898 ^ _2127;
  wire _5143 = uncoded_block[1038] ^ uncoded_block[1040];
  wire _5144 = _1342 ^ _5143;
  wire _5145 = _5142 ^ _5144;
  wire _5146 = _512 ^ _3681;
  wire _5147 = uncoded_block[1051] ^ uncoded_block[1053];
  wire _5148 = _1357 ^ _5147;
  wire _5149 = _5146 ^ _5148;
  wire _5150 = _5145 ^ _5149;
  wire _5151 = _5141 ^ _5150;
  wire _5152 = _4430 ^ _519;
  wire _5153 = uncoded_block[1061] ^ uncoded_block[1064];
  wire _5154 = _1363 ^ _5153;
  wire _5155 = _5152 ^ _5154;
  wire _5156 = uncoded_block[1069] ^ uncoded_block[1071];
  wire _5157 = _2921 ^ _5156;
  wire _5158 = uncoded_block[1072] ^ uncoded_block[1073];
  wire _5159 = _5158 ^ _2924;
  wire _5160 = _5157 ^ _5159;
  wire _5161 = _5155 ^ _5160;
  wire _5162 = uncoded_block[1078] ^ uncoded_block[1079];
  wire _5163 = uncoded_block[1080] ^ uncoded_block[1083];
  wire _5164 = _5162 ^ _5163;
  wire _5165 = uncoded_block[1085] ^ uncoded_block[1093];
  wire _5166 = uncoded_block[1094] ^ uncoded_block[1097];
  wire _5167 = _5165 ^ _5166;
  wire _5168 = _5164 ^ _5167;
  wire _5169 = uncoded_block[1099] ^ uncoded_block[1100];
  wire _5170 = _5169 ^ _2161;
  wire _5171 = _5170 ^ _2166;
  wire _5172 = _5168 ^ _5171;
  wire _5173 = _5161 ^ _5172;
  wire _5174 = _5151 ^ _5173;
  wire _5175 = uncoded_block[1116] ^ uncoded_block[1118];
  wire _5176 = uncoded_block[1121] ^ uncoded_block[1123];
  wire _5177 = _5175 ^ _5176;
  wire _5178 = uncoded_block[1124] ^ uncoded_block[1130];
  wire _5179 = _5178 ^ _1393;
  wire _5180 = _5177 ^ _5179;
  wire _5181 = uncoded_block[1135] ^ uncoded_block[1138];
  wire _5182 = uncoded_block[1139] ^ uncoded_block[1141];
  wire _5183 = _5181 ^ _5182;
  wire _5184 = uncoded_block[1146] ^ uncoded_block[1149];
  wire _5185 = _1400 ^ _5184;
  wire _5186 = _5183 ^ _5185;
  wire _5187 = _5180 ^ _5186;
  wire _5188 = uncoded_block[1154] ^ uncoded_block[1156];
  wire _5189 = _4468 ^ _5188;
  wire _5190 = uncoded_block[1157] ^ uncoded_block[1158];
  wire _5191 = _5190 ^ _3733;
  wire _5192 = _5189 ^ _5191;
  wire _5193 = uncoded_block[1166] ^ uncoded_block[1167];
  wire _5194 = _1407 ^ _5193;
  wire _5195 = uncoded_block[1175] ^ uncoded_block[1178];
  wire _5196 = _5195 ^ _590;
  wire _5197 = _5194 ^ _5196;
  wire _5198 = _5192 ^ _5197;
  wire _5199 = _5187 ^ _5198;
  wire _5200 = uncoded_block[1183] ^ uncoded_block[1184];
  wire _5201 = uncoded_block[1186] ^ uncoded_block[1187];
  wire _5202 = _5200 ^ _5201;
  wire _5203 = uncoded_block[1189] ^ uncoded_block[1191];
  wire _5204 = _5203 ^ _1420;
  wire _5205 = _5202 ^ _5204;
  wire _5206 = uncoded_block[1197] ^ uncoded_block[1201];
  wire _5207 = uncoded_block[1202] ^ uncoded_block[1205];
  wire _5208 = _5206 ^ _5207;
  wire _5209 = uncoded_block[1208] ^ uncoded_block[1209];
  wire _5210 = _5209 ^ _1427;
  wire _5211 = _5208 ^ _5210;
  wire _5212 = _5205 ^ _5211;
  wire _5213 = uncoded_block[1212] ^ uncoded_block[1216];
  wire _5214 = _5213 ^ _2220;
  wire _5215 = uncoded_block[1220] ^ uncoded_block[1221];
  wire _5216 = _5215 ^ _1435;
  wire _5217 = _5214 ^ _5216;
  wire _5218 = uncoded_block[1229] ^ uncoded_block[1231];
  wire _5219 = uncoded_block[1233] ^ uncoded_block[1234];
  wire _5220 = _5218 ^ _5219;
  wire _5221 = uncoded_block[1238] ^ uncoded_block[1239];
  wire _5222 = _2989 ^ _5221;
  wire _5223 = _5220 ^ _5222;
  wire _5224 = _5217 ^ _5223;
  wire _5225 = _5212 ^ _5224;
  wire _5226 = _5199 ^ _5225;
  wire _5227 = _5174 ^ _5226;
  wire _5228 = uncoded_block[1240] ^ uncoded_block[1245];
  wire _5229 = uncoded_block[1247] ^ uncoded_block[1249];
  wire _5230 = _5228 ^ _5229;
  wire _5231 = uncoded_block[1252] ^ uncoded_block[1253];
  wire _5232 = _5231 ^ _3001;
  wire _5233 = _5230 ^ _5232;
  wire _5234 = uncoded_block[1258] ^ uncoded_block[1259];
  wire _5235 = uncoded_block[1262] ^ uncoded_block[1263];
  wire _5236 = _5234 ^ _5235;
  wire _5237 = uncoded_block[1265] ^ uncoded_block[1270];
  wire _5238 = _5237 ^ _1463;
  wire _5239 = _5236 ^ _5238;
  wire _5240 = _5233 ^ _5239;
  wire _5241 = uncoded_block[1278] ^ uncoded_block[1282];
  wire _5242 = _5241 ^ _638;
  wire _5243 = uncoded_block[1285] ^ uncoded_block[1286];
  wire _5244 = _5243 ^ _1468;
  wire _5245 = _5242 ^ _5244;
  wire _5246 = uncoded_block[1297] ^ uncoded_block[1300];
  wire _5247 = _3015 ^ _5246;
  wire _5248 = uncoded_block[1301] ^ uncoded_block[1308];
  wire _5249 = _5248 ^ _2261;
  wire _5250 = _5247 ^ _5249;
  wire _5251 = _5245 ^ _5250;
  wire _5252 = _5240 ^ _5251;
  wire _5253 = uncoded_block[1315] ^ uncoded_block[1318];
  wire _5254 = uncoded_block[1320] ^ uncoded_block[1322];
  wire _5255 = _5253 ^ _5254;
  wire _5256 = uncoded_block[1330] ^ uncoded_block[1333];
  wire _5257 = _1490 ^ _5256;
  wire _5258 = _5255 ^ _5257;
  wire _5259 = uncoded_block[1336] ^ uncoded_block[1337];
  wire _5260 = _4551 ^ _5259;
  wire _5261 = uncoded_block[1338] ^ uncoded_block[1340];
  wire _5262 = uncoded_block[1341] ^ uncoded_block[1342];
  wire _5263 = _5261 ^ _5262;
  wire _5264 = _5260 ^ _5263;
  wire _5265 = _5258 ^ _5264;
  wire _5266 = uncoded_block[1343] ^ uncoded_block[1344];
  wire _5267 = _5266 ^ _4556;
  wire _5268 = uncoded_block[1347] ^ uncoded_block[1348];
  wire _5269 = uncoded_block[1349] ^ uncoded_block[1350];
  wire _5270 = _5268 ^ _5269;
  wire _5271 = _5267 ^ _5270;
  wire _5272 = uncoded_block[1354] ^ uncoded_block[1355];
  wire _5273 = uncoded_block[1358] ^ uncoded_block[1359];
  wire _5274 = _5272 ^ _5273;
  wire _5275 = uncoded_block[1361] ^ uncoded_block[1362];
  wire _5276 = _5275 ^ _2283;
  wire _5277 = _5274 ^ _5276;
  wire _5278 = _5271 ^ _5277;
  wire _5279 = _5265 ^ _5278;
  wire _5280 = _5252 ^ _5279;
  wire _5281 = uncoded_block[1367] ^ uncoded_block[1369];
  wire _5282 = uncoded_block[1370] ^ uncoded_block[1375];
  wire _5283 = _5281 ^ _5282;
  wire _5284 = uncoded_block[1376] ^ uncoded_block[1377];
  wire _5285 = uncoded_block[1378] ^ uncoded_block[1380];
  wire _5286 = _5284 ^ _5285;
  wire _5287 = _5283 ^ _5286;
  wire _5288 = uncoded_block[1383] ^ uncoded_block[1387];
  wire _5289 = _5288 ^ _691;
  wire _5290 = _4569 ^ _3065;
  wire _5291 = _5289 ^ _5290;
  wire _5292 = _5287 ^ _5291;
  wire _5293 = uncoded_block[1401] ^ uncoded_block[1402];
  wire _5294 = uncoded_block[1407] ^ uncoded_block[1411];
  wire _5295 = _5293 ^ _5294;
  wire _5296 = uncoded_block[1412] ^ uncoded_block[1416];
  wire _5297 = _5296 ^ _705;
  wire _5298 = _5295 ^ _5297;
  wire _5299 = uncoded_block[1430] ^ uncoded_block[1432];
  wire _5300 = _1530 ^ _5299;
  wire _5301 = _1528 ^ _5300;
  wire _5302 = _5298 ^ _5301;
  wire _5303 = _5292 ^ _5302;
  wire _5304 = uncoded_block[1440] ^ uncoded_block[1442];
  wire _5305 = uncoded_block[1444] ^ uncoded_block[1445];
  wire _5306 = _5304 ^ _5305;
  wire _5307 = _2315 ^ _5306;
  wire _5308 = _3864 ^ _2328;
  wire _5309 = uncoded_block[1455] ^ uncoded_block[1456];
  wire _5310 = _5309 ^ _723;
  wire _5311 = _5308 ^ _5310;
  wire _5312 = _5307 ^ _5311;
  wire _5313 = uncoded_block[1459] ^ uncoded_block[1463];
  wire _5314 = uncoded_block[1465] ^ uncoded_block[1468];
  wire _5315 = _5313 ^ _5314;
  wire _5316 = uncoded_block[1474] ^ uncoded_block[1476];
  wire _5317 = _732 ^ _5316;
  wire _5318 = _5315 ^ _5317;
  wire _5319 = _2342 ^ _2344;
  wire _5320 = uncoded_block[1483] ^ uncoded_block[1484];
  wire _5321 = uncoded_block[1485] ^ uncoded_block[1488];
  wire _5322 = _5320 ^ _5321;
  wire _5323 = _5319 ^ _5322;
  wire _5324 = _5318 ^ _5323;
  wire _5325 = _5312 ^ _5324;
  wire _5326 = _5303 ^ _5325;
  wire _5327 = _5280 ^ _5326;
  wire _5328 = _5227 ^ _5327;
  wire _5329 = uncoded_block[1491] ^ uncoded_block[1493];
  wire _5330 = _5329 ^ _3890;
  wire _5331 = _4614 ^ _3112;
  wire _5332 = _5330 ^ _5331;
  wire _5333 = uncoded_block[1508] ^ uncoded_block[1509];
  wire _5334 = uncoded_block[1510] ^ uncoded_block[1511];
  wire _5335 = _5333 ^ _5334;
  wire _5336 = uncoded_block[1513] ^ uncoded_block[1515];
  wire _5337 = uncoded_block[1516] ^ uncoded_block[1517];
  wire _5338 = _5336 ^ _5337;
  wire _5339 = _5335 ^ _5338;
  wire _5340 = _5332 ^ _5339;
  wire _5341 = uncoded_block[1519] ^ uncoded_block[1522];
  wire _5342 = _5341 ^ _3118;
  wire _5343 = uncoded_block[1527] ^ uncoded_block[1528];
  wire _5344 = uncoded_block[1529] ^ uncoded_block[1531];
  wire _5345 = _5343 ^ _5344;
  wire _5346 = _5342 ^ _5345;
  wire _5347 = uncoded_block[1534] ^ uncoded_block[1535];
  wire _5348 = uncoded_block[1536] ^ uncoded_block[1539];
  wire _5349 = _5347 ^ _5348;
  wire _5350 = uncoded_block[1540] ^ uncoded_block[1541];
  wire _5351 = _5350 ^ _1590;
  wire _5352 = _5349 ^ _5351;
  wire _5353 = _5346 ^ _5352;
  wire _5354 = _5340 ^ _5353;
  wire _5355 = uncoded_block[1545] ^ uncoded_block[1546];
  wire _5356 = uncoded_block[1547] ^ uncoded_block[1551];
  wire _5357 = _5355 ^ _5356;
  wire _5358 = uncoded_block[1553] ^ uncoded_block[1555];
  wire _5359 = _5358 ^ _1596;
  wire _5360 = _5357 ^ _5359;
  wire _5361 = uncoded_block[1563] ^ uncoded_block[1564];
  wire _5362 = _5361 ^ _1606;
  wire _5363 = uncoded_block[1570] ^ uncoded_block[1571];
  wire _5364 = _5363 ^ _781;
  wire _5365 = _5362 ^ _5364;
  wire _5366 = _5360 ^ _5365;
  wire _5367 = _782 ^ _2383;
  wire _5368 = uncoded_block[1587] ^ uncoded_block[1588];
  wire _5369 = _3925 ^ _5368;
  wire _5370 = _5367 ^ _5369;
  wire _5371 = uncoded_block[1589] ^ uncoded_block[1592];
  wire _5372 = _5371 ^ _4654;
  wire _5373 = uncoded_block[1599] ^ uncoded_block[1601];
  wire _5374 = _1620 ^ _5373;
  wire _5375 = _5372 ^ _5374;
  wire _5376 = _5370 ^ _5375;
  wire _5377 = _5366 ^ _5376;
  wire _5378 = _5354 ^ _5377;
  wire _5379 = uncoded_block[1602] ^ uncoded_block[1608];
  wire _5380 = uncoded_block[1609] ^ uncoded_block[1610];
  wire _5381 = _5379 ^ _5380;
  wire _5382 = uncoded_block[1612] ^ uncoded_block[1615];
  wire _5383 = uncoded_block[1616] ^ uncoded_block[1620];
  wire _5384 = _5382 ^ _5383;
  wire _5385 = _5381 ^ _5384;
  wire _5386 = uncoded_block[1624] ^ uncoded_block[1627];
  wire _5387 = _5386 ^ _808;
  wire _5388 = uncoded_block[1631] ^ uncoded_block[1632];
  wire _5389 = _5388 ^ _1641;
  wire _5390 = _5387 ^ _5389;
  wire _5391 = _5385 ^ _5390;
  wire _5392 = uncoded_block[1637] ^ uncoded_block[1639];
  wire _5393 = _5392 ^ _1646;
  wire _5394 = uncoded_block[1644] ^ uncoded_block[1645];
  wire _5395 = uncoded_block[1646] ^ uncoded_block[1651];
  wire _5396 = _5394 ^ _5395;
  wire _5397 = _5393 ^ _5396;
  wire _5398 = uncoded_block[1656] ^ uncoded_block[1661];
  wire _5399 = uncoded_block[1666] ^ uncoded_block[1667];
  wire _5400 = _5398 ^ _5399;
  wire _5401 = uncoded_block[1675] ^ uncoded_block[1677];
  wire _5402 = _2423 ^ _5401;
  wire _5403 = _5400 ^ _5402;
  wire _5404 = _5397 ^ _5403;
  wire _5405 = _5391 ^ _5404;
  wire _5406 = uncoded_block[1678] ^ uncoded_block[1681];
  wire _5407 = uncoded_block[1683] ^ uncoded_block[1688];
  wire _5408 = _5406 ^ _5407;
  wire _5409 = uncoded_block[1697] ^ uncoded_block[1698];
  wire _5410 = _3967 ^ _5409;
  wire _5411 = _5408 ^ _5410;
  wire _5412 = uncoded_block[1705] ^ uncoded_block[1708];
  wire _5413 = _3973 ^ _5412;
  wire _5414 = _5413 ^ _3201;
  wire _5415 = _5411 ^ _5414;
  wire _5416 = _860 ^ uncoded_block[1722];
  wire _5417 = _5415 ^ _5416;
  wire _5418 = _5405 ^ _5417;
  wire _5419 = _5378 ^ _5418;
  wire _5420 = _5328 ^ _5419;
  wire _5421 = _5128 ^ _5420;
  wire _5422 = _1 ^ _3993;
  wire _5423 = uncoded_block[15] ^ uncoded_block[16];
  wire _5424 = _4713 ^ _5423;
  wire _5425 = _5422 ^ _5424;
  wire _5426 = uncoded_block[18] ^ uncoded_block[22];
  wire _5427 = uncoded_block[24] ^ uncoded_block[28];
  wire _5428 = _5426 ^ _5427;
  wire _5429 = uncoded_block[29] ^ uncoded_block[32];
  wire _5430 = _5429 ^ _880;
  wire _5431 = _5428 ^ _5430;
  wire _5432 = _5425 ^ _5431;
  wire _5433 = uncoded_block[47] ^ uncoded_block[50];
  wire _5434 = _4009 ^ _5433;
  wire _5435 = uncoded_block[51] ^ uncoded_block[52];
  wire _5436 = uncoded_block[54] ^ uncoded_block[55];
  wire _5437 = _5435 ^ _5436;
  wire _5438 = _5434 ^ _5437;
  wire _5439 = uncoded_block[57] ^ uncoded_block[65];
  wire _5440 = uncoded_block[68] ^ uncoded_block[70];
  wire _5441 = _5439 ^ _5440;
  wire _5442 = uncoded_block[71] ^ uncoded_block[73];
  wire _5443 = uncoded_block[75] ^ uncoded_block[77];
  wire _5444 = _5442 ^ _5443;
  wire _5445 = _5441 ^ _5444;
  wire _5446 = _5438 ^ _5445;
  wire _5447 = _5432 ^ _5446;
  wire _5448 = _4735 ^ _903;
  wire _5449 = uncoded_block[97] ^ uncoded_block[102];
  wire _5450 = _4026 ^ _5449;
  wire _5451 = _5448 ^ _5450;
  wire _5452 = uncoded_block[103] ^ uncoded_block[108];
  wire _5453 = uncoded_block[110] ^ uncoded_block[111];
  wire _5454 = _5452 ^ _5453;
  wire _5455 = uncoded_block[114] ^ uncoded_block[119];
  wire _5456 = _5455 ^ _2502;
  wire _5457 = _5454 ^ _5456;
  wire _5458 = _5451 ^ _5457;
  wire _5459 = _924 ^ _3263;
  wire _5460 = _4755 ^ _5459;
  wire _5461 = uncoded_block[141] ^ uncoded_block[142];
  wire _5462 = _3265 ^ _5461;
  wire _5463 = uncoded_block[144] ^ uncoded_block[147];
  wire _5464 = _5463 ^ _70;
  wire _5465 = _5462 ^ _5464;
  wire _5466 = _5460 ^ _5465;
  wire _5467 = _5458 ^ _5466;
  wire _5468 = _5447 ^ _5467;
  wire _5469 = uncoded_block[153] ^ uncoded_block[154];
  wire _5470 = uncoded_block[156] ^ uncoded_block[158];
  wire _5471 = _5469 ^ _5470;
  wire _5472 = uncoded_block[162] ^ uncoded_block[165];
  wire _5473 = uncoded_block[169] ^ uncoded_block[170];
  wire _5474 = _5472 ^ _5473;
  wire _5475 = _5471 ^ _5474;
  wire _5476 = uncoded_block[174] ^ uncoded_block[178];
  wire _5477 = uncoded_block[179] ^ uncoded_block[180];
  wire _5478 = _5476 ^ _5477;
  wire _5479 = uncoded_block[181] ^ uncoded_block[182];
  wire _5480 = _5479 ^ _86;
  wire _5481 = _5478 ^ _5480;
  wire _5482 = _5475 ^ _5481;
  wire _5483 = uncoded_block[190] ^ uncoded_block[191];
  wire _5484 = _4772 ^ _5483;
  wire _5485 = uncoded_block[196] ^ uncoded_block[199];
  wire _5486 = uncoded_block[202] ^ uncoded_block[207];
  wire _5487 = _5485 ^ _5486;
  wire _5488 = _5484 ^ _5487;
  wire _5489 = uncoded_block[208] ^ uncoded_block[210];
  wire _5490 = _5489 ^ _956;
  wire _5491 = uncoded_block[214] ^ uncoded_block[217];
  wire _5492 = uncoded_block[220] ^ uncoded_block[221];
  wire _5493 = _5491 ^ _5492;
  wire _5494 = _5490 ^ _5493;
  wire _5495 = _5488 ^ _5494;
  wire _5496 = _5482 ^ _5495;
  wire _5497 = uncoded_block[222] ^ uncoded_block[223];
  wire _5498 = uncoded_block[224] ^ uncoded_block[228];
  wire _5499 = _5497 ^ _5498;
  wire _5500 = uncoded_block[238] ^ uncoded_block[240];
  wire _5501 = _2550 ^ _5500;
  wire _5502 = _5499 ^ _5501;
  wire _5503 = uncoded_block[241] ^ uncoded_block[242];
  wire _5504 = _5503 ^ _4797;
  wire _5505 = uncoded_block[245] ^ uncoded_block[248];
  wire _5506 = _5505 ^ _2559;
  wire _5507 = _5504 ^ _5506;
  wire _5508 = _5502 ^ _5507;
  wire _5509 = _4096 ^ _4098;
  wire _5510 = _4099 ^ _4102;
  wire _5511 = _5509 ^ _5510;
  wire _5512 = uncoded_block[274] ^ uncoded_block[275];
  wire _5513 = uncoded_block[276] ^ uncoded_block[278];
  wire _5514 = _5512 ^ _5513;
  wire _5515 = uncoded_block[280] ^ uncoded_block[281];
  wire _5516 = _5515 ^ _4105;
  wire _5517 = _5514 ^ _5516;
  wire _5518 = _5511 ^ _5517;
  wire _5519 = _5508 ^ _5518;
  wire _5520 = _5496 ^ _5519;
  wire _5521 = _5468 ^ _5520;
  wire _5522 = uncoded_block[287] ^ uncoded_block[288];
  wire _5523 = _5522 ^ _994;
  wire _5524 = uncoded_block[293] ^ uncoded_block[296];
  wire _5525 = uncoded_block[297] ^ uncoded_block[303];
  wire _5526 = _5524 ^ _5525;
  wire _5527 = _5523 ^ _5526;
  wire _5528 = uncoded_block[308] ^ uncoded_block[311];
  wire _5529 = _4114 ^ _5528;
  wire _5530 = uncoded_block[319] ^ uncoded_block[323];
  wire _5531 = _4117 ^ _5530;
  wire _5532 = _5529 ^ _5531;
  wire _5533 = _5527 ^ _5532;
  wire _5534 = uncoded_block[328] ^ uncoded_block[330];
  wire _5535 = _5534 ^ _1821;
  wire _5536 = uncoded_block[334] ^ uncoded_block[335];
  wire _5537 = _5536 ^ _2592;
  wire _5538 = _5535 ^ _5537;
  wire _5539 = uncoded_block[344] ^ uncoded_block[347];
  wire _5540 = _4840 ^ _5539;
  wire _5541 = uncoded_block[349] ^ uncoded_block[350];
  wire _5542 = _5541 ^ _1024;
  wire _5543 = _5540 ^ _5542;
  wire _5544 = _5538 ^ _5543;
  wire _5545 = _5533 ^ _5544;
  wire _5546 = uncoded_block[356] ^ uncoded_block[361];
  wire _5547 = _1028 ^ _5546;
  wire _5548 = uncoded_block[363] ^ uncoded_block[364];
  wire _5549 = uncoded_block[365] ^ uncoded_block[379];
  wire _5550 = _5548 ^ _5549;
  wire _5551 = _5547 ^ _5550;
  wire _5552 = uncoded_block[384] ^ uncoded_block[387];
  wire _5553 = _4857 ^ _5552;
  wire _5554 = uncoded_block[391] ^ uncoded_block[392];
  wire _5555 = _3381 ^ _5554;
  wire _5556 = _5553 ^ _5555;
  wire _5557 = _5551 ^ _5556;
  wire _5558 = uncoded_block[395] ^ uncoded_block[400];
  wire _5559 = uncoded_block[401] ^ uncoded_block[402];
  wire _5560 = _5558 ^ _5559;
  wire _5561 = uncoded_block[404] ^ uncoded_block[406];
  wire _5562 = _5561 ^ _190;
  wire _5563 = _5560 ^ _5562;
  wire _5564 = uncoded_block[411] ^ uncoded_block[414];
  wire _5565 = uncoded_block[415] ^ uncoded_block[416];
  wire _5566 = _5564 ^ _5565;
  wire _5567 = uncoded_block[424] ^ uncoded_block[428];
  wire _5568 = _1854 ^ _5567;
  wire _5569 = _5566 ^ _5568;
  wire _5570 = _5563 ^ _5569;
  wire _5571 = _5557 ^ _5570;
  wire _5572 = _5545 ^ _5571;
  wire _5573 = _4167 ^ _2638;
  wire _5574 = uncoded_block[438] ^ uncoded_block[439];
  wire _5575 = _2640 ^ _5574;
  wire _5576 = _5573 ^ _5575;
  wire _5577 = uncoded_block[440] ^ uncoded_block[441];
  wire _5578 = uncoded_block[442] ^ uncoded_block[443];
  wire _5579 = _5577 ^ _5578;
  wire _5580 = uncoded_block[444] ^ uncoded_block[447];
  wire _5581 = _5580 ^ _2645;
  wire _5582 = _5579 ^ _5581;
  wire _5583 = _5576 ^ _5582;
  wire _5584 = uncoded_block[455] ^ uncoded_block[457];
  wire _5585 = _5584 ^ _3415;
  wire _5586 = uncoded_block[460] ^ uncoded_block[462];
  wire _5587 = uncoded_block[463] ^ uncoded_block[470];
  wire _5588 = _5586 ^ _5587;
  wire _5589 = _5585 ^ _5588;
  wire _5590 = uncoded_block[476] ^ uncoded_block[477];
  wire _5591 = _1083 ^ _5590;
  wire _5592 = uncoded_block[478] ^ uncoded_block[479];
  wire _5593 = uncoded_block[480] ^ uncoded_block[481];
  wire _5594 = _5592 ^ _5593;
  wire _5595 = _5591 ^ _5594;
  wire _5596 = _5589 ^ _5595;
  wire _5597 = _5583 ^ _5596;
  wire _5598 = uncoded_block[482] ^ uncoded_block[484];
  wire _5599 = _5598 ^ _2660;
  wire _5600 = uncoded_block[488] ^ uncoded_block[490];
  wire _5601 = _5600 ^ _4902;
  wire _5602 = _5599 ^ _5601;
  wire _5603 = uncoded_block[495] ^ uncoded_block[496];
  wire _5604 = uncoded_block[497] ^ uncoded_block[498];
  wire _5605 = _5603 ^ _5604;
  wire _5606 = uncoded_block[500] ^ uncoded_block[503];
  wire _5607 = uncoded_block[504] ^ uncoded_block[506];
  wire _5608 = _5606 ^ _5607;
  wire _5609 = _5605 ^ _5608;
  wire _5610 = _5602 ^ _5609;
  wire _5611 = uncoded_block[507] ^ uncoded_block[508];
  wire _5612 = _5611 ^ _4908;
  wire _5613 = uncoded_block[512] ^ uncoded_block[516];
  wire _5614 = _5613 ^ _2681;
  wire _5615 = _5612 ^ _5614;
  wire _5616 = uncoded_block[524] ^ uncoded_block[530];
  wire _5617 = uncoded_block[533] ^ uncoded_block[536];
  wire _5618 = _5616 ^ _5617;
  wire _5619 = uncoded_block[537] ^ uncoded_block[538];
  wire _5620 = uncoded_block[539] ^ uncoded_block[543];
  wire _5621 = _5619 ^ _5620;
  wire _5622 = _5618 ^ _5621;
  wire _5623 = _5615 ^ _5622;
  wire _5624 = _5610 ^ _5623;
  wire _5625 = _5597 ^ _5624;
  wire _5626 = _5572 ^ _5625;
  wire _5627 = _5521 ^ _5626;
  wire _5628 = uncoded_block[546] ^ uncoded_block[547];
  wire _5629 = _1117 ^ _5628;
  wire _5630 = uncoded_block[551] ^ uncoded_block[553];
  wire _5631 = _4933 ^ _5630;
  wire _5632 = _5629 ^ _5631;
  wire _5633 = uncoded_block[561] ^ uncoded_block[563];
  wire _5634 = _1122 ^ _5633;
  wire _5635 = uncoded_block[565] ^ uncoded_block[567];
  wire _5636 = _5635 ^ _3468;
  wire _5637 = _5634 ^ _5636;
  wire _5638 = _5632 ^ _5637;
  wire _5639 = uncoded_block[571] ^ uncoded_block[576];
  wire _5640 = _5639 ^ _1133;
  wire _5641 = uncoded_block[581] ^ uncoded_block[584];
  wire _5642 = _5641 ^ _4947;
  wire _5643 = _5640 ^ _5642;
  wire _5644 = uncoded_block[588] ^ uncoded_block[596];
  wire _5645 = _5644 ^ _4953;
  wire _5646 = uncoded_block[601] ^ uncoded_block[603];
  wire _5647 = uncoded_block[604] ^ uncoded_block[609];
  wire _5648 = _5646 ^ _5647;
  wire _5649 = _5645 ^ _5648;
  wire _5650 = _5643 ^ _5649;
  wire _5651 = _5638 ^ _5650;
  wire _5652 = uncoded_block[613] ^ uncoded_block[614];
  wire _5653 = uncoded_block[615] ^ uncoded_block[617];
  wire _5654 = _5652 ^ _5653;
  wire _5655 = uncoded_block[622] ^ uncoded_block[625];
  wire _5656 = _4243 ^ _5655;
  wire _5657 = _5654 ^ _5656;
  wire _5658 = uncoded_block[628] ^ uncoded_block[629];
  wire _5659 = _1154 ^ _5658;
  wire _5660 = uncoded_block[630] ^ uncoded_block[634];
  wire _5661 = uncoded_block[635] ^ uncoded_block[636];
  wire _5662 = _5660 ^ _5661;
  wire _5663 = _5659 ^ _5662;
  wire _5664 = _5657 ^ _5663;
  wire _5665 = uncoded_block[638] ^ uncoded_block[640];
  wire _5666 = _5665 ^ _294;
  wire _5667 = _1164 ^ _297;
  wire _5668 = _5666 ^ _5667;
  wire _5669 = _1170 ^ _3513;
  wire _5670 = uncoded_block[660] ^ uncoded_block[663];
  wire _5671 = uncoded_block[664] ^ uncoded_block[668];
  wire _5672 = _5670 ^ _5671;
  wire _5673 = _5669 ^ _5672;
  wire _5674 = _5668 ^ _5673;
  wire _5675 = _5664 ^ _5674;
  wire _5676 = _5651 ^ _5675;
  wire _5677 = _2744 ^ _3522;
  wire _5678 = uncoded_block[683] ^ uncoded_block[685];
  wire _5679 = _5678 ^ _322;
  wire _5680 = _5677 ^ _5679;
  wire _5681 = _325 ^ _4272;
  wire _5682 = _328 ^ _3529;
  wire _5683 = _5681 ^ _5682;
  wire _5684 = _5680 ^ _5683;
  wire _5685 = uncoded_block[703] ^ uncoded_block[705];
  wire _5686 = _333 ^ _5685;
  wire _5687 = uncoded_block[711] ^ uncoded_block[718];
  wire _5688 = _4996 ^ _5687;
  wire _5689 = _5686 ^ _5688;
  wire _5690 = uncoded_block[719] ^ uncoded_block[721];
  wire _5691 = uncoded_block[722] ^ uncoded_block[725];
  wire _5692 = _5690 ^ _5691;
  wire _5693 = uncoded_block[726] ^ uncoded_block[728];
  wire _5694 = _5693 ^ _1991;
  wire _5695 = _5692 ^ _5694;
  wire _5696 = _5689 ^ _5695;
  wire _5697 = _5684 ^ _5696;
  wire _5698 = _3547 ^ _1995;
  wire _5699 = uncoded_block[742] ^ uncoded_block[743];
  wire _5700 = _1996 ^ _5699;
  wire _5701 = _5698 ^ _5700;
  wire _5702 = uncoded_block[744] ^ uncoded_block[745];
  wire _5703 = _5702 ^ _1999;
  wire _5704 = uncoded_block[748] ^ uncoded_block[749];
  wire _5705 = _5704 ^ _2778;
  wire _5706 = _5703 ^ _5705;
  wire _5707 = _5701 ^ _5706;
  wire _5708 = uncoded_block[757] ^ uncoded_block[763];
  wire _5709 = uncoded_block[766] ^ uncoded_block[768];
  wire _5710 = _5708 ^ _5709;
  wire _5711 = uncoded_block[774] ^ uncoded_block[775];
  wire _5712 = _1218 ^ _5711;
  wire _5713 = _5710 ^ _5712;
  wire _5714 = _2014 ^ _368;
  wire _5715 = uncoded_block[781] ^ uncoded_block[784];
  wire _5716 = _5715 ^ _2018;
  wire _5717 = _5714 ^ _5716;
  wire _5718 = _5713 ^ _5717;
  wire _5719 = _5707 ^ _5718;
  wire _5720 = _5697 ^ _5719;
  wire _5721 = _5676 ^ _5720;
  wire _5722 = _5033 ^ _374;
  wire _5723 = uncoded_block[793] ^ uncoded_block[796];
  wire _5724 = _5723 ^ _385;
  wire _5725 = _5722 ^ _5724;
  wire _5726 = uncoded_block[802] ^ uncoded_block[804];
  wire _5727 = uncoded_block[805] ^ uncoded_block[808];
  wire _5728 = _5726 ^ _5727;
  wire _5729 = uncoded_block[811] ^ uncoded_block[814];
  wire _5730 = _392 ^ _5729;
  wire _5731 = _5728 ^ _5730;
  wire _5732 = _5725 ^ _5731;
  wire _5733 = uncoded_block[818] ^ uncoded_block[826];
  wire _5734 = uncoded_block[828] ^ uncoded_block[830];
  wire _5735 = _5733 ^ _5734;
  wire _5736 = uncoded_block[833] ^ uncoded_block[838];
  wire _5737 = uncoded_block[840] ^ uncoded_block[842];
  wire _5738 = _5736 ^ _5737;
  wire _5739 = _5735 ^ _5738;
  wire _5740 = _3597 ^ _1257;
  wire _5741 = uncoded_block[848] ^ uncoded_block[851];
  wire _5742 = uncoded_block[856] ^ uncoded_block[858];
  wire _5743 = _5741 ^ _5742;
  wire _5744 = _5740 ^ _5743;
  wire _5745 = _5739 ^ _5744;
  wire _5746 = _5732 ^ _5745;
  wire _5747 = uncoded_block[859] ^ uncoded_block[860];
  wire _5748 = _5747 ^ _2824;
  wire _5749 = uncoded_block[868] ^ uncoded_block[870];
  wire _5750 = _2827 ^ _5749;
  wire _5751 = _5748 ^ _5750;
  wire _5752 = uncoded_block[871] ^ uncoded_block[876];
  wire _5753 = uncoded_block[877] ^ uncoded_block[881];
  wire _5754 = _5752 ^ _5753;
  wire _5755 = _4352 ^ _2061;
  wire _5756 = _5754 ^ _5755;
  wire _5757 = _5751 ^ _5756;
  wire _5758 = uncoded_block[896] ^ uncoded_block[897];
  wire _5759 = uncoded_block[898] ^ uncoded_block[901];
  wire _5760 = _5758 ^ _5759;
  wire _5761 = uncoded_block[905] ^ uncoded_block[909];
  wire _5762 = uncoded_block[912] ^ uncoded_block[914];
  wire _5763 = _5761 ^ _5762;
  wire _5764 = _5760 ^ _5763;
  wire _5765 = _3629 ^ _3631;
  wire _5766 = uncoded_block[923] ^ uncoded_block[924];
  wire _5767 = _3632 ^ _5766;
  wire _5768 = _5765 ^ _5767;
  wire _5769 = _5764 ^ _5768;
  wire _5770 = _5757 ^ _5769;
  wire _5771 = _5746 ^ _5770;
  wire _5772 = uncoded_block[925] ^ uncoded_block[929];
  wire _5773 = uncoded_block[930] ^ uncoded_block[933];
  wire _5774 = _5772 ^ _5773;
  wire _5775 = _5774 ^ _5102;
  wire _5776 = uncoded_block[942] ^ uncoded_block[947];
  wire _5777 = uncoded_block[948] ^ uncoded_block[949];
  wire _5778 = _5776 ^ _5777;
  wire _5779 = uncoded_block[952] ^ uncoded_block[953];
  wire _5780 = _5779 ^ _4384;
  wire _5781 = _5778 ^ _5780;
  wire _5782 = _5775 ^ _5781;
  wire _5783 = uncoded_block[961] ^ uncoded_block[963];
  wire _5784 = _5783 ^ _2092;
  wire _5785 = uncoded_block[967] ^ uncoded_block[969];
  wire _5786 = uncoded_block[970] ^ uncoded_block[975];
  wire _5787 = _5785 ^ _5786;
  wire _5788 = _5784 ^ _5787;
  wire _5789 = uncoded_block[977] ^ uncoded_block[978];
  wire _5790 = uncoded_block[980] ^ uncoded_block[981];
  wire _5791 = _5789 ^ _5790;
  wire _5792 = uncoded_block[982] ^ uncoded_block[983];
  wire _5793 = _5792 ^ _2882;
  wire _5794 = _5791 ^ _5793;
  wire _5795 = _5788 ^ _5794;
  wire _5796 = _5782 ^ _5795;
  wire _5797 = uncoded_block[992] ^ uncoded_block[997];
  wire _5798 = uncoded_block[998] ^ uncoded_block[999];
  wire _5799 = _5797 ^ _5798;
  wire _5800 = uncoded_block[1001] ^ uncoded_block[1007];
  wire _5801 = uncoded_block[1008] ^ uncoded_block[1015];
  wire _5802 = _5800 ^ _5801;
  wire _5803 = _5799 ^ _5802;
  wire _5804 = uncoded_block[1016] ^ uncoded_block[1019];
  wire _5805 = _5804 ^ _2120;
  wire _5806 = uncoded_block[1030] ^ uncoded_block[1032];
  wire _5807 = _2121 ^ _5806;
  wire _5808 = _5805 ^ _5807;
  wire _5809 = _5803 ^ _5808;
  wire _5810 = uncoded_block[1037] ^ uncoded_block[1039];
  wire _5811 = _1342 ^ _5810;
  wire _5812 = uncoded_block[1040] ^ uncoded_block[1044];
  wire _5813 = _5812 ^ _2133;
  wire _5814 = _5811 ^ _5813;
  wire _5815 = _515 ^ _1357;
  wire _5816 = uncoded_block[1056] ^ uncoded_block[1060];
  wire _5817 = _2136 ^ _5816;
  wire _5818 = _5815 ^ _5817;
  wire _5819 = _5814 ^ _5818;
  wire _5820 = _5809 ^ _5819;
  wire _5821 = _5796 ^ _5820;
  wire _5822 = _5771 ^ _5821;
  wire _5823 = _5721 ^ _5822;
  wire _5824 = _5627 ^ _5823;
  wire _5825 = uncoded_block[1061] ^ uncoded_block[1062];
  wire _5826 = uncoded_block[1063] ^ uncoded_block[1066];
  wire _5827 = _5825 ^ _5826;
  wire _5828 = uncoded_block[1067] ^ uncoded_block[1070];
  wire _5829 = _5828 ^ _527;
  wire _5830 = _5827 ^ _5829;
  wire _5831 = uncoded_block[1073] ^ uncoded_block[1074];
  wire _5832 = uncoded_block[1075] ^ uncoded_block[1078];
  wire _5833 = _5831 ^ _5832;
  wire _5834 = uncoded_block[1079] ^ uncoded_block[1080];
  wire _5835 = uncoded_block[1081] ^ uncoded_block[1084];
  wire _5836 = _5834 ^ _5835;
  wire _5837 = _5833 ^ _5836;
  wire _5838 = _5830 ^ _5837;
  wire _5839 = uncoded_block[1086] ^ uncoded_block[1089];
  wire _5840 = uncoded_block[1091] ^ uncoded_block[1092];
  wire _5841 = _5839 ^ _5840;
  wire _5842 = uncoded_block[1093] ^ uncoded_block[1095];
  wire _5843 = uncoded_block[1096] ^ uncoded_block[1097];
  wire _5844 = _5842 ^ _5843;
  wire _5845 = _5841 ^ _5844;
  wire _5846 = uncoded_block[1098] ^ uncoded_block[1100];
  wire _5847 = _5846 ^ _2160;
  wire _5848 = uncoded_block[1115] ^ uncoded_block[1118];
  wire _5849 = _1386 ^ _5848;
  wire _5850 = _5847 ^ _5849;
  wire _5851 = _5845 ^ _5850;
  wire _5852 = _5838 ^ _5851;
  wire _5853 = uncoded_block[1119] ^ uncoded_block[1122];
  wire _5854 = uncoded_block[1125] ^ uncoded_block[1126];
  wire _5855 = _5853 ^ _5854;
  wire _5856 = uncoded_block[1134] ^ uncoded_block[1135];
  wire _5857 = _560 ^ _5856;
  wire _5858 = _5855 ^ _5857;
  wire _5859 = uncoded_block[1141] ^ uncoded_block[1142];
  wire _5860 = _565 ^ _5859;
  wire _5861 = uncoded_block[1143] ^ uncoded_block[1145];
  wire _5862 = uncoded_block[1146] ^ uncoded_block[1148];
  wire _5863 = _5861 ^ _5862;
  wire _5864 = _5860 ^ _5863;
  wire _5865 = _5858 ^ _5864;
  wire _5866 = uncoded_block[1149] ^ uncoded_block[1154];
  wire _5867 = _5866 ^ _5190;
  wire _5868 = _5867 ^ _2959;
  wire _5869 = uncoded_block[1163] ^ uncoded_block[1168];
  wire _5870 = uncoded_block[1169] ^ uncoded_block[1171];
  wire _5871 = _5869 ^ _5870;
  wire _5872 = uncoded_block[1176] ^ uncoded_block[1177];
  wire _5873 = uncoded_block[1178] ^ uncoded_block[1181];
  wire _5874 = _5872 ^ _5873;
  wire _5875 = _5871 ^ _5874;
  wire _5876 = _5868 ^ _5875;
  wire _5877 = _5865 ^ _5876;
  wire _5878 = _5852 ^ _5877;
  wire _5879 = _592 ^ _4486;
  wire _5880 = _2200 ^ _596;
  wire _5881 = _5879 ^ _5880;
  wire _5882 = uncoded_block[1196] ^ uncoded_block[1199];
  wire _5883 = uncoded_block[1200] ^ uncoded_block[1204];
  wire _5884 = _5882 ^ _5883;
  wire _5885 = uncoded_block[1205] ^ uncoded_block[1207];
  wire _5886 = _5885 ^ _1428;
  wire _5887 = _5884 ^ _5886;
  wire _5888 = _5881 ^ _5887;
  wire _5889 = uncoded_block[1214] ^ uncoded_block[1216];
  wire _5890 = _5889 ^ _4499;
  wire _5891 = uncoded_block[1224] ^ uncoded_block[1226];
  wire _5892 = _4502 ^ _5891;
  wire _5893 = _5890 ^ _5892;
  wire _5894 = uncoded_block[1228] ^ uncoded_block[1230];
  wire _5895 = _5894 ^ _1442;
  wire _5896 = _1443 ^ _1448;
  wire _5897 = _5895 ^ _5896;
  wire _5898 = _5893 ^ _5897;
  wire _5899 = _5888 ^ _5898;
  wire _5900 = _3777 ^ _1451;
  wire _5901 = uncoded_block[1250] ^ uncoded_block[1252];
  wire _5902 = uncoded_block[1254] ^ uncoded_block[1258];
  wire _5903 = _5901 ^ _5902;
  wire _5904 = _5900 ^ _5903;
  wire _5905 = uncoded_block[1271] ^ uncoded_block[1273];
  wire _5906 = _2238 ^ _5905;
  wire _5907 = uncoded_block[1274] ^ uncoded_block[1276];
  wire _5908 = uncoded_block[1277] ^ uncoded_block[1278];
  wire _5909 = _5907 ^ _5908;
  wire _5910 = _5906 ^ _5909;
  wire _5911 = _5904 ^ _5910;
  wire _5912 = _631 ^ _3797;
  wire _5913 = uncoded_block[1286] ^ uncoded_block[1288];
  wire _5914 = _5913 ^ _641;
  wire _5915 = _5912 ^ _5914;
  wire _5916 = uncoded_block[1292] ^ uncoded_block[1298];
  wire _5917 = uncoded_block[1300] ^ uncoded_block[1306];
  wire _5918 = _5916 ^ _5917;
  wire _5919 = uncoded_block[1312] ^ uncoded_block[1314];
  wire _5920 = _3807 ^ _5919;
  wire _5921 = _5918 ^ _5920;
  wire _5922 = _5915 ^ _5921;
  wire _5923 = _5911 ^ _5922;
  wire _5924 = _5899 ^ _5923;
  wire _5925 = _5878 ^ _5924;
  wire _5926 = uncoded_block[1316] ^ uncoded_block[1318];
  wire _5927 = uncoded_block[1320] ^ uncoded_block[1323];
  wire _5928 = _5926 ^ _5927;
  wire _5929 = _656 ^ _4545;
  wire _5930 = _5928 ^ _5929;
  wire _5931 = uncoded_block[1331] ^ uncoded_block[1333];
  wire _5932 = uncoded_block[1334] ^ uncoded_block[1336];
  wire _5933 = _5931 ^ _5932;
  wire _5934 = _2277 ^ _5266;
  wire _5935 = _5933 ^ _5934;
  wire _5936 = _5930 ^ _5935;
  wire _5937 = uncoded_block[1345] ^ uncoded_block[1350];
  wire _5938 = uncoded_block[1351] ^ uncoded_block[1353];
  wire _5939 = _5937 ^ _5938;
  wire _5940 = uncoded_block[1357] ^ uncoded_block[1358];
  wire _5941 = _5272 ^ _5940;
  wire _5942 = _5939 ^ _5941;
  wire _5943 = uncoded_block[1360] ^ uncoded_block[1364];
  wire _5944 = uncoded_block[1365] ^ uncoded_block[1373];
  wire _5945 = _5943 ^ _5944;
  wire _5946 = _2289 ^ _3055;
  wire _5947 = _5945 ^ _5946;
  wire _5948 = _5942 ^ _5947;
  wire _5949 = _5936 ^ _5948;
  wire _5950 = uncoded_block[1387] ^ uncoded_block[1388];
  wire _5951 = _3061 ^ _5950;
  wire _5952 = uncoded_block[1392] ^ uncoded_block[1393];
  wire _5953 = _5952 ^ _694;
  wire _5954 = _5951 ^ _5953;
  wire _5955 = uncoded_block[1397] ^ uncoded_block[1398];
  wire _5956 = _5955 ^ _1519;
  wire _5957 = uncoded_block[1408] ^ uncoded_block[1409];
  wire _5958 = _2300 ^ _5957;
  wire _5959 = _5956 ^ _5958;
  wire _5960 = _5954 ^ _5959;
  wire _5961 = uncoded_block[1410] ^ uncoded_block[1411];
  wire _5962 = uncoded_block[1412] ^ uncoded_block[1414];
  wire _5963 = _5961 ^ _5962;
  wire _5964 = uncoded_block[1418] ^ uncoded_block[1421];
  wire _5965 = _2306 ^ _5964;
  wire _5966 = _5963 ^ _5965;
  wire _5967 = uncoded_block[1424] ^ uncoded_block[1427];
  wire _5968 = uncoded_block[1429] ^ uncoded_block[1430];
  wire _5969 = _5967 ^ _5968;
  wire _5970 = uncoded_block[1442] ^ uncoded_block[1445];
  wire _5971 = _1540 ^ _5970;
  wire _5972 = _5969 ^ _5971;
  wire _5973 = _5966 ^ _5972;
  wire _5974 = _5960 ^ _5973;
  wire _5975 = _5949 ^ _5974;
  wire _5976 = uncoded_block[1449] ^ uncoded_block[1452];
  wire _5977 = _2322 ^ _5976;
  wire _5978 = uncoded_block[1454] ^ uncoded_block[1458];
  wire _5979 = _5978 ^ _726;
  wire _5980 = _5977 ^ _5979;
  wire _5981 = uncoded_block[1463] ^ uncoded_block[1466];
  wire _5982 = _5981 ^ _1550;
  wire _5983 = uncoded_block[1470] ^ uncoded_block[1471];
  wire _5984 = uncoded_block[1473] ^ uncoded_block[1481];
  wire _5985 = _5983 ^ _5984;
  wire _5986 = _5982 ^ _5985;
  wire _5987 = _5980 ^ _5986;
  wire _5988 = uncoded_block[1484] ^ uncoded_block[1485];
  wire _5989 = _1559 ^ _5988;
  wire _5990 = uncoded_block[1488] ^ uncoded_block[1492];
  wire _5991 = _739 ^ _5990;
  wire _5992 = _5989 ^ _5991;
  wire _5993 = uncoded_block[1499] ^ uncoded_block[1502];
  wire _5994 = _1566 ^ _5993;
  wire _5995 = _1572 ^ _5334;
  wire _5996 = _5994 ^ _5995;
  wire _5997 = _5992 ^ _5996;
  wire _5998 = _5987 ^ _5997;
  wire _5999 = uncoded_block[1519] ^ uncoded_block[1524];
  wire _6000 = _751 ^ _5999;
  wire _6001 = uncoded_block[1526] ^ uncoded_block[1529];
  wire _6002 = uncoded_block[1530] ^ uncoded_block[1531];
  wire _6003 = _6001 ^ _6002;
  wire _6004 = _6000 ^ _6003;
  wire _6005 = uncoded_block[1532] ^ uncoded_block[1533];
  wire _6006 = uncoded_block[1535] ^ uncoded_block[1538];
  wire _6007 = _6005 ^ _6006;
  wire _6008 = uncoded_block[1542] ^ uncoded_block[1543];
  wire _6009 = _5350 ^ _6008;
  wire _6010 = _6007 ^ _6009;
  wire _6011 = _6004 ^ _6010;
  wire _6012 = uncoded_block[1544] ^ uncoded_block[1547];
  wire _6013 = uncoded_block[1548] ^ uncoded_block[1550];
  wire _6014 = _6012 ^ _6013;
  wire _6015 = uncoded_block[1551] ^ uncoded_block[1556];
  wire _6016 = uncoded_block[1557] ^ uncoded_block[1559];
  wire _6017 = _6015 ^ _6016;
  wire _6018 = _6014 ^ _6017;
  wire _6019 = uncoded_block[1564] ^ uncoded_block[1566];
  wire _6020 = _4640 ^ _6019;
  wire _6021 = _1606 ^ _4645;
  wire _6022 = _6020 ^ _6021;
  wire _6023 = _6018 ^ _6022;
  wire _6024 = _6011 ^ _6023;
  wire _6025 = _5998 ^ _6024;
  wire _6026 = _5975 ^ _6025;
  wire _6027 = _5925 ^ _6026;
  wire _6028 = uncoded_block[1573] ^ uncoded_block[1576];
  wire _6029 = uncoded_block[1577] ^ uncoded_block[1580];
  wire _6030 = _6028 ^ _6029;
  wire _6031 = uncoded_block[1581] ^ uncoded_block[1582];
  wire _6032 = _6031 ^ _785;
  wire _6033 = _6030 ^ _6032;
  wire _6034 = uncoded_block[1585] ^ uncoded_block[1589];
  wire _6035 = _6034 ^ _3146;
  wire _6036 = _4654 ^ _5373;
  wire _6037 = _6035 ^ _6036;
  wire _6038 = _6033 ^ _6037;
  wire _6039 = uncoded_block[1602] ^ uncoded_block[1603];
  wire _6040 = uncoded_block[1608] ^ uncoded_block[1609];
  wire _6041 = _6039 ^ _6040;
  wire _6042 = uncoded_block[1613] ^ uncoded_block[1614];
  wire _6043 = uncoded_block[1615] ^ uncoded_block[1619];
  wire _6044 = _6042 ^ _6043;
  wire _6045 = _6041 ^ _6044;
  wire _6046 = uncoded_block[1624] ^ uncoded_block[1625];
  wire _6047 = _6046 ^ _3161;
  wire _6048 = uncoded_block[1630] ^ uncoded_block[1633];
  wire _6049 = uncoded_block[1634] ^ uncoded_block[1638];
  wire _6050 = _6048 ^ _6049;
  wire _6051 = _6047 ^ _6050;
  wire _6052 = _6045 ^ _6051;
  wire _6053 = _6038 ^ _6052;
  wire _6054 = _4674 ^ _4677;
  wire _6055 = uncoded_block[1660] ^ uncoded_block[1661];
  wire _6056 = _3174 ^ _6055;
  wire _6057 = _6054 ^ _6056;
  wire _6058 = uncoded_block[1667] ^ uncoded_block[1670];
  wire _6059 = uncoded_block[1671] ^ uncoded_block[1674];
  wire _6060 = _6058 ^ _6059;
  wire _6061 = uncoded_block[1682] ^ uncoded_block[1684];
  wire _6062 = _5406 ^ _6061;
  wire _6063 = _6060 ^ _6062;
  wire _6064 = _6057 ^ _6063;
  wire _6065 = uncoded_block[1686] ^ uncoded_block[1691];
  wire _6066 = uncoded_block[1693] ^ uncoded_block[1694];
  wire _6067 = _6065 ^ _6066;
  wire _6068 = uncoded_block[1700] ^ uncoded_block[1701];
  wire _6069 = _844 ^ _6068;
  wire _6070 = _6067 ^ _6069;
  wire _6071 = uncoded_block[1706] ^ uncoded_block[1711];
  wire _6072 = uncoded_block[1714] ^ uncoded_block[1717];
  wire _6073 = _6071 ^ _6072;
  wire _6074 = _6073 ^ _5416;
  wire _6075 = _6070 ^ _6074;
  wire _6076 = _6064 ^ _6075;
  wire _6077 = _6053 ^ _6076;
  wire _6078 = _6027 ^ _6077;
  wire _6079 = _5824 ^ _6078;
  wire _6080 = uncoded_block[4] ^ uncoded_block[5];
  wire _6081 = _3210 ^ _6080;
  wire _6082 = uncoded_block[6] ^ uncoded_block[8];
  wire _6083 = uncoded_block[10] ^ uncoded_block[11];
  wire _6084 = _6082 ^ _6083;
  wire _6085 = _6081 ^ _6084;
  wire _6086 = uncoded_block[13] ^ uncoded_block[15];
  wire _6087 = uncoded_block[17] ^ uncoded_block[18];
  wire _6088 = _6086 ^ _6087;
  wire _6089 = uncoded_block[23] ^ uncoded_block[26];
  wire _6090 = _3217 ^ _6089;
  wire _6091 = _6088 ^ _6090;
  wire _6092 = _6085 ^ _6091;
  wire _6093 = uncoded_block[27] ^ uncoded_block[29];
  wire _6094 = _6093 ^ _875;
  wire _6095 = uncoded_block[33] ^ uncoded_block[34];
  wire _6096 = uncoded_block[39] ^ uncoded_block[42];
  wire _6097 = _6095 ^ _6096;
  wire _6098 = _6094 ^ _6097;
  wire _6099 = uncoded_block[47] ^ uncoded_block[48];
  wire _6100 = _4009 ^ _6099;
  wire _6101 = uncoded_block[49] ^ uncoded_block[51];
  wire _6102 = _6101 ^ _25;
  wire _6103 = _6100 ^ _6102;
  wire _6104 = _6098 ^ _6103;
  wire _6105 = _6092 ^ _6104;
  wire _6106 = uncoded_block[57] ^ uncoded_block[62];
  wire _6107 = uncoded_block[65] ^ uncoded_block[70];
  wire _6108 = _6106 ^ _6107;
  wire _6109 = uncoded_block[75] ^ uncoded_block[79];
  wire _6110 = _5442 ^ _6109;
  wire _6111 = _6108 ^ _6110;
  wire _6112 = uncoded_block[80] ^ uncoded_block[86];
  wire _6113 = uncoded_block[87] ^ uncoded_block[90];
  wire _6114 = _6112 ^ _6113;
  wire _6115 = uncoded_block[93] ^ uncoded_block[94];
  wire _6116 = uncoded_block[97] ^ uncoded_block[100];
  wire _6117 = _6115 ^ _6116;
  wire _6118 = _6114 ^ _6117;
  wire _6119 = _6111 ^ _6118;
  wire _6120 = uncoded_block[104] ^ uncoded_block[105];
  wire _6121 = _4028 ^ _6120;
  wire _6122 = uncoded_block[106] ^ uncoded_block[107];
  wire _6123 = uncoded_block[109] ^ uncoded_block[110];
  wire _6124 = _6122 ^ _6123;
  wire _6125 = _6121 ^ _6124;
  wire _6126 = uncoded_block[111] ^ uncoded_block[113];
  wire _6127 = _6126 ^ _2495;
  wire _6128 = uncoded_block[117] ^ uncoded_block[119];
  wire _6129 = _6128 ^ _1730;
  wire _6130 = _6127 ^ _6129;
  wire _6131 = _6125 ^ _6130;
  wire _6132 = _6119 ^ _6131;
  wire _6133 = _6105 ^ _6132;
  wire _6134 = _3262 ^ _4754;
  wire _6135 = _6134 ^ _5459;
  wire _6136 = uncoded_block[138] ^ uncoded_block[140];
  wire _6137 = _6136 ^ _5461;
  wire _6138 = uncoded_block[143] ^ uncoded_block[144];
  wire _6139 = uncoded_block[145] ^ uncoded_block[151];
  wire _6140 = _6138 ^ _6139;
  wire _6141 = _6137 ^ _6140;
  wire _6142 = _6135 ^ _6141;
  wire _6143 = _5469 ^ _1748;
  wire _6144 = uncoded_block[160] ^ uncoded_block[162];
  wire _6145 = _6144 ^ _1749;
  wire _6146 = _6143 ^ _6145;
  wire _6147 = uncoded_block[170] ^ uncoded_block[174];
  wire _6148 = _4056 ^ _6147;
  wire _6149 = uncoded_block[175] ^ uncoded_block[176];
  wire _6150 = _6149 ^ _4060;
  wire _6151 = _6148 ^ _6150;
  wire _6152 = _6146 ^ _6151;
  wire _6153 = _6142 ^ _6152;
  wire _6154 = _944 ^ _4772;
  wire _6155 = uncoded_block[191] ^ uncoded_block[195];
  wire _6156 = _4773 ^ _6155;
  wire _6157 = _6154 ^ _6156;
  wire _6158 = uncoded_block[200] ^ uncoded_block[204];
  wire _6159 = _2532 ^ _6158;
  wire _6160 = uncoded_block[205] ^ uncoded_block[210];
  wire _6161 = uncoded_block[212] ^ uncoded_block[215];
  wire _6162 = _6160 ^ _6161;
  wire _6163 = _6159 ^ _6162;
  wire _6164 = _6157 ^ _6163;
  wire _6165 = _4074 ^ _4787;
  wire _6166 = _4788 ^ _4076;
  wire _6167 = _6165 ^ _6166;
  wire _6168 = uncoded_block[226] ^ uncoded_block[227];
  wire _6169 = uncoded_block[228] ^ uncoded_block[230];
  wire _6170 = _6168 ^ _6169;
  wire _6171 = uncoded_block[231] ^ uncoded_block[236];
  wire _6172 = uncoded_block[241] ^ uncoded_block[243];
  wire _6173 = _6171 ^ _6172;
  wire _6174 = _6170 ^ _6173;
  wire _6175 = _6167 ^ _6174;
  wire _6176 = _6164 ^ _6175;
  wire _6177 = _6153 ^ _6176;
  wire _6178 = _6133 ^ _6177;
  wire _6179 = uncoded_block[244] ^ uncoded_block[245];
  wire _6180 = uncoded_block[246] ^ uncoded_block[247];
  wire _6181 = _6179 ^ _6180;
  wire _6182 = uncoded_block[250] ^ uncoded_block[254];
  wire _6183 = _6182 ^ _3311;
  wire _6184 = _6181 ^ _6183;
  wire _6185 = uncoded_block[261] ^ uncoded_block[262];
  wire _6186 = _1788 ^ _6185;
  wire _6187 = uncoded_block[263] ^ uncoded_block[264];
  wire _6188 = uncoded_block[265] ^ uncoded_block[266];
  wire _6189 = _6187 ^ _6188;
  wire _6190 = _6186 ^ _6189;
  wire _6191 = _6184 ^ _6190;
  wire _6192 = uncoded_block[272] ^ uncoded_block[275];
  wire _6193 = _2566 ^ _6192;
  wire _6194 = uncoded_block[279] ^ uncoded_block[280];
  wire _6195 = _1795 ^ _6194;
  wire _6196 = _6193 ^ _6195;
  wire _6197 = uncoded_block[283] ^ uncoded_block[287];
  wire _6198 = _6197 ^ _135;
  wire _6199 = _3328 ^ _137;
  wire _6200 = _6198 ^ _6199;
  wire _6201 = _6196 ^ _6200;
  wire _6202 = _6191 ^ _6201;
  wire _6203 = _1807 ^ _1810;
  wire _6204 = _4826 ^ _3334;
  wire _6205 = _6203 ^ _6204;
  wire _6206 = uncoded_block[309] ^ uncoded_block[314];
  wire _6207 = _6206 ^ _1006;
  wire _6208 = uncoded_block[318] ^ uncoded_block[320];
  wire _6209 = uncoded_block[321] ^ uncoded_block[325];
  wire _6210 = _6208 ^ _6209;
  wire _6211 = _6207 ^ _6210;
  wire _6212 = _6205 ^ _6211;
  wire _6213 = uncoded_block[327] ^ uncoded_block[331];
  wire _6214 = _6213 ^ _5536;
  wire _6215 = _2592 ^ _1825;
  wire _6216 = _6214 ^ _6215;
  wire _6217 = uncoded_block[340] ^ uncoded_block[341];
  wire _6218 = uncoded_block[344] ^ uncoded_block[345];
  wire _6219 = _6217 ^ _6218;
  wire _6220 = uncoded_block[348] ^ uncoded_block[353];
  wire _6221 = uncoded_block[355] ^ uncoded_block[357];
  wire _6222 = _6220 ^ _6221;
  wire _6223 = _6219 ^ _6222;
  wire _6224 = _6216 ^ _6223;
  wire _6225 = _6212 ^ _6224;
  wire _6226 = _6202 ^ _6225;
  wire _6227 = uncoded_block[358] ^ uncoded_block[360];
  wire _6228 = uncoded_block[361] ^ uncoded_block[362];
  wire _6229 = _6227 ^ _6228;
  wire _6230 = _4851 ^ _1835;
  wire _6231 = _6229 ^ _6230;
  wire _6232 = uncoded_block[371] ^ uncoded_block[375];
  wire _6233 = uncoded_block[376] ^ uncoded_block[377];
  wire _6234 = _6232 ^ _6233;
  wire _6235 = uncoded_block[379] ^ uncoded_block[382];
  wire _6236 = _6235 ^ _2613;
  wire _6237 = _6234 ^ _6236;
  wire _6238 = _6231 ^ _6237;
  wire _6239 = uncoded_block[389] ^ uncoded_block[390];
  wire _6240 = _6239 ^ _5554;
  wire _6241 = uncoded_block[396] ^ uncoded_block[403];
  wire _6242 = _1847 ^ _6241;
  wire _6243 = _6240 ^ _6242;
  wire _6244 = uncoded_block[404] ^ uncoded_block[405];
  wire _6245 = _6244 ^ _184;
  wire _6246 = _6245 ^ _2631;
  wire _6247 = _6243 ^ _6246;
  wire _6248 = _6238 ^ _6247;
  wire _6249 = uncoded_block[418] ^ uncoded_block[419];
  wire _6250 = _4871 ^ _6249;
  wire _6251 = uncoded_block[421] ^ uncoded_block[425];
  wire _6252 = _6251 ^ _1062;
  wire _6253 = _6250 ^ _6252;
  wire _6254 = uncoded_block[431] ^ uncoded_block[433];
  wire _6255 = uncoded_block[435] ^ uncoded_block[436];
  wire _6256 = _6254 ^ _6255;
  wire _6257 = _6256 ^ _1865;
  wire _6258 = _6253 ^ _6257;
  wire _6259 = uncoded_block[447] ^ uncoded_block[449];
  wire _6260 = _6259 ^ _4883;
  wire _6261 = uncoded_block[454] ^ uncoded_block[456];
  wire _6262 = _2645 ^ _6261;
  wire _6263 = _6260 ^ _6262;
  wire _6264 = uncoded_block[457] ^ uncoded_block[461];
  wire _6265 = _6264 ^ _4185;
  wire _6266 = uncoded_block[471] ^ uncoded_block[474];
  wire _6267 = _3416 ^ _6266;
  wire _6268 = _6265 ^ _6267;
  wire _6269 = _6263 ^ _6268;
  wire _6270 = _6258 ^ _6269;
  wire _6271 = _6248 ^ _6270;
  wire _6272 = _6226 ^ _6271;
  wire _6273 = _6178 ^ _6272;
  wire _6274 = _4895 ^ _1090;
  wire _6275 = _2658 ^ _6274;
  wire _6276 = uncoded_block[487] ^ uncoded_block[488];
  wire _6277 = uncoded_block[491] ^ uncoded_block[494];
  wire _6278 = _6276 ^ _6277;
  wire _6279 = uncoded_block[500] ^ uncoded_block[502];
  wire _6280 = _1094 ^ _6279;
  wire _6281 = _6278 ^ _6280;
  wire _6282 = _6275 ^ _6281;
  wire _6283 = uncoded_block[506] ^ uncoded_block[509];
  wire _6284 = _2671 ^ _6283;
  wire _6285 = uncoded_block[510] ^ uncoded_block[513];
  wire _6286 = uncoded_block[516] ^ uncoded_block[520];
  wire _6287 = _6285 ^ _6286;
  wire _6288 = _6284 ^ _6287;
  wire _6289 = uncoded_block[523] ^ uncoded_block[524];
  wire _6290 = uncoded_block[528] ^ uncoded_block[532];
  wire _6291 = _6289 ^ _6290;
  wire _6292 = uncoded_block[534] ^ uncoded_block[536];
  wire _6293 = uncoded_block[539] ^ uncoded_block[541];
  wire _6294 = _6292 ^ _6293;
  wire _6295 = _6291 ^ _6294;
  wire _6296 = _6288 ^ _6295;
  wire _6297 = _6282 ^ _6296;
  wire _6298 = uncoded_block[542] ^ uncoded_block[544];
  wire _6299 = _6298 ^ _1909;
  wire _6300 = uncoded_block[547] ^ uncoded_block[548];
  wire _6301 = uncoded_block[549] ^ uncoded_block[553];
  wire _6302 = _6300 ^ _6301;
  wire _6303 = _6299 ^ _6302;
  wire _6304 = uncoded_block[554] ^ uncoded_block[556];
  wire _6305 = uncoded_block[557] ^ uncoded_block[560];
  wire _6306 = _6304 ^ _6305;
  wire _6307 = _6306 ^ _3466;
  wire _6308 = _6303 ^ _6307;
  wire _6309 = uncoded_block[568] ^ uncoded_block[569];
  wire _6310 = uncoded_block[570] ^ uncoded_block[578];
  wire _6311 = _6309 ^ _6310;
  wire _6312 = uncoded_block[579] ^ uncoded_block[583];
  wire _6313 = _6312 ^ _1139;
  wire _6314 = _6311 ^ _6313;
  wire _6315 = uncoded_block[588] ^ uncoded_block[592];
  wire _6316 = uncoded_block[593] ^ uncoded_block[594];
  wire _6317 = _6315 ^ _6316;
  wire _6318 = _1142 ^ _3487;
  wire _6319 = _6317 ^ _6318;
  wire _6320 = _6314 ^ _6319;
  wire _6321 = _6308 ^ _6320;
  wire _6322 = _6297 ^ _6321;
  wire _6323 = uncoded_block[608] ^ uncoded_block[609];
  wire _6324 = _2710 ^ _6323;
  wire _6325 = uncoded_block[612] ^ uncoded_block[614];
  wire _6326 = _6325 ^ _5653;
  wire _6327 = _6324 ^ _6326;
  wire _6328 = uncoded_block[618] ^ uncoded_block[622];
  wire _6329 = _6328 ^ _1953;
  wire _6330 = uncoded_block[632] ^ uncoded_block[633];
  wire _6331 = uncoded_block[634] ^ uncoded_block[635];
  wire _6332 = _6330 ^ _6331;
  wire _6333 = _6329 ^ _6332;
  wire _6334 = _6327 ^ _6333;
  wire _6335 = uncoded_block[639] ^ uncoded_block[641];
  wire _6336 = uncoded_block[642] ^ uncoded_block[643];
  wire _6337 = _6335 ^ _6336;
  wire _6338 = uncoded_block[646] ^ uncoded_block[647];
  wire _6339 = _2729 ^ _6338;
  wire _6340 = _6337 ^ _6339;
  wire _6341 = uncoded_block[649] ^ uncoded_block[652];
  wire _6342 = uncoded_block[654] ^ uncoded_block[660];
  wire _6343 = _6341 ^ _6342;
  wire _6344 = uncoded_block[661] ^ uncoded_block[665];
  wire _6345 = _6344 ^ _309;
  wire _6346 = _6343 ^ _6345;
  wire _6347 = _6340 ^ _6346;
  wire _6348 = _6334 ^ _6347;
  wire _6349 = uncoded_block[676] ^ uncoded_block[678];
  wire _6350 = _2748 ^ _6349;
  wire _6351 = _1179 ^ _6350;
  wire _6352 = uncoded_block[679] ^ uncoded_block[680];
  wire _6353 = uncoded_block[682] ^ uncoded_block[683];
  wire _6354 = _6352 ^ _6353;
  wire _6355 = _6354 ^ _323;
  wire _6356 = _6351 ^ _6355;
  wire _6357 = uncoded_block[689] ^ uncoded_block[691];
  wire _6358 = uncoded_block[693] ^ uncoded_block[695];
  wire _6359 = _6357 ^ _6358;
  wire _6360 = uncoded_block[698] ^ uncoded_block[699];
  wire _6361 = uncoded_block[703] ^ uncoded_block[704];
  wire _6362 = _6360 ^ _6361;
  wire _6363 = _6359 ^ _6362;
  wire _6364 = uncoded_block[705] ^ uncoded_block[707];
  wire _6365 = _6364 ^ _2762;
  wire _6366 = uncoded_block[713] ^ uncoded_block[716];
  wire _6367 = uncoded_block[719] ^ uncoded_block[720];
  wire _6368 = _6366 ^ _6367;
  wire _6369 = _6365 ^ _6368;
  wire _6370 = _6363 ^ _6369;
  wire _6371 = _6356 ^ _6370;
  wire _6372 = _6348 ^ _6371;
  wire _6373 = _6322 ^ _6372;
  wire _6374 = uncoded_block[723] ^ uncoded_block[724];
  wire _6375 = uncoded_block[725] ^ uncoded_block[734];
  wire _6376 = _6374 ^ _6375;
  wire _6377 = uncoded_block[736] ^ uncoded_block[745];
  wire _6378 = uncoded_block[748] ^ uncoded_block[753];
  wire _6379 = _6377 ^ _6378;
  wire _6380 = _6376 ^ _6379;
  wire _6381 = _1215 ^ _5019;
  wire _6382 = uncoded_block[771] ^ uncoded_block[772];
  wire _6383 = _2783 ^ _6382;
  wire _6384 = _6381 ^ _6383;
  wire _6385 = _6380 ^ _6384;
  wire _6386 = uncoded_block[777] ^ uncoded_block[782];
  wire _6387 = _6386 ^ _4309;
  wire _6388 = uncoded_block[785] ^ uncoded_block[789];
  wire _6389 = _6388 ^ _1232;
  wire _6390 = _6387 ^ _6389;
  wire _6391 = uncoded_block[795] ^ uncoded_block[796];
  wire _6392 = _6391 ^ _3576;
  wire _6393 = uncoded_block[803] ^ uncoded_block[809];
  wire _6394 = _6393 ^ _5042;
  wire _6395 = _6392 ^ _6394;
  wire _6396 = _6390 ^ _6395;
  wire _6397 = _6385 ^ _6396;
  wire _6398 = uncoded_block[816] ^ uncoded_block[819];
  wire _6399 = uncoded_block[822] ^ uncoded_block[825];
  wire _6400 = _6398 ^ _6399;
  wire _6401 = uncoded_block[827] ^ uncoded_block[828];
  wire _6402 = uncoded_block[829] ^ uncoded_block[835];
  wire _6403 = _6401 ^ _6402;
  wire _6404 = _6400 ^ _6403;
  wire _6405 = _2815 ^ _5060;
  wire _6406 = uncoded_block[851] ^ uncoded_block[852];
  wire _6407 = _4340 ^ _6406;
  wire _6408 = _6405 ^ _6407;
  wire _6409 = _6404 ^ _6408;
  wire _6410 = uncoded_block[859] ^ uncoded_block[861];
  wire _6411 = _5742 ^ _6410;
  wire _6412 = uncoded_block[862] ^ uncoded_block[864];
  wire _6413 = _6412 ^ _2827;
  wire _6414 = _6411 ^ _6413;
  wire _6415 = uncoded_block[870] ^ uncoded_block[871];
  wire _6416 = uncoded_block[873] ^ uncoded_block[874];
  wire _6417 = _6415 ^ _6416;
  wire _6418 = _3608 ^ _421;
  wire _6419 = _6417 ^ _6418;
  wire _6420 = _6414 ^ _6419;
  wire _6421 = _6409 ^ _6420;
  wire _6422 = _6397 ^ _6421;
  wire _6423 = _1273 ^ _1277;
  wire _6424 = uncoded_block[899] ^ uncoded_block[901];
  wire _6425 = uncoded_block[902] ^ uncoded_block[906];
  wire _6426 = _6424 ^ _6425;
  wire _6427 = _6423 ^ _6426;
  wire _6428 = uncoded_block[909] ^ uncoded_block[910];
  wire _6429 = _1284 ^ _6428;
  wire _6430 = uncoded_block[912] ^ uncoded_block[915];
  wire _6431 = _6430 ^ _2852;
  wire _6432 = _6429 ^ _6431;
  wire _6433 = _6427 ^ _6432;
  wire _6434 = uncoded_block[918] ^ uncoded_block[922];
  wire _6435 = uncoded_block[923] ^ uncoded_block[929];
  wire _6436 = _6434 ^ _6435;
  wire _6437 = _5096 ^ _452;
  wire _6438 = _6436 ^ _6437;
  wire _6439 = uncoded_block[941] ^ uncoded_block[942];
  wire _6440 = _4375 ^ _6439;
  wire _6441 = uncoded_block[954] ^ uncoded_block[958];
  wire _6442 = _455 ^ _6441;
  wire _6443 = _6440 ^ _6442;
  wire _6444 = _6438 ^ _6443;
  wire _6445 = _6433 ^ _6444;
  wire _6446 = _1308 ^ _5783;
  wire _6447 = uncoded_block[968] ^ uncoded_block[970];
  wire _6448 = _6447 ^ _2877;
  wire _6449 = _6446 ^ _6448;
  wire _6450 = uncoded_block[978] ^ uncoded_block[982];
  wire _6451 = uncoded_block[984] ^ uncoded_block[987];
  wire _6452 = _6450 ^ _6451;
  wire _6453 = uncoded_block[995] ^ uncoded_block[996];
  wire _6454 = _1318 ^ _6453;
  wire _6455 = _6452 ^ _6454;
  wire _6456 = _6449 ^ _6455;
  wire _6457 = uncoded_block[997] ^ uncoded_block[999];
  wire _6458 = _6457 ^ _4404;
  wire _6459 = uncoded_block[1005] ^ uncoded_block[1007];
  wire _6460 = _6459 ^ _4409;
  wire _6461 = _6458 ^ _6460;
  wire _6462 = uncoded_block[1011] ^ uncoded_block[1016];
  wire _6463 = _6462 ^ _2893;
  wire _6464 = _5135 ^ _5137;
  wire _6465 = _6463 ^ _6464;
  wire _6466 = _6461 ^ _6465;
  wire _6467 = _6456 ^ _6466;
  wire _6468 = _6445 ^ _6467;
  wire _6469 = _6422 ^ _6468;
  wire _6470 = _6373 ^ _6469;
  wire _6471 = _6273 ^ _6470;
  wire _6472 = uncoded_block[1027] ^ uncoded_block[1031];
  wire _6473 = _6472 ^ _4418;
  wire _6474 = uncoded_block[1034] ^ uncoded_block[1037];
  wire _6475 = uncoded_block[1039] ^ uncoded_block[1040];
  wire _6476 = _6474 ^ _6475;
  wire _6477 = _6473 ^ _6476;
  wire _6478 = uncoded_block[1041] ^ uncoded_block[1042];
  wire _6479 = _6478 ^ _2134;
  wire _6480 = _518 ^ _3682;
  wire _6481 = _6479 ^ _6480;
  wire _6482 = _6477 ^ _6481;
  wire _6483 = uncoded_block[1059] ^ uncoded_block[1060];
  wire _6484 = _6483 ^ _2917;
  wire _6485 = uncoded_block[1065] ^ uncoded_block[1070];
  wire _6486 = uncoded_block[1076] ^ uncoded_block[1077];
  wire _6487 = _6485 ^ _6486;
  wire _6488 = _6484 ^ _6487;
  wire _6489 = _1370 ^ _534;
  wire _6490 = _536 ^ _5842;
  wire _6491 = _6489 ^ _6490;
  wire _6492 = _6488 ^ _6491;
  wire _6493 = _6482 ^ _6492;
  wire _6494 = uncoded_block[1107] ^ uncoded_block[1110];
  wire _6495 = _546 ^ _6494;
  wire _6496 = uncoded_block[1118] ^ uncoded_block[1121];
  wire _6497 = _6496 ^ _2944;
  wire _6498 = _6495 ^ _6497;
  wire _6499 = uncoded_block[1128] ^ uncoded_block[1129];
  wire _6500 = _4459 ^ _6499;
  wire _6501 = uncoded_block[1134] ^ uncoded_block[1136];
  wire _6502 = _6501 ^ _5859;
  wire _6503 = _6500 ^ _6502;
  wire _6504 = _6498 ^ _6503;
  wire _6505 = uncoded_block[1148] ^ uncoded_block[1149];
  wire _6506 = _2953 ^ _6505;
  wire _6507 = uncoded_block[1153] ^ uncoded_block[1156];
  wire _6508 = _4466 ^ _6507;
  wire _6509 = _6506 ^ _6508;
  wire _6510 = uncoded_block[1157] ^ uncoded_block[1160];
  wire _6511 = uncoded_block[1164] ^ uncoded_block[1165];
  wire _6512 = _6510 ^ _6511;
  wire _6513 = uncoded_block[1167] ^ uncoded_block[1171];
  wire _6514 = _6513 ^ _5872;
  wire _6515 = _6512 ^ _6514;
  wire _6516 = _6509 ^ _6515;
  wire _6517 = _6504 ^ _6516;
  wire _6518 = _6493 ^ _6517;
  wire _6519 = uncoded_block[1178] ^ uncoded_block[1179];
  wire _6520 = uncoded_block[1182] ^ uncoded_block[1184];
  wire _6521 = _6519 ^ _6520;
  wire _6522 = uncoded_block[1190] ^ uncoded_block[1192];
  wire _6523 = _5201 ^ _6522;
  wire _6524 = _6521 ^ _6523;
  wire _6525 = uncoded_block[1194] ^ uncoded_block[1195];
  wire _6526 = _6525 ^ _597;
  wire _6527 = _6526 ^ _2208;
  wire _6528 = _6524 ^ _6527;
  wire _6529 = uncoded_block[1203] ^ uncoded_block[1205];
  wire _6530 = uncoded_block[1206] ^ uncoded_block[1207];
  wire _6531 = _6529 ^ _6530;
  wire _6532 = uncoded_block[1222] ^ uncoded_block[1224];
  wire _6533 = _4496 ^ _6532;
  wire _6534 = _6531 ^ _6533;
  wire _6535 = uncoded_block[1225] ^ uncoded_block[1236];
  wire _6536 = uncoded_block[1240] ^ uncoded_block[1241];
  wire _6537 = _6535 ^ _6536;
  wire _6538 = uncoded_block[1245] ^ uncoded_block[1246];
  wire _6539 = _1448 ^ _6538;
  wire _6540 = _6537 ^ _6539;
  wire _6541 = _6534 ^ _6540;
  wire _6542 = _6528 ^ _6541;
  wire _6543 = uncoded_block[1249] ^ uncoded_block[1250];
  wire _6544 = _2232 ^ _6543;
  wire _6545 = uncoded_block[1251] ^ uncoded_block[1253];
  wire _6546 = uncoded_block[1254] ^ uncoded_block[1255];
  wire _6547 = _6545 ^ _6546;
  wire _6548 = _6544 ^ _6547;
  wire _6549 = _5234 ^ _3784;
  wire _6550 = uncoded_block[1264] ^ uncoded_block[1265];
  wire _6551 = _5235 ^ _6550;
  wire _6552 = _6549 ^ _6551;
  wire _6553 = _6548 ^ _6552;
  wire _6554 = uncoded_block[1269] ^ uncoded_block[1273];
  wire _6555 = _6554 ^ _630;
  wire _6556 = uncoded_block[1278] ^ uncoded_block[1281];
  wire _6557 = uncoded_block[1282] ^ uncoded_block[1283];
  wire _6558 = _6556 ^ _6557;
  wire _6559 = _6555 ^ _6558;
  wire _6560 = uncoded_block[1284] ^ uncoded_block[1285];
  wire _6561 = uncoded_block[1287] ^ uncoded_block[1291];
  wire _6562 = _6560 ^ _6561;
  wire _6563 = uncoded_block[1294] ^ uncoded_block[1297];
  wire _6564 = uncoded_block[1299] ^ uncoded_block[1300];
  wire _6565 = _6563 ^ _6564;
  wire _6566 = _6562 ^ _6565;
  wire _6567 = _6559 ^ _6566;
  wire _6568 = _6553 ^ _6567;
  wire _6569 = _6542 ^ _6568;
  wire _6570 = _6518 ^ _6569;
  wire _6571 = uncoded_block[1304] ^ uncoded_block[1306];
  wire _6572 = uncoded_block[1308] ^ uncoded_block[1309];
  wire _6573 = _6571 ^ _6572;
  wire _6574 = uncoded_block[1314] ^ uncoded_block[1317];
  wire _6575 = _3808 ^ _6574;
  wire _6576 = _6573 ^ _6575;
  wire _6577 = _4540 ^ _1487;
  wire _6578 = uncoded_block[1330] ^ uncoded_block[1332];
  wire _6579 = _4545 ^ _6578;
  wire _6580 = _6577 ^ _6579;
  wire _6581 = _6576 ^ _6580;
  wire _6582 = _5932 ^ _3822;
  wire _6583 = uncoded_block[1340] ^ uncoded_block[1344];
  wire _6584 = uncoded_block[1345] ^ uncoded_block[1353];
  wire _6585 = _6583 ^ _6584;
  wire _6586 = _6582 ^ _6585;
  wire _6587 = uncoded_block[1356] ^ uncoded_block[1357];
  wire _6588 = uncoded_block[1359] ^ uncoded_block[1360];
  wire _6589 = _6587 ^ _6588;
  wire _6590 = _5275 ^ _677;
  wire _6591 = _6589 ^ _6590;
  wire _6592 = _6586 ^ _6591;
  wire _6593 = _6581 ^ _6592;
  wire _6594 = uncoded_block[1369] ^ uncoded_block[1374];
  wire _6595 = _6594 ^ _687;
  wire _6596 = uncoded_block[1384] ^ uncoded_block[1386];
  wire _6597 = uncoded_block[1389] ^ uncoded_block[1392];
  wire _6598 = _6596 ^ _6597;
  wire _6599 = _6595 ^ _6598;
  wire _6600 = uncoded_block[1398] ^ uncoded_block[1400];
  wire _6601 = _4569 ^ _6600;
  wire _6602 = uncoded_block[1401] ^ uncoded_block[1405];
  wire _6603 = _6602 ^ _701;
  wire _6604 = _6601 ^ _6603;
  wire _6605 = _6599 ^ _6604;
  wire _6606 = uncoded_block[1409] ^ uncoded_block[1413];
  wire _6607 = uncoded_block[1417] ^ uncoded_block[1419];
  wire _6608 = _6606 ^ _6607;
  wire _6609 = uncoded_block[1420] ^ uncoded_block[1426];
  wire _6610 = _6609 ^ _5968;
  wire _6611 = _6608 ^ _6610;
  wire _6612 = _3857 ^ _3861;
  wire _6613 = uncoded_block[1442] ^ uncoded_block[1443];
  wire _6614 = _6613 ^ _5305;
  wire _6615 = _6612 ^ _6614;
  wire _6616 = _6611 ^ _6615;
  wire _6617 = _6605 ^ _6616;
  wire _6618 = _6593 ^ _6617;
  wire _6619 = uncoded_block[1446] ^ uncoded_block[1449];
  wire _6620 = uncoded_block[1450] ^ uncoded_block[1451];
  wire _6621 = _6619 ^ _6620;
  wire _6622 = uncoded_block[1454] ^ uncoded_block[1455];
  wire _6623 = uncoded_block[1456] ^ uncoded_block[1463];
  wire _6624 = _6622 ^ _6623;
  wire _6625 = _6621 ^ _6624;
  wire _6626 = _3094 ^ _3879;
  wire _6627 = uncoded_block[1473] ^ uncoded_block[1476];
  wire _6628 = _6627 ^ _3884;
  wire _6629 = _6626 ^ _6628;
  wire _6630 = _6625 ^ _6629;
  wire _6631 = uncoded_block[1494] ^ uncoded_block[1495];
  wire _6632 = _6631 ^ _743;
  wire _6633 = _3104 ^ _6632;
  wire _6634 = uncoded_block[1498] ^ uncoded_block[1499];
  wire _6635 = uncoded_block[1500] ^ uncoded_block[1503];
  wire _6636 = _6634 ^ _6635;
  wire _6637 = uncoded_block[1508] ^ uncoded_block[1510];
  wire _6638 = _3894 ^ _6637;
  wire _6639 = _6636 ^ _6638;
  wire _6640 = _6633 ^ _6639;
  wire _6641 = _6630 ^ _6640;
  wire _6642 = uncoded_block[1511] ^ uncoded_block[1514];
  wire _6643 = uncoded_block[1516] ^ uncoded_block[1518];
  wire _6644 = _6642 ^ _6643;
  wire _6645 = _4621 ^ _3123;
  wire _6646 = _6644 ^ _6645;
  wire _6647 = uncoded_block[1530] ^ uncoded_block[1532];
  wire _6648 = uncoded_block[1535] ^ uncoded_block[1536];
  wire _6649 = _6647 ^ _6648;
  wire _6650 = uncoded_block[1537] ^ uncoded_block[1538];
  wire _6651 = uncoded_block[1539] ^ uncoded_block[1540];
  wire _6652 = _6650 ^ _6651;
  wire _6653 = _6649 ^ _6652;
  wire _6654 = _6646 ^ _6653;
  wire _6655 = uncoded_block[1546] ^ uncoded_block[1551];
  wire _6656 = _1590 ^ _6655;
  wire _6657 = uncoded_block[1552] ^ uncoded_block[1553];
  wire _6658 = _6657 ^ _770;
  wire _6659 = _6656 ^ _6658;
  wire _6660 = uncoded_block[1559] ^ uncoded_block[1568];
  wire _6661 = uncoded_block[1569] ^ uncoded_block[1572];
  wire _6662 = _6660 ^ _6661;
  wire _6663 = uncoded_block[1577] ^ uncoded_block[1578];
  wire _6664 = _4648 ^ _6663;
  wire _6665 = _6662 ^ _6664;
  wire _6666 = _6659 ^ _6665;
  wire _6667 = _6654 ^ _6666;
  wire _6668 = _6641 ^ _6667;
  wire _6669 = _6618 ^ _6668;
  wire _6670 = _6570 ^ _6669;
  wire _6671 = uncoded_block[1580] ^ uncoded_block[1586];
  wire _6672 = _6671 ^ _789;
  wire _6673 = uncoded_block[1593] ^ uncoded_block[1594];
  wire _6674 = uncoded_block[1596] ^ uncoded_block[1599];
  wire _6675 = _6673 ^ _6674;
  wire _6676 = _6672 ^ _6675;
  wire _6677 = uncoded_block[1606] ^ uncoded_block[1608];
  wire _6678 = _6677 ^ _801;
  wire _6679 = uncoded_block[1614] ^ uncoded_block[1615];
  wire _6680 = uncoded_block[1616] ^ uncoded_block[1618];
  wire _6681 = _6679 ^ _6680;
  wire _6682 = _6678 ^ _6681;
  wire _6683 = _6676 ^ _6682;
  wire _6684 = uncoded_block[1621] ^ uncoded_block[1623];
  wire _6685 = uncoded_block[1624] ^ uncoded_block[1629];
  wire _6686 = _6684 ^ _6685;
  wire _6687 = _5388 ^ _2405;
  wire _6688 = _6686 ^ _6687;
  wire _6689 = uncoded_block[1640] ^ uncoded_block[1641];
  wire _6690 = _5392 ^ _6689;
  wire _6691 = uncoded_block[1647] ^ uncoded_block[1649];
  wire _6692 = _6691 ^ _4677;
  wire _6693 = _6690 ^ _6692;
  wire _6694 = _6688 ^ _6693;
  wire _6695 = _6683 ^ _6694;
  wire _6696 = uncoded_block[1655] ^ uncoded_block[1658];
  wire _6697 = _4678 ^ _6696;
  wire _6698 = _4680 ^ _5399;
  wire _6699 = _6697 ^ _6698;
  wire _6700 = uncoded_block[1672] ^ uncoded_block[1673];
  wire _6701 = _3182 ^ _6700;
  wire _6702 = _830 ^ _832;
  wire _6703 = _6701 ^ _6702;
  wire _6704 = _6699 ^ _6703;
  wire _6705 = uncoded_block[1685] ^ uncoded_block[1687];
  wire _6706 = _833 ^ _6705;
  wire _6707 = uncoded_block[1691] ^ uncoded_block[1692];
  wire _6708 = _837 ^ _6707;
  wire _6709 = _6706 ^ _6708;
  wire _6710 = uncoded_block[1694] ^ uncoded_block[1697];
  wire _6711 = uncoded_block[1698] ^ uncoded_block[1702];
  wire _6712 = _6710 ^ _6711;
  wire _6713 = uncoded_block[1710] ^ uncoded_block[1716];
  wire _6714 = _2435 ^ _6713;
  wire _6715 = _6712 ^ _6714;
  wire _6716 = _6709 ^ _6715;
  wire _6717 = _6704 ^ _6716;
  wire _6718 = _6695 ^ _6717;
  wire _6719 = uncoded_block[1718] ^ uncoded_block[1721];
  wire _6720 = _6719 ^ uncoded_block[1722];
  wire _6721 = _6718 ^ _6720;
  wire _6722 = _6670 ^ _6721;
  wire _6723 = _6471 ^ _6722;
  wire _6724 = uncoded_block[7] ^ uncoded_block[8];
  wire _6725 = _4712 ^ _6724;
  wire _6726 = _4711 ^ _6725;
  wire _6727 = _3213 ^ _5423;
  wire _6728 = uncoded_block[26] ^ uncoded_block[29];
  wire _6729 = _4716 ^ _6728;
  wire _6730 = _6727 ^ _6729;
  wire _6731 = _6726 ^ _6730;
  wire _6732 = uncoded_block[34] ^ uncoded_block[37];
  wire _6733 = _3225 ^ _6732;
  wire _6734 = _2466 ^ _4008;
  wire _6735 = _6733 ^ _6734;
  wire _6736 = uncoded_block[43] ^ uncoded_block[45];
  wire _6737 = _6736 ^ _885;
  wire _6738 = _886 ^ _1703;
  wire _6739 = _6737 ^ _6738;
  wire _6740 = _6735 ^ _6739;
  wire _6741 = _6731 ^ _6740;
  wire _6742 = uncoded_block[60] ^ uncoded_block[63];
  wire _6743 = _26 ^ _6742;
  wire _6744 = uncoded_block[66] ^ uncoded_block[68];
  wire _6745 = uncoded_block[69] ^ uncoded_block[72];
  wire _6746 = _6744 ^ _6745;
  wire _6747 = _6743 ^ _6746;
  wire _6748 = _4733 ^ _1712;
  wire _6749 = uncoded_block[79] ^ uncoded_block[80];
  wire _6750 = uncoded_block[81] ^ uncoded_block[82];
  wire _6751 = _6749 ^ _6750;
  wire _6752 = _6748 ^ _6751;
  wire _6753 = _6747 ^ _6752;
  wire _6754 = uncoded_block[83] ^ uncoded_block[86];
  wire _6755 = uncoded_block[87] ^ uncoded_block[88];
  wire _6756 = _6754 ^ _6755;
  wire _6757 = uncoded_block[89] ^ uncoded_block[93];
  wire _6758 = uncoded_block[95] ^ uncoded_block[97];
  wire _6759 = _6757 ^ _6758;
  wire _6760 = _6756 ^ _6759;
  wire _6761 = _910 ^ _1721;
  wire _6762 = uncoded_block[106] ^ uncoded_block[111];
  wire _6763 = uncoded_block[112] ^ uncoded_block[113];
  wire _6764 = _6762 ^ _6763;
  wire _6765 = _6761 ^ _6764;
  wire _6766 = _6760 ^ _6765;
  wire _6767 = _6753 ^ _6766;
  wire _6768 = _6741 ^ _6767;
  wire _6769 = uncoded_block[114] ^ uncoded_block[116];
  wire _6770 = _6769 ^ _4750;
  wire _6771 = uncoded_block[120] ^ uncoded_block[125];
  wire _6772 = _6771 ^ _4753;
  wire _6773 = _6770 ^ _6772;
  wire _6774 = uncoded_block[128] ^ uncoded_block[130];
  wire _6775 = _6774 ^ _924;
  wire _6776 = uncoded_block[139] ^ uncoded_block[141];
  wire _6777 = _2510 ^ _6776;
  wire _6778 = _6775 ^ _6777;
  wire _6779 = _6773 ^ _6778;
  wire _6780 = uncoded_block[147] ^ uncoded_block[148];
  wire _6781 = _2511 ^ _6780;
  wire _6782 = _70 ^ _5469;
  wire _6783 = _6781 ^ _6782;
  wire _6784 = uncoded_block[155] ^ uncoded_block[158];
  wire _6785 = uncoded_block[161] ^ uncoded_block[163];
  wire _6786 = _6784 ^ _6785;
  wire _6787 = uncoded_block[165] ^ uncoded_block[167];
  wire _6788 = uncoded_block[168] ^ uncoded_block[169];
  wire _6789 = _6787 ^ _6788;
  wire _6790 = _6786 ^ _6789;
  wire _6791 = _6783 ^ _6790;
  wire _6792 = _6779 ^ _6791;
  wire _6793 = _81 ^ _2522;
  wire _6794 = uncoded_block[177] ^ uncoded_block[182];
  wire _6795 = _6794 ^ _944;
  wire _6796 = _6793 ^ _6795;
  wire _6797 = uncoded_block[186] ^ uncoded_block[190];
  wire _6798 = uncoded_block[191] ^ uncoded_block[192];
  wire _6799 = _6797 ^ _6798;
  wire _6800 = uncoded_block[194] ^ uncoded_block[197];
  wire _6801 = uncoded_block[198] ^ uncoded_block[199];
  wire _6802 = _6800 ^ _6801;
  wire _6803 = _6799 ^ _6802;
  wire _6804 = _6796 ^ _6803;
  wire _6805 = uncoded_block[201] ^ uncoded_block[202];
  wire _6806 = uncoded_block[205] ^ uncoded_block[207];
  wire _6807 = _6805 ^ _6806;
  wire _6808 = uncoded_block[208] ^ uncoded_block[212];
  wire _6809 = _6808 ^ _959;
  wire _6810 = _6807 ^ _6809;
  wire _6811 = uncoded_block[215] ^ uncoded_block[219];
  wire _6812 = uncoded_block[220] ^ uncoded_block[222];
  wire _6813 = _6811 ^ _6812;
  wire _6814 = uncoded_block[226] ^ uncoded_block[228];
  wire _6815 = _2545 ^ _6814;
  wire _6816 = _6813 ^ _6815;
  wire _6817 = _6810 ^ _6816;
  wire _6818 = _6804 ^ _6817;
  wire _6819 = _6792 ^ _6818;
  wire _6820 = _6768 ^ _6819;
  wire _6821 = uncoded_block[229] ^ uncoded_block[231];
  wire _6822 = uncoded_block[234] ^ uncoded_block[236];
  wire _6823 = _6821 ^ _6822;
  wire _6824 = uncoded_block[237] ^ uncoded_block[240];
  wire _6825 = _6824 ^ _5503;
  wire _6826 = _6823 ^ _6825;
  wire _6827 = _6179 ^ _4087;
  wire _6828 = _1786 ^ _4095;
  wire _6829 = _6827 ^ _6828;
  wire _6830 = _6826 ^ _6829;
  wire _6831 = uncoded_block[262] ^ uncoded_block[264];
  wire _6832 = _6831 ^ _4099;
  wire _6833 = uncoded_block[275] ^ uncoded_block[276];
  wire _6834 = uncoded_block[277] ^ uncoded_block[281];
  wire _6835 = _6833 ^ _6834;
  wire _6836 = _6832 ^ _6835;
  wire _6837 = uncoded_block[286] ^ uncoded_block[289];
  wire _6838 = uncoded_block[290] ^ uncoded_block[293];
  wire _6839 = _6837 ^ _6838;
  wire _6840 = _137 ^ _1807;
  wire _6841 = _6839 ^ _6840;
  wire _6842 = _6836 ^ _6841;
  wire _6843 = _6830 ^ _6842;
  wire _6844 = _142 ^ _4826;
  wire _6845 = uncoded_block[305] ^ uncoded_block[306];
  wire _6846 = uncoded_block[309] ^ uncoded_block[313];
  wire _6847 = _6845 ^ _6846;
  wire _6848 = _6844 ^ _6847;
  wire _6849 = uncoded_block[315] ^ uncoded_block[319];
  wire _6850 = uncoded_block[320] ^ uncoded_block[321];
  wire _6851 = _6849 ^ _6850;
  wire _6852 = uncoded_block[322] ^ uncoded_block[326];
  wire _6853 = uncoded_block[329] ^ uncoded_block[333];
  wire _6854 = _6852 ^ _6853;
  wire _6855 = _6851 ^ _6854;
  wire _6856 = _6848 ^ _6855;
  wire _6857 = uncoded_block[335] ^ uncoded_block[336];
  wire _6858 = _6857 ^ _1018;
  wire _6859 = uncoded_block[342] ^ uncoded_block[345];
  wire _6860 = uncoded_block[348] ^ uncoded_block[352];
  wire _6861 = _6859 ^ _6860;
  wire _6862 = _6858 ^ _6861;
  wire _6863 = uncoded_block[353] ^ uncoded_block[357];
  wire _6864 = uncoded_block[358] ^ uncoded_block[359];
  wire _6865 = _6863 ^ _6864;
  wire _6866 = uncoded_block[360] ^ uncoded_block[363];
  wire _6867 = uncoded_block[364] ^ uncoded_block[370];
  wire _6868 = _6866 ^ _6867;
  wire _6869 = _6865 ^ _6868;
  wire _6870 = _6862 ^ _6869;
  wire _6871 = _6856 ^ _6870;
  wire _6872 = _6843 ^ _6871;
  wire _6873 = uncoded_block[371] ^ uncoded_block[372];
  wire _6874 = uncoded_block[374] ^ uncoded_block[378];
  wire _6875 = _6873 ^ _6874;
  wire _6876 = uncoded_block[382] ^ uncoded_block[383];
  wire _6877 = _6876 ^ _3380;
  wire _6878 = _6875 ^ _6877;
  wire _6879 = uncoded_block[391] ^ uncoded_block[393];
  wire _6880 = _176 ^ _6879;
  wire _6881 = uncoded_block[394] ^ uncoded_block[396];
  wire _6882 = _6881 ^ _1048;
  wire _6883 = _6880 ^ _6882;
  wire _6884 = _6878 ^ _6883;
  wire _6885 = _181 ^ _6244;
  wire _6886 = _190 ^ _4871;
  wire _6887 = _6885 ^ _6886;
  wire _6888 = _6249 ^ _4163;
  wire _6889 = uncoded_block[422] ^ uncoded_block[425];
  wire _6890 = _6889 ^ _1062;
  wire _6891 = _6888 ^ _6890;
  wire _6892 = _6887 ^ _6891;
  wire _6893 = _6884 ^ _6892;
  wire _6894 = uncoded_block[428] ^ uncoded_block[429];
  wire _6895 = _6894 ^ _2638;
  wire _6896 = _201 ^ _2641;
  wire _6897 = _6895 ^ _6896;
  wire _6898 = uncoded_block[442] ^ uncoded_block[445];
  wire _6899 = _6898 ^ _1069;
  wire _6900 = uncoded_block[450] ^ uncoded_block[453];
  wire _6901 = _6900 ^ _2650;
  wire _6902 = _6899 ^ _6901;
  wire _6903 = _6897 ^ _6902;
  wire _6904 = uncoded_block[460] ^ uncoded_block[465];
  wire _6905 = _3415 ^ _6904;
  wire _6906 = uncoded_block[469] ^ uncoded_block[471];
  wire _6907 = _3416 ^ _6906;
  wire _6908 = _6905 ^ _6907;
  wire _6909 = uncoded_block[474] ^ uncoded_block[482];
  wire _6910 = _4188 ^ _6909;
  wire _6911 = uncoded_block[483] ^ uncoded_block[490];
  wire _6912 = _6911 ^ _6277;
  wire _6913 = _6910 ^ _6912;
  wire _6914 = _6908 ^ _6913;
  wire _6915 = _6903 ^ _6914;
  wire _6916 = _6893 ^ _6915;
  wire _6917 = _6872 ^ _6916;
  wire _6918 = _6820 ^ _6917;
  wire _6919 = uncoded_block[495] ^ uncoded_block[497];
  wire _6920 = _6919 ^ _6279;
  wire _6921 = uncoded_block[503] ^ uncoded_block[504];
  wire _6922 = uncoded_block[505] ^ uncoded_block[508];
  wire _6923 = _6921 ^ _6922;
  wire _6924 = _6920 ^ _6923;
  wire _6925 = uncoded_block[510] ^ uncoded_block[515];
  wire _6926 = _6925 ^ _4208;
  wire _6927 = _6926 ^ _1109;
  wire _6928 = _6924 ^ _6927;
  wire _6929 = uncoded_block[528] ^ uncoded_block[529];
  wire _6930 = _1110 ^ _6929;
  wire _6931 = uncoded_block[531] ^ uncoded_block[533];
  wire _6932 = uncoded_block[535] ^ uncoded_block[536];
  wire _6933 = _6931 ^ _6932;
  wire _6934 = _6930 ^ _6933;
  wire _6935 = _1115 ^ _6298;
  wire _6936 = _246 ^ _6304;
  wire _6937 = _6935 ^ _6936;
  wire _6938 = _6934 ^ _6937;
  wire _6939 = _6928 ^ _6938;
  wire _6940 = uncoded_block[557] ^ uncoded_block[559];
  wire _6941 = _6940 ^ _5633;
  wire _6942 = uncoded_block[570] ^ uncoded_block[571];
  wire _6943 = _3467 ^ _6942;
  wire _6944 = _6941 ^ _6943;
  wire _6945 = uncoded_block[573] ^ uncoded_block[575];
  wire _6946 = _6945 ^ _263;
  wire _6947 = uncoded_block[580] ^ uncoded_block[581];
  wire _6948 = uncoded_block[583] ^ uncoded_block[588];
  wire _6949 = _6947 ^ _6948;
  wire _6950 = _6946 ^ _6949;
  wire _6951 = _6944 ^ _6950;
  wire _6952 = uncoded_block[595] ^ uncoded_block[597];
  wire _6953 = _6952 ^ _3487;
  wire _6954 = uncoded_block[603] ^ uncoded_block[607];
  wire _6955 = _6954 ^ _6323;
  wire _6956 = _6953 ^ _6955;
  wire _6957 = uncoded_block[610] ^ uncoded_block[612];
  wire _6958 = _6957 ^ _280;
  wire _6959 = uncoded_block[617] ^ uncoded_block[618];
  wire _6960 = uncoded_block[619] ^ uncoded_block[620];
  wire _6961 = _6959 ^ _6960;
  wire _6962 = _6958 ^ _6961;
  wire _6963 = _6956 ^ _6962;
  wire _6964 = _6951 ^ _6963;
  wire _6965 = _6939 ^ _6964;
  wire _6966 = uncoded_block[627] ^ uncoded_block[628];
  wire _6967 = _286 ^ _6966;
  wire _6968 = uncoded_block[629] ^ uncoded_block[636];
  wire _6969 = uncoded_block[638] ^ uncoded_block[641];
  wire _6970 = _6968 ^ _6969;
  wire _6971 = _6967 ^ _6970;
  wire _6972 = _6336 ^ _1164;
  wire _6973 = uncoded_block[648] ^ uncoded_block[651];
  wire _6974 = uncoded_block[652] ^ uncoded_block[654];
  wire _6975 = _6973 ^ _6974;
  wire _6976 = _6972 ^ _6975;
  wire _6977 = _6971 ^ _6976;
  wire _6978 = uncoded_block[669] ^ uncoded_block[675];
  wire _6979 = _308 ^ _6978;
  wire _6980 = uncoded_block[676] ^ uncoded_block[681];
  wire _6981 = _6980 ^ _3526;
  wire _6982 = _6979 ^ _6981;
  wire _6983 = uncoded_block[686] ^ uncoded_block[687];
  wire _6984 = _6983 ^ _2751;
  wire _6985 = uncoded_block[693] ^ uncoded_block[694];
  wire _6986 = _326 ^ _6985;
  wire _6987 = _6984 ^ _6986;
  wire _6988 = _6982 ^ _6987;
  wire _6989 = _6977 ^ _6988;
  wire _6990 = uncoded_block[695] ^ uncoded_block[697];
  wire _6991 = _6990 ^ _6360;
  wire _6992 = uncoded_block[701] ^ uncoded_block[702];
  wire _6993 = _6992 ^ _5685;
  wire _6994 = _6991 ^ _6993;
  wire _6995 = _3536 ^ _2763;
  wire _6996 = _4997 ^ _6995;
  wire _6997 = _6994 ^ _6996;
  wire _6998 = uncoded_block[719] ^ uncoded_block[723];
  wire _6999 = uncoded_block[725] ^ uncoded_block[727];
  wire _7000 = _6998 ^ _6999;
  wire _7001 = uncoded_block[728] ^ uncoded_block[729];
  wire _7002 = uncoded_block[732] ^ uncoded_block[733];
  wire _7003 = _7001 ^ _7002;
  wire _7004 = _7000 ^ _7003;
  wire _7005 = uncoded_block[737] ^ uncoded_block[738];
  wire _7006 = uncoded_block[741] ^ uncoded_block[743];
  wire _7007 = _7005 ^ _7006;
  wire _7008 = _7007 ^ _5014;
  wire _7009 = _7004 ^ _7008;
  wire _7010 = _6997 ^ _7009;
  wire _7011 = _6989 ^ _7010;
  wire _7012 = _6965 ^ _7011;
  wire _7013 = uncoded_block[753] ^ uncoded_block[754];
  wire _7014 = _4295 ^ _7013;
  wire _7015 = uncoded_block[755] ^ uncoded_block[757];
  wire _7016 = uncoded_block[760] ^ uncoded_block[763];
  wire _7017 = _7015 ^ _7016;
  wire _7018 = _7014 ^ _7017;
  wire _7019 = uncoded_block[772] ^ uncoded_block[775];
  wire _7020 = _5709 ^ _7019;
  wire _7021 = uncoded_block[778] ^ uncoded_block[780];
  wire _7022 = _7021 ^ _2794;
  wire _7023 = _7020 ^ _7022;
  wire _7024 = _7018 ^ _7023;
  wire _7025 = _2795 ^ _4311;
  wire _7026 = uncoded_block[793] ^ uncoded_block[798];
  wire _7027 = _374 ^ _7026;
  wire _7028 = _7025 ^ _7027;
  wire _7029 = uncoded_block[799] ^ uncoded_block[800];
  wire _7030 = uncoded_block[802] ^ uncoded_block[806];
  wire _7031 = _7029 ^ _7030;
  wire _7032 = uncoded_block[808] ^ uncoded_block[815];
  wire _7033 = _7032 ^ _4325;
  wire _7034 = _7031 ^ _7033;
  wire _7035 = _7028 ^ _7034;
  wire _7036 = _7024 ^ _7035;
  wire _7037 = uncoded_block[821] ^ uncoded_block[822];
  wire _7038 = _1242 ^ _7037;
  wire _7039 = uncoded_block[829] ^ uncoded_block[830];
  wire _7040 = _6401 ^ _7039;
  wire _7041 = _7038 ^ _7040;
  wire _7042 = _4331 ^ _4336;
  wire _7043 = uncoded_block[838] ^ uncoded_block[840];
  wire _7044 = _7043 ^ _2036;
  wire _7045 = _7042 ^ _7044;
  wire _7046 = _7041 ^ _7045;
  wire _7047 = uncoded_block[845] ^ uncoded_block[847];
  wire _7048 = _1256 ^ _7047;
  wire _7049 = uncoded_block[854] ^ uncoded_block[856];
  wire _7050 = _2044 ^ _7049;
  wire _7051 = _7048 ^ _7050;
  wire _7052 = uncoded_block[857] ^ uncoded_block[861];
  wire _7053 = _7052 ^ _5069;
  wire _7054 = uncoded_block[867] ^ uncoded_block[869];
  wire _7055 = _7054 ^ _6415;
  wire _7056 = _7053 ^ _7055;
  wire _7057 = _7051 ^ _7056;
  wire _7058 = _7046 ^ _7057;
  wire _7059 = _7036 ^ _7058;
  wire _7060 = uncoded_block[877] ^ uncoded_block[880];
  wire _7061 = _417 ^ _7060;
  wire _7062 = uncoded_block[882] ^ uncoded_block[883];
  wire _7063 = _7062 ^ _423;
  wire _7064 = _7061 ^ _7063;
  wire _7065 = _4354 ^ _5083;
  wire _7066 = uncoded_block[899] ^ uncoded_block[903];
  wire _7067 = _428 ^ _7066;
  wire _7068 = _7065 ^ _7067;
  wire _7069 = _7064 ^ _7068;
  wire _7070 = uncoded_block[906] ^ uncoded_block[908];
  wire _7071 = _7070 ^ _6428;
  wire _7072 = _7071 ^ _2853;
  wire _7073 = uncoded_block[919] ^ uncoded_block[924];
  wire _7074 = _7073 ^ _4370;
  wire _7075 = uncoded_block[928] ^ uncoded_block[930];
  wire _7076 = _7075 ^ _3637;
  wire _7077 = _7074 ^ _7076;
  wire _7078 = _7072 ^ _7077;
  wire _7079 = _7069 ^ _7078;
  wire _7080 = uncoded_block[938] ^ uncoded_block[939];
  wire _7081 = _2079 ^ _7080;
  wire _7082 = uncoded_block[941] ^ uncoded_block[951];
  wire _7083 = uncoded_block[953] ^ uncoded_block[957];
  wire _7084 = _7082 ^ _7083;
  wire _7085 = _7081 ^ _7084;
  wire _7086 = uncoded_block[961] ^ uncoded_block[964];
  wire _7087 = _7086 ^ _2092;
  wire _7088 = uncoded_block[969] ^ uncoded_block[970];
  wire _7089 = _2093 ^ _7088;
  wire _7090 = _7087 ^ _7089;
  wire _7091 = _7085 ^ _7090;
  wire _7092 = _5112 ^ _5789;
  wire _7093 = uncoded_block[984] ^ uncoded_block[985];
  wire _7094 = uncoded_block[987] ^ uncoded_block[990];
  wire _7095 = _7093 ^ _7094;
  wire _7096 = _7092 ^ _7095;
  wire _7097 = uncoded_block[993] ^ uncoded_block[1001];
  wire _7098 = _7097 ^ _4404;
  wire _7099 = _2886 ^ _1330;
  wire _7100 = _7098 ^ _7099;
  wire _7101 = _7096 ^ _7100;
  wire _7102 = _7091 ^ _7101;
  wire _7103 = _7079 ^ _7102;
  wire _7104 = _7059 ^ _7103;
  wire _7105 = _7012 ^ _7104;
  wire _7106 = _6918 ^ _7105;
  wire _7107 = uncoded_block[1014] ^ uncoded_block[1017];
  wire _7108 = uncoded_block[1020] ^ uncoded_block[1022];
  wire _7109 = _7107 ^ _7108;
  wire _7110 = uncoded_block[1023] ^ uncoded_block[1029];
  wire _7111 = _7110 ^ _499;
  wire _7112 = _7109 ^ _7111;
  wire _7113 = _2127 ^ _6475;
  wire _7114 = _512 ^ _1356;
  wire _7115 = _7113 ^ _7114;
  wire _7116 = _7112 ^ _7115;
  wire _7117 = uncoded_block[1057] ^ uncoded_block[1058];
  wire _7118 = _5147 ^ _7117;
  wire _7119 = uncoded_block[1060] ^ uncoded_block[1068];
  wire _7120 = uncoded_block[1069] ^ uncoded_block[1077];
  wire _7121 = _7119 ^ _7120;
  wire _7122 = _7118 ^ _7121;
  wire _7123 = _5162 ^ _530;
  wire _7124 = uncoded_block[1087] ^ uncoded_block[1092];
  wire _7125 = _1371 ^ _7124;
  wire _7126 = _7123 ^ _7125;
  wire _7127 = _7122 ^ _7126;
  wire _7128 = _7116 ^ _7127;
  wire _7129 = uncoded_block[1093] ^ uncoded_block[1096];
  wire _7130 = _7129 ^ _5169;
  wire _7131 = _7130 ^ _3709;
  wire _7132 = uncoded_block[1110] ^ uncoded_block[1111];
  wire _7133 = uncoded_block[1113] ^ uncoded_block[1114];
  wire _7134 = _7132 ^ _7133;
  wire _7135 = _553 ^ _2942;
  wire _7136 = _7134 ^ _7135;
  wire _7137 = _7131 ^ _7136;
  wire _7138 = _1392 ^ _560;
  wire _7139 = _3721 ^ _5859;
  wire _7140 = _7138 ^ _7139;
  wire _7141 = uncoded_block[1144] ^ uncoded_block[1147];
  wire _7142 = _7141 ^ _6505;
  wire _7143 = uncoded_block[1150] ^ uncoded_block[1152];
  wire _7144 = _7143 ^ _2186;
  wire _7145 = _7142 ^ _7144;
  wire _7146 = _7140 ^ _7145;
  wire _7147 = _7137 ^ _7146;
  wire _7148 = _7128 ^ _7147;
  wire _7149 = uncoded_block[1160] ^ uncoded_block[1163];
  wire _7150 = _5190 ^ _7149;
  wire _7151 = uncoded_block[1165] ^ uncoded_block[1168];
  wire _7152 = _7151 ^ _1408;
  wire _7153 = _7150 ^ _7152;
  wire _7154 = uncoded_block[1171] ^ uncoded_block[1172];
  wire _7155 = _7154 ^ _2967;
  wire _7156 = _5200 ^ _2201;
  wire _7157 = _7155 ^ _7156;
  wire _7158 = _7153 ^ _7157;
  wire _7159 = uncoded_block[1191] ^ uncoded_block[1194];
  wire _7160 = uncoded_block[1197] ^ uncoded_block[1199];
  wire _7161 = _7159 ^ _7160;
  wire _7162 = uncoded_block[1200] ^ uncoded_block[1201];
  wire _7163 = uncoded_block[1202] ^ uncoded_block[1204];
  wire _7164 = _7162 ^ _7163;
  wire _7165 = _7161 ^ _7164;
  wire _7166 = uncoded_block[1208] ^ uncoded_block[1212];
  wire _7167 = _7166 ^ _605;
  wire _7168 = uncoded_block[1222] ^ uncoded_block[1223];
  wire _7169 = uncoded_block[1229] ^ uncoded_block[1233];
  wire _7170 = _7168 ^ _7169;
  wire _7171 = _7167 ^ _7170;
  wire _7172 = _7165 ^ _7171;
  wire _7173 = _7158 ^ _7172;
  wire _7174 = uncoded_block[1236] ^ uncoded_block[1238];
  wire _7175 = _1442 ^ _7174;
  wire _7176 = _2994 ^ _2997;
  wire _7177 = _7175 ^ _7176;
  wire _7178 = uncoded_block[1261] ^ uncoded_block[1264];
  wire _7179 = uncoded_block[1268] ^ uncoded_block[1270];
  wire _7180 = _7178 ^ _7179;
  wire _7181 = _5903 ^ _7180;
  wire _7182 = _7177 ^ _7181;
  wire _7183 = uncoded_block[1278] ^ uncoded_block[1280];
  wire _7184 = _7183 ^ _4525;
  wire _7185 = _4524 ^ _7184;
  wire _7186 = _3797 ^ _5913;
  wire _7187 = _4529 ^ _3800;
  wire _7188 = _7186 ^ _7187;
  wire _7189 = _7185 ^ _7188;
  wire _7190 = _7182 ^ _7189;
  wire _7191 = _7173 ^ _7190;
  wire _7192 = _7148 ^ _7191;
  wire _7193 = uncoded_block[1293] ^ uncoded_block[1295];
  wire _7194 = uncoded_block[1296] ^ uncoded_block[1299];
  wire _7195 = _7193 ^ _7194;
  wire _7196 = uncoded_block[1304] ^ uncoded_block[1310];
  wire _7197 = uncoded_block[1311] ^ uncoded_block[1317];
  wire _7198 = _7196 ^ _7197;
  wire _7199 = _7195 ^ _7198;
  wire _7200 = _3028 ^ _4543;
  wire _7201 = uncoded_block[1325] ^ uncoded_block[1327];
  wire _7202 = _7201 ^ _1490;
  wire _7203 = _7200 ^ _7202;
  wire _7204 = _7199 ^ _7203;
  wire _7205 = uncoded_block[1334] ^ uncoded_block[1341];
  wire _7206 = uncoded_block[1344] ^ uncoded_block[1347];
  wire _7207 = _7205 ^ _7206;
  wire _7208 = _669 ^ _3042;
  wire _7209 = _7207 ^ _7208;
  wire _7210 = _5272 ^ _673;
  wire _7211 = uncoded_block[1363] ^ uncoded_block[1365];
  wire _7212 = _5275 ^ _7211;
  wire _7213 = _7210 ^ _7212;
  wire _7214 = _7209 ^ _7213;
  wire _7215 = _7204 ^ _7214;
  wire _7216 = uncoded_block[1366] ^ uncoded_block[1375];
  wire _7217 = uncoded_block[1376] ^ uncoded_block[1379];
  wire _7218 = _7216 ^ _7217;
  wire _7219 = uncoded_block[1380] ^ uncoded_block[1381];
  wire _7220 = _7219 ^ _3835;
  wire _7221 = _7218 ^ _7220;
  wire _7222 = uncoded_block[1386] ^ uncoded_block[1387];
  wire _7223 = _7222 ^ _1513;
  wire _7224 = _7223 ^ _4570;
  wire _7225 = _7221 ^ _7224;
  wire _7226 = _4571 ^ _5955;
  wire _7227 = _3066 ^ _4578;
  wire _7228 = _7226 ^ _7227;
  wire _7229 = uncoded_block[1410] ^ uncoded_block[1412];
  wire _7230 = _2300 ^ _7229;
  wire _7231 = _705 ^ _1526;
  wire _7232 = _7230 ^ _7231;
  wire _7233 = _7228 ^ _7232;
  wire _7234 = _7225 ^ _7233;
  wire _7235 = _7215 ^ _7234;
  wire _7236 = _2308 ^ _5299;
  wire _7237 = uncoded_block[1434] ^ uncoded_block[1437];
  wire _7238 = uncoded_block[1438] ^ uncoded_block[1453];
  wire _7239 = _7237 ^ _7238;
  wire _7240 = _7236 ^ _7239;
  wire _7241 = uncoded_block[1458] ^ uncoded_block[1460];
  wire _7242 = _3868 ^ _7241;
  wire _7243 = uncoded_block[1461] ^ uncoded_block[1464];
  wire _7244 = _7243 ^ _1548;
  wire _7245 = _7242 ^ _7244;
  wire _7246 = _7240 ^ _7245;
  wire _7247 = uncoded_block[1468] ^ uncoded_block[1469];
  wire _7248 = _7247 ^ _4603;
  wire _7249 = _735 ^ _3884;
  wire _7250 = _7248 ^ _7249;
  wire _7251 = uncoded_block[1487] ^ uncoded_block[1489];
  wire _7252 = _3885 ^ _7251;
  wire _7253 = _3103 ^ _1565;
  wire _7254 = _7252 ^ _7253;
  wire _7255 = _7250 ^ _7254;
  wire _7256 = _7246 ^ _7255;
  wire _7257 = _743 ^ _6634;
  wire _7258 = uncoded_block[1500] ^ uncoded_block[1502];
  wire _7259 = uncoded_block[1504] ^ uncoded_block[1505];
  wire _7260 = _7258 ^ _7259;
  wire _7261 = _7257 ^ _7260;
  wire _7262 = uncoded_block[1506] ^ uncoded_block[1508];
  wire _7263 = _7262 ^ _5334;
  wire _7264 = uncoded_block[1512] ^ uncoded_block[1515];
  wire _7265 = uncoded_block[1517] ^ uncoded_block[1518];
  wire _7266 = _7264 ^ _7265;
  wire _7267 = _7263 ^ _7266;
  wire _7268 = _7261 ^ _7267;
  wire _7269 = uncoded_block[1521] ^ uncoded_block[1522];
  wire _7270 = uncoded_block[1531] ^ uncoded_block[1537];
  wire _7271 = _7269 ^ _7270;
  wire _7272 = _6651 ^ _6008;
  wire _7273 = _7271 ^ _7272;
  wire _7274 = uncoded_block[1544] ^ uncoded_block[1546];
  wire _7275 = uncoded_block[1547] ^ uncoded_block[1549];
  wire _7276 = _7274 ^ _7275;
  wire _7277 = uncoded_block[1550] ^ uncoded_block[1552];
  wire _7278 = _7277 ^ _5358;
  wire _7279 = _7276 ^ _7278;
  wire _7280 = _7273 ^ _7279;
  wire _7281 = _7268 ^ _7280;
  wire _7282 = _7256 ^ _7281;
  wire _7283 = _7235 ^ _7282;
  wire _7284 = _7192 ^ _7283;
  wire _7285 = uncoded_block[1568] ^ uncoded_block[1571];
  wire _7286 = _776 ^ _7285;
  wire _7287 = _3915 ^ _7286;
  wire _7288 = _4648 ^ _2383;
  wire _7289 = _2384 ^ _2386;
  wire _7290 = _7288 ^ _7289;
  wire _7291 = _7287 ^ _7290;
  wire _7292 = uncoded_block[1587] ^ uncoded_block[1595];
  wire _7293 = _7292 ^ _1620;
  wire _7294 = uncoded_block[1604] ^ uncoded_block[1611];
  wire _7295 = _3151 ^ _7294;
  wire _7296 = _7293 ^ _7295;
  wire _7297 = uncoded_block[1615] ^ uncoded_block[1618];
  wire _7298 = uncoded_block[1619] ^ uncoded_block[1621];
  wire _7299 = _7297 ^ _7298;
  wire _7300 = uncoded_block[1622] ^ uncoded_block[1623];
  wire _7301 = _7300 ^ _5386;
  wire _7302 = _7299 ^ _7301;
  wire _7303 = _7296 ^ _7302;
  wire _7304 = _7291 ^ _7303;
  wire _7305 = uncoded_block[1631] ^ uncoded_block[1634];
  wire _7306 = uncoded_block[1635] ^ uncoded_block[1636];
  wire _7307 = _7305 ^ _7306;
  wire _7308 = uncoded_block[1638] ^ uncoded_block[1639];
  wire _7309 = uncoded_block[1640] ^ uncoded_block[1642];
  wire _7310 = _7308 ^ _7309;
  wire _7311 = _7307 ^ _7310;
  wire _7312 = uncoded_block[1645] ^ uncoded_block[1647];
  wire _7313 = _7312 ^ _1649;
  wire _7314 = uncoded_block[1650] ^ uncoded_block[1656];
  wire _7315 = _7314 ^ _1653;
  wire _7316 = _7313 ^ _7315;
  wire _7317 = _7311 ^ _7316;
  wire _7318 = _823 ^ _1654;
  wire _7319 = uncoded_block[1665] ^ uncoded_block[1666];
  wire _7320 = _7319 ^ _4687;
  wire _7321 = _7318 ^ _7320;
  wire _7322 = uncoded_block[1669] ^ uncoded_block[1672];
  wire _7323 = uncoded_block[1673] ^ uncoded_block[1674];
  wire _7324 = _7322 ^ _7323;
  wire _7325 = uncoded_block[1677] ^ uncoded_block[1679];
  wire _7326 = _7325 ^ _6061;
  wire _7327 = _7324 ^ _7326;
  wire _7328 = _7321 ^ _7327;
  wire _7329 = _7317 ^ _7328;
  wire _7330 = _7304 ^ _7329;
  wire _7331 = uncoded_block[1690] ^ uncoded_block[1691];
  wire _7332 = _3189 ^ _7331;
  wire _7333 = _3968 ^ _5409;
  wire _7334 = _7332 ^ _7333;
  wire _7335 = uncoded_block[1707] ^ uncoded_block[1710];
  wire _7336 = _3973 ^ _7335;
  wire _7337 = uncoded_block[1711] ^ uncoded_block[1712];
  wire _7338 = _7337 ^ _854;
  wire _7339 = _7336 ^ _7338;
  wire _7340 = _7334 ^ _7339;
  wire _7341 = uncoded_block[1716] ^ uncoded_block[1720];
  wire _7342 = _7341 ^ uncoded_block[1721];
  wire _7343 = _7340 ^ _7342;
  wire _7344 = _7330 ^ _7343;
  wire _7345 = _7284 ^ _7344;
  wire _7346 = _7106 ^ _7345;
  wire _7347 = uncoded_block[2] ^ uncoded_block[5];
  wire _7348 = _7347 ^ _3993;
  wire _7349 = _3995 ^ _6083;
  wire _7350 = _7348 ^ _7349;
  wire _7351 = uncoded_block[16] ^ uncoded_block[19];
  wire _7352 = _6086 ^ _7351;
  wire _7353 = uncoded_block[22] ^ uncoded_block[24];
  wire _7354 = _7353 ^ _3224;
  wire _7355 = _7352 ^ _7354;
  wire _7356 = _7350 ^ _7355;
  wire _7357 = _875 ^ _879;
  wire _7358 = _7357 ^ _2467;
  wire _7359 = uncoded_block[46] ^ uncoded_block[48];
  wire _7360 = _22 ^ _7359;
  wire _7361 = _7360 ^ _5437;
  wire _7362 = _7358 ^ _7361;
  wire _7363 = _7356 ^ _7362;
  wire _7364 = uncoded_block[59] ^ uncoded_block[60];
  wire _7365 = uncoded_block[61] ^ uncoded_block[63];
  wire _7366 = _7364 ^ _7365;
  wire _7367 = uncoded_block[69] ^ uncoded_block[70];
  wire _7368 = _1706 ^ _7367;
  wire _7369 = _7366 ^ _7368;
  wire _7370 = _5442 ^ _1714;
  wire _7371 = _4735 ^ _6755;
  wire _7372 = _7370 ^ _7371;
  wire _7373 = _7369 ^ _7372;
  wire _7374 = uncoded_block[91] ^ uncoded_block[95];
  wire _7375 = uncoded_block[96] ^ uncoded_block[99];
  wire _7376 = _7374 ^ _7375;
  wire _7377 = uncoded_block[100] ^ uncoded_block[102];
  wire _7378 = _7377 ^ _4031;
  wire _7379 = _7376 ^ _7378;
  wire _7380 = _6123 ^ _914;
  wire _7381 = _915 ^ _1729;
  wire _7382 = _7380 ^ _7381;
  wire _7383 = _7379 ^ _7382;
  wire _7384 = _7373 ^ _7383;
  wire _7385 = _7363 ^ _7384;
  wire _7386 = uncoded_block[124] ^ uncoded_block[126];
  wire _7387 = _3255 ^ _7386;
  wire _7388 = uncoded_block[130] ^ uncoded_block[133];
  wire _7389 = _57 ^ _7388;
  wire _7390 = _7387 ^ _7389;
  wire _7391 = uncoded_block[137] ^ uncoded_block[143];
  wire _7392 = uncoded_block[144] ^ uncoded_block[145];
  wire _7393 = _7391 ^ _7392;
  wire _7394 = _67 ^ _70;
  wire _7395 = _7393 ^ _7394;
  wire _7396 = _7390 ^ _7395;
  wire _7397 = uncoded_block[154] ^ uncoded_block[155];
  wire _7398 = _7397 ^ _1748;
  wire _7399 = uncoded_block[168] ^ uncoded_block[170];
  wire _7400 = _933 ^ _7399;
  wire _7401 = _7398 ^ _7400;
  wire _7402 = _938 ^ _3278;
  wire _7403 = uncoded_block[178] ^ uncoded_block[180];
  wire _7404 = _82 ^ _7403;
  wire _7405 = _7402 ^ _7404;
  wire _7406 = _7401 ^ _7405;
  wire _7407 = _7396 ^ _7406;
  wire _7408 = uncoded_block[183] ^ uncoded_block[186];
  wire _7409 = uncoded_block[188] ^ uncoded_block[190];
  wire _7410 = _7408 ^ _7409;
  wire _7411 = uncoded_block[194] ^ uncoded_block[196];
  wire _7412 = _6798 ^ _7411;
  wire _7413 = _7410 ^ _7412;
  wire _7414 = _95 ^ _4070;
  wire _7415 = uncoded_block[209] ^ uncoded_block[211];
  wire _7416 = _4780 ^ _7415;
  wire _7417 = _7414 ^ _7416;
  wire _7418 = _7413 ^ _7417;
  wire _7419 = uncoded_block[222] ^ uncoded_block[224];
  wire _7420 = _5491 ^ _7419;
  wire _7421 = _7420 ^ _4082;
  wire _7422 = uncoded_block[232] ^ uncoded_block[234];
  wire _7423 = uncoded_block[236] ^ uncoded_block[237];
  wire _7424 = _7422 ^ _7423;
  wire _7425 = uncoded_block[238] ^ uncoded_block[241];
  wire _7426 = _7425 ^ _113;
  wire _7427 = _7424 ^ _7426;
  wire _7428 = _7421 ^ _7427;
  wire _7429 = _7418 ^ _7428;
  wire _7430 = _7407 ^ _7429;
  wire _7431 = _7385 ^ _7430;
  wire _7432 = uncoded_block[248] ^ uncoded_block[249];
  wire _7433 = _6180 ^ _7432;
  wire _7434 = uncoded_block[250] ^ uncoded_block[252];
  wire _7435 = uncoded_block[253] ^ uncoded_block[257];
  wire _7436 = _7434 ^ _7435;
  wire _7437 = _7433 ^ _7436;
  wire _7438 = uncoded_block[260] ^ uncoded_block[261];
  wire _7439 = _7438 ^ _977;
  wire _7440 = uncoded_block[267] ^ uncoded_block[268];
  wire _7441 = uncoded_block[269] ^ uncoded_block[272];
  wire _7442 = _7440 ^ _7441;
  wire _7443 = _7439 ^ _7442;
  wire _7444 = _7437 ^ _7443;
  wire _7445 = uncoded_block[278] ^ uncoded_block[279];
  wire _7446 = uncoded_block[282] ^ uncoded_block[284];
  wire _7447 = _7445 ^ _7446;
  wire _7448 = uncoded_block[285] ^ uncoded_block[289];
  wire _7449 = uncoded_block[292] ^ uncoded_block[296];
  wire _7450 = _7448 ^ _7449;
  wire _7451 = _7447 ^ _7450;
  wire _7452 = uncoded_block[297] ^ uncoded_block[301];
  wire _7453 = uncoded_block[302] ^ uncoded_block[305];
  wire _7454 = _7452 ^ _7453;
  wire _7455 = _3334 ^ _3337;
  wire _7456 = _7454 ^ _7455;
  wire _7457 = _7451 ^ _7456;
  wire _7458 = _7444 ^ _7457;
  wire _7459 = uncoded_block[311] ^ uncoded_block[317];
  wire _7460 = _7459 ^ _1008;
  wire _7461 = _4123 ^ _4125;
  wire _7462 = _7460 ^ _7461;
  wire _7463 = uncoded_block[337] ^ uncoded_block[338];
  wire _7464 = _3352 ^ _7463;
  wire _7465 = uncoded_block[345] ^ uncoded_block[347];
  wire _7466 = _7465 ^ _1028;
  wire _7467 = _7464 ^ _7466;
  wire _7468 = _7462 ^ _7467;
  wire _7469 = _3361 ^ _6864;
  wire _7470 = uncoded_block[365] ^ uncoded_block[366];
  wire _7471 = _1031 ^ _7470;
  wire _7472 = _7469 ^ _7471;
  wire _7473 = uncoded_block[368] ^ uncoded_block[375];
  wire _7474 = uncoded_block[376] ^ uncoded_block[378];
  wire _7475 = _7473 ^ _7474;
  wire _7476 = uncoded_block[379] ^ uncoded_block[380];
  wire _7477 = _7476 ^ _1038;
  wire _7478 = _7475 ^ _7477;
  wire _7479 = _7472 ^ _7478;
  wire _7480 = _7468 ^ _7479;
  wire _7481 = _7458 ^ _7480;
  wire _7482 = _3377 ^ _4149;
  wire _7483 = uncoded_block[388] ^ uncoded_block[391];
  wire _7484 = _7483 ^ _3383;
  wire _7485 = _7482 ^ _7484;
  wire _7486 = _6881 ^ _1849;
  wire _7487 = uncoded_block[403] ^ uncoded_block[404];
  wire _7488 = _181 ^ _7487;
  wire _7489 = _7486 ^ _7488;
  wire _7490 = _7485 ^ _7489;
  wire _7491 = _3391 ^ _3394;
  wire _7492 = uncoded_block[416] ^ uncoded_block[421];
  wire _7493 = _7492 ^ _2633;
  wire _7494 = _7491 ^ _7493;
  wire _7495 = uncoded_block[430] ^ uncoded_block[431];
  wire _7496 = _6894 ^ _7495;
  wire _7497 = uncoded_block[435] ^ uncoded_block[438];
  wire _7498 = uncoded_block[445] ^ uncoded_block[447];
  wire _7499 = _7497 ^ _7498;
  wire _7500 = _7496 ^ _7499;
  wire _7501 = _7494 ^ _7500;
  wire _7502 = _7490 ^ _7501;
  wire _7503 = _6900 ^ _212;
  wire _7504 = uncoded_block[457] ^ uncoded_block[459];
  wire _7505 = _7504 ^ _5586;
  wire _7506 = _7503 ^ _7505;
  wire _7507 = uncoded_block[464] ^ uncoded_block[466];
  wire _7508 = _7507 ^ _3418;
  wire _7509 = uncoded_block[472] ^ uncoded_block[474];
  wire _7510 = _7509 ^ _2657;
  wire _7511 = _7508 ^ _7510;
  wire _7512 = _7506 ^ _7511;
  wire _7513 = uncoded_block[478] ^ uncoded_block[480];
  wire _7514 = _7513 ^ _3423;
  wire _7515 = uncoded_block[486] ^ uncoded_block[487];
  wire _7516 = uncoded_block[488] ^ uncoded_block[489];
  wire _7517 = _7515 ^ _7516;
  wire _7518 = _7514 ^ _7517;
  wire _7519 = _2664 ^ _3432;
  wire _7520 = uncoded_block[495] ^ uncoded_block[499];
  wire _7521 = uncoded_block[501] ^ uncoded_block[503];
  wire _7522 = _7520 ^ _7521;
  wire _7523 = _7519 ^ _7522;
  wire _7524 = _7518 ^ _7523;
  wire _7525 = _7512 ^ _7524;
  wire _7526 = _7502 ^ _7525;
  wire _7527 = _7481 ^ _7526;
  wire _7528 = _7431 ^ _7527;
  wire _7529 = uncoded_block[506] ^ uncoded_block[508];
  wire _7530 = _2671 ^ _7529;
  wire _7531 = uncoded_block[509] ^ uncoded_block[511];
  wire _7532 = _7531 ^ _3439;
  wire _7533 = _7530 ^ _7532;
  wire _7534 = uncoded_block[526] ^ uncoded_block[529];
  wire _7535 = _1895 ^ _7534;
  wire _7536 = uncoded_block[538] ^ uncoded_block[539];
  wire _7537 = _4926 ^ _7536;
  wire _7538 = _7535 ^ _7537;
  wire _7539 = _7533 ^ _7538;
  wire _7540 = uncoded_block[540] ^ uncoded_block[542];
  wire _7541 = uncoded_block[543] ^ uncoded_block[546];
  wire _7542 = _7540 ^ _7541;
  wire _7543 = _1912 ^ _2688;
  wire _7544 = _7542 ^ _7543;
  wire _7545 = uncoded_block[562] ^ uncoded_block[565];
  wire _7546 = _3461 ^ _7545;
  wire _7547 = _1917 ^ _7546;
  wire _7548 = _7544 ^ _7547;
  wire _7549 = _7539 ^ _7548;
  wire _7550 = uncoded_block[567] ^ uncoded_block[568];
  wire _7551 = uncoded_block[570] ^ uncoded_block[573];
  wire _7552 = _7550 ^ _7551;
  wire _7553 = _6312 ^ _266;
  wire _7554 = _7552 ^ _7553;
  wire _7555 = uncoded_block[586] ^ uncoded_block[591];
  wire _7556 = uncoded_block[593] ^ uncoded_block[597];
  wire _7557 = _7555 ^ _7556;
  wire _7558 = uncoded_block[600] ^ uncoded_block[602];
  wire _7559 = _7558 ^ _3489;
  wire _7560 = _7557 ^ _7559;
  wire _7561 = _7554 ^ _7560;
  wire _7562 = _1146 ^ _278;
  wire _7563 = uncoded_block[612] ^ uncoded_block[613];
  wire _7564 = uncoded_block[614] ^ uncoded_block[615];
  wire _7565 = _7563 ^ _7564;
  wire _7566 = _7562 ^ _7565;
  wire _7567 = uncoded_block[616] ^ uncoded_block[618];
  wire _7568 = uncoded_block[620] ^ uncoded_block[622];
  wire _7569 = _7567 ^ _7568;
  wire _7570 = uncoded_block[624] ^ uncoded_block[626];
  wire _7571 = _7570 ^ _5658;
  wire _7572 = _7569 ^ _7571;
  wire _7573 = _7566 ^ _7572;
  wire _7574 = _7561 ^ _7573;
  wire _7575 = _7549 ^ _7574;
  wire _7576 = uncoded_block[630] ^ uncoded_block[633];
  wire _7577 = uncoded_block[634] ^ uncoded_block[636];
  wire _7578 = _7576 ^ _7577;
  wire _7579 = _5665 ^ _2727;
  wire _7580 = _7578 ^ _7579;
  wire _7581 = _6973 ^ _2738;
  wire _7582 = uncoded_block[663] ^ uncoded_block[665];
  wire _7583 = _2739 ^ _7582;
  wire _7584 = _7581 ^ _7583;
  wire _7585 = _7580 ^ _7584;
  wire _7586 = uncoded_block[668] ^ uncoded_block[671];
  wire _7587 = _309 ^ _7586;
  wire _7588 = _2748 ^ _319;
  wire _7589 = _7587 ^ _7588;
  wire _7590 = _1972 ^ _1974;
  wire _7591 = _326 ^ _328;
  wire _7592 = _7590 ^ _7591;
  wire _7593 = _7589 ^ _7592;
  wire _7594 = _7585 ^ _7593;
  wire _7595 = uncoded_block[703] ^ uncoded_block[707];
  wire _7596 = _3532 ^ _7595;
  wire _7597 = uncoded_block[709] ^ uncoded_block[712];
  wire _7598 = _7597 ^ _1983;
  wire _7599 = _7596 ^ _7598;
  wire _7600 = _5690 ^ _343;
  wire _7601 = _7600 ^ _3545;
  wire _7602 = _7599 ^ _7601;
  wire _7603 = uncoded_block[729] ^ uncoded_block[731];
  wire _7604 = _7603 ^ _3547;
  wire _7605 = uncoded_block[735] ^ uncoded_block[737];
  wire _7606 = _7605 ^ _352;
  wire _7607 = _7604 ^ _7606;
  wire _7608 = _1210 ^ _7015;
  wire _7609 = _5703 ^ _7608;
  wire _7610 = _7607 ^ _7609;
  wire _7611 = _7602 ^ _7610;
  wire _7612 = _7594 ^ _7611;
  wire _7613 = _7575 ^ _7612;
  wire _7614 = uncoded_block[758] ^ uncoded_block[762];
  wire _7615 = _7614 ^ _1217;
  wire _7616 = uncoded_block[765] ^ uncoded_block[768];
  wire _7617 = uncoded_block[769] ^ uncoded_block[771];
  wire _7618 = _7616 ^ _7617;
  wire _7619 = _7615 ^ _7618;
  wire _7620 = uncoded_block[773] ^ uncoded_block[776];
  wire _7621 = _7620 ^ _368;
  wire _7622 = uncoded_block[786] ^ uncoded_block[789];
  wire _7623 = _3568 ^ _7622;
  wire _7624 = _7621 ^ _7623;
  wire _7625 = _7619 ^ _7624;
  wire _7626 = uncoded_block[790] ^ uncoded_block[792];
  wire _7627 = _7626 ^ _5723;
  wire _7628 = uncoded_block[797] ^ uncoded_block[799];
  wire _7629 = uncoded_block[801] ^ uncoded_block[804];
  wire _7630 = _7628 ^ _7629;
  wire _7631 = _7627 ^ _7630;
  wire _7632 = uncoded_block[811] ^ uncoded_block[815];
  wire _7633 = _1238 ^ _7632;
  wire _7634 = uncoded_block[818] ^ uncoded_block[820];
  wire _7635 = _7634 ^ _3587;
  wire _7636 = _7633 ^ _7635;
  wire _7637 = _7631 ^ _7636;
  wire _7638 = _7625 ^ _7637;
  wire _7639 = _1249 ^ _4336;
  wire _7640 = uncoded_block[841] ^ uncoded_block[843];
  wire _7641 = _4337 ^ _7640;
  wire _7642 = _7639 ^ _7641;
  wire _7643 = uncoded_block[849] ^ uncoded_block[850];
  wire _7644 = uncoded_block[851] ^ uncoded_block[854];
  wire _7645 = _7643 ^ _7644;
  wire _7646 = _5061 ^ _7645;
  wire _7647 = _7642 ^ _7646;
  wire _7648 = _3600 ^ _5066;
  wire _7649 = uncoded_block[860] ^ uncoded_block[863];
  wire _7650 = uncoded_block[864] ^ uncoded_block[866];
  wire _7651 = _7649 ^ _7650;
  wire _7652 = _7648 ^ _7651;
  wire _7653 = _5072 ^ _416;
  wire _7654 = uncoded_block[875] ^ uncoded_block[880];
  wire _7655 = _7654 ^ _2836;
  wire _7656 = _7653 ^ _7655;
  wire _7657 = _7652 ^ _7656;
  wire _7658 = _7647 ^ _7657;
  wire _7659 = _7638 ^ _7658;
  wire _7660 = uncoded_block[887] ^ uncoded_block[888];
  wire _7661 = _7660 ^ _3614;
  wire _7662 = _7661 ^ _5086;
  wire _7663 = uncoded_block[902] ^ uncoded_block[908];
  wire _7664 = _7663 ^ _6428;
  wire _7665 = uncoded_block[912] ^ uncoded_block[913];
  wire _7666 = _7665 ^ _3629;
  wire _7667 = _7664 ^ _7666;
  wire _7668 = _7662 ^ _7667;
  wire _7669 = _5766 ^ _4370;
  wire _7670 = uncoded_block[929] ^ uncoded_block[933];
  wire _7671 = _7670 ^ _5101;
  wire _7672 = _7669 ^ _7671;
  wire _7673 = uncoded_block[938] ^ uncoded_block[940];
  wire _7674 = _7673 ^ _6439;
  wire _7675 = uncoded_block[945] ^ uncoded_block[950];
  wire _7676 = _7675 ^ _7083;
  wire _7677 = _7674 ^ _7676;
  wire _7678 = _7672 ^ _7677;
  wire _7679 = _7668 ^ _7678;
  wire _7680 = uncoded_block[958] ^ uncoded_block[959];
  wire _7681 = _7680 ^ _5783;
  wire _7682 = uncoded_block[965] ^ uncoded_block[968];
  wire _7683 = _7682 ^ _7088;
  wire _7684 = _7681 ^ _7683;
  wire _7685 = _468 ^ _470;
  wire _7686 = _471 ^ _476;
  wire _7687 = _7685 ^ _7686;
  wire _7688 = _7684 ^ _7687;
  wire _7689 = uncoded_block[983] ^ uncoded_block[985];
  wire _7690 = _7689 ^ _1317;
  wire _7691 = uncoded_block[1000] ^ uncoded_block[1001];
  wire _7692 = _6453 ^ _7691;
  wire _7693 = _7690 ^ _7692;
  wire _7694 = _4404 ^ _2886;
  wire _7695 = _487 ^ _491;
  wire _7696 = _7694 ^ _7695;
  wire _7697 = _7693 ^ _7696;
  wire _7698 = _7688 ^ _7697;
  wire _7699 = _7679 ^ _7698;
  wire _7700 = _7659 ^ _7699;
  wire _7701 = _7613 ^ _7700;
  wire _7702 = _7528 ^ _7701;
  wire _7703 = uncoded_block[1015] ^ uncoded_block[1017];
  wire _7704 = _7703 ^ _1338;
  wire _7705 = _495 ^ _498;
  wire _7706 = _7704 ^ _7705;
  wire _7707 = uncoded_block[1034] ^ uncoded_block[1036];
  wire _7708 = _4417 ^ _7707;
  wire _7709 = _2129 ^ _1346;
  wire _7710 = _7708 ^ _7709;
  wire _7711 = _7706 ^ _7710;
  wire _7712 = uncoded_block[1046] ^ uncoded_block[1049];
  wire _7713 = _514 ^ _7712;
  wire _7714 = uncoded_block[1050] ^ uncoded_block[1053];
  wire _7715 = _7714 ^ _4430;
  wire _7716 = _7713 ^ _7715;
  wire _7717 = uncoded_block[1060] ^ uncoded_block[1064];
  wire _7718 = _7117 ^ _7717;
  wire _7719 = _7718 ^ _3690;
  wire _7720 = _7716 ^ _7719;
  wire _7721 = _7711 ^ _7720;
  wire _7722 = uncoded_block[1072] ^ uncoded_block[1074];
  wire _7723 = _7722 ^ _3695;
  wire _7724 = uncoded_block[1081] ^ uncoded_block[1082];
  wire _7725 = uncoded_block[1084] ^ uncoded_block[1088];
  wire _7726 = _7724 ^ _7725;
  wire _7727 = _7723 ^ _7726;
  wire _7728 = _5843 ^ _5846;
  wire _7729 = _4443 ^ _7728;
  wire _7730 = _7727 ^ _7729;
  wire _7731 = uncoded_block[1101] ^ uncoded_block[1103];
  wire _7732 = _7731 ^ _3707;
  wire _7733 = _549 ^ _7132;
  wire _7734 = _7732 ^ _7733;
  wire _7735 = _7133 ^ _3713;
  wire _7736 = uncoded_block[1120] ^ uncoded_block[1121];
  wire _7737 = uncoded_block[1125] ^ uncoded_block[1136];
  wire _7738 = _7736 ^ _7737;
  wire _7739 = _7735 ^ _7738;
  wire _7740 = _7734 ^ _7739;
  wire _7741 = _7730 ^ _7740;
  wire _7742 = _7721 ^ _7741;
  wire _7743 = uncoded_block[1142] ^ uncoded_block[1146];
  wire _7744 = _3721 ^ _7743;
  wire _7745 = _6505 ^ _4468;
  wire _7746 = _7744 ^ _7745;
  wire _7747 = _3728 ^ _578;
  wire _7748 = uncoded_block[1160] ^ uncoded_block[1161];
  wire _7749 = uncoded_block[1162] ^ uncoded_block[1165];
  wire _7750 = _7748 ^ _7749;
  wire _7751 = _7747 ^ _7750;
  wire _7752 = _7746 ^ _7751;
  wire _7753 = _2967 ^ _4481;
  wire _7754 = _590 ^ _3746;
  wire _7755 = _7753 ^ _7754;
  wire _7756 = uncoded_block[1190] ^ uncoded_block[1193];
  wire _7757 = _7756 ^ _6525;
  wire _7758 = uncoded_block[1198] ^ uncoded_block[1200];
  wire _7759 = _1421 ^ _7758;
  wire _7760 = _7757 ^ _7759;
  wire _7761 = _7755 ^ _7760;
  wire _7762 = _7752 ^ _7761;
  wire _7763 = uncoded_block[1201] ^ uncoded_block[1203];
  wire _7764 = _7763 ^ _4491;
  wire _7765 = uncoded_block[1209] ^ uncoded_block[1211];
  wire _7766 = uncoded_block[1212] ^ uncoded_block[1217];
  wire _7767 = _7765 ^ _7766;
  wire _7768 = _7764 ^ _7767;
  wire _7769 = _606 ^ _1433;
  wire _7770 = _612 ^ _1439;
  wire _7771 = _7769 ^ _7770;
  wire _7772 = _7768 ^ _7771;
  wire _7773 = uncoded_block[1231] ^ uncoded_block[1235];
  wire _7774 = uncoded_block[1236] ^ uncoded_block[1240];
  wire _7775 = _7773 ^ _7774;
  wire _7776 = _1448 ^ _2232;
  wire _7777 = _7775 ^ _7776;
  wire _7778 = uncoded_block[1251] ^ uncoded_block[1252];
  wire _7779 = _7778 ^ _3780;
  wire _7780 = uncoded_block[1257] ^ uncoded_block[1258];
  wire _7781 = uncoded_block[1259] ^ uncoded_block[1260];
  wire _7782 = _7780 ^ _7781;
  wire _7783 = _7779 ^ _7782;
  wire _7784 = _7777 ^ _7783;
  wire _7785 = _7772 ^ _7784;
  wire _7786 = _7762 ^ _7785;
  wire _7787 = _7742 ^ _7786;
  wire _7788 = uncoded_block[1267] ^ uncoded_block[1270];
  wire _7789 = _7788 ^ _628;
  wire _7790 = _3005 ^ _7789;
  wire _7791 = uncoded_block[1273] ^ uncoded_block[1275];
  wire _7792 = uncoded_block[1276] ^ uncoded_block[1277];
  wire _7793 = _7791 ^ _7792;
  wire _7794 = _631 ^ _4525;
  wire _7795 = _7793 ^ _7794;
  wire _7796 = _7790 ^ _7795;
  wire _7797 = uncoded_block[1286] ^ uncoded_block[1291];
  wire _7798 = _638 ^ _7797;
  wire _7799 = uncoded_block[1297] ^ uncoded_block[1299];
  wire _7800 = _3801 ^ _7799;
  wire _7801 = _7798 ^ _7800;
  wire _7802 = uncoded_block[1307] ^ uncoded_block[1310];
  wire _7803 = _648 ^ _7802;
  wire _7804 = uncoded_block[1311] ^ uncoded_block[1315];
  wire _7805 = uncoded_block[1318] ^ uncoded_block[1321];
  wire _7806 = _7804 ^ _7805;
  wire _7807 = _7803 ^ _7806;
  wire _7808 = _7801 ^ _7807;
  wire _7809 = _7796 ^ _7808;
  wire _7810 = _4543 ^ _1489;
  wire _7811 = uncoded_block[1328] ^ uncoded_block[1334];
  wire _7812 = _7811 ^ _3034;
  wire _7813 = _7810 ^ _7812;
  wire _7814 = uncoded_block[1338] ^ uncoded_block[1341];
  wire _7815 = uncoded_block[1342] ^ uncoded_block[1343];
  wire _7816 = _7814 ^ _7815;
  wire _7817 = uncoded_block[1352] ^ uncoded_block[1358];
  wire _7818 = _1498 ^ _7817;
  wire _7819 = _7816 ^ _7818;
  wire _7820 = _7813 ^ _7819;
  wire _7821 = uncoded_block[1359] ^ uncoded_block[1361];
  wire _7822 = _7821 ^ _3828;
  wire _7823 = uncoded_block[1372] ^ uncoded_block[1375];
  wire _7824 = uncoded_block[1376] ^ uncoded_block[1378];
  wire _7825 = _7823 ^ _7824;
  wire _7826 = _7822 ^ _7825;
  wire _7827 = _7219 ^ _3059;
  wire _7828 = uncoded_block[1391] ^ uncoded_block[1393];
  wire _7829 = _691 ^ _7828;
  wire _7830 = _7827 ^ _7829;
  wire _7831 = _7826 ^ _7830;
  wire _7832 = _7820 ^ _7831;
  wire _7833 = _7809 ^ _7832;
  wire _7834 = uncoded_block[1395] ^ uncoded_block[1398];
  wire _7835 = _7834 ^ _3841;
  wire _7836 = _3846 ^ _2300;
  wire _7837 = _7835 ^ _7836;
  wire _7838 = _3849 ^ _702;
  wire _7839 = _704 ^ _3850;
  wire _7840 = _7838 ^ _7839;
  wire _7841 = _7837 ^ _7840;
  wire _7842 = uncoded_block[1421] ^ uncoded_block[1422];
  wire _7843 = _7842 ^ _1527;
  wire _7844 = uncoded_block[1426] ^ uncoded_block[1427];
  wire _7845 = _7844 ^ _5968;
  wire _7846 = _7843 ^ _7845;
  wire _7847 = _2313 ^ _3083;
  wire _7848 = _3862 ^ _3864;
  wire _7849 = _7847 ^ _7848;
  wire _7850 = _7846 ^ _7849;
  wire _7851 = _7841 ^ _7850;
  wire _7852 = uncoded_block[1451] ^ uncoded_block[1455];
  wire _7853 = _3865 ^ _7852;
  wire _7854 = _3088 ^ _7241;
  wire _7855 = _7853 ^ _7854;
  wire _7856 = _3871 ^ _1548;
  wire _7857 = _1551 ^ _1555;
  wire _7858 = _7856 ^ _7857;
  wire _7859 = _7855 ^ _7858;
  wire _7860 = _3884 ^ _1559;
  wire _7861 = uncoded_block[1484] ^ uncoded_block[1486];
  wire _7862 = _7861 ^ _7251;
  wire _7863 = _7860 ^ _7862;
  wire _7864 = uncoded_block[1496] ^ uncoded_block[1498];
  wire _7865 = _7864 ^ _747;
  wire _7866 = uncoded_block[1501] ^ uncoded_block[1502];
  wire _7867 = _7866 ^ _1572;
  wire _7868 = _7865 ^ _7867;
  wire _7869 = _7863 ^ _7868;
  wire _7870 = _7859 ^ _7869;
  wire _7871 = _7851 ^ _7870;
  wire _7872 = _7833 ^ _7871;
  wire _7873 = _7787 ^ _7872;
  wire _7874 = uncoded_block[1505] ^ uncoded_block[1508];
  wire _7875 = uncoded_block[1511] ^ uncoded_block[1512];
  wire _7876 = _7874 ^ _7875;
  wire _7877 = _3115 ^ _6643;
  wire _7878 = _7876 ^ _7877;
  wire _7879 = _2357 ^ _3900;
  wire _7880 = _5343 ^ _757;
  wire _7881 = _7879 ^ _7880;
  wire _7882 = _7878 ^ _7881;
  wire _7883 = uncoded_block[1541] ^ uncoded_block[1544];
  wire _7884 = _6651 ^ _7883;
  wire _7885 = uncoded_block[1552] ^ uncoded_block[1554];
  wire _7886 = _2367 ^ _7885;
  wire _7887 = _7884 ^ _7886;
  wire _7888 = uncoded_block[1559] ^ uncoded_block[1561];
  wire _7889 = uncoded_block[1562] ^ uncoded_block[1564];
  wire _7890 = _7888 ^ _7889;
  wire _7891 = uncoded_block[1568] ^ uncoded_block[1570];
  wire _7892 = uncoded_block[1571] ^ uncoded_block[1575];
  wire _7893 = _7891 ^ _7892;
  wire _7894 = _7890 ^ _7893;
  wire _7895 = _7887 ^ _7894;
  wire _7896 = _7882 ^ _7895;
  wire _7897 = uncoded_block[1581] ^ uncoded_block[1584];
  wire _7898 = _6029 ^ _7897;
  wire _7899 = _2386 ^ _5368;
  wire _7900 = _7898 ^ _7899;
  wire _7901 = _3146 ^ _792;
  wire _7902 = uncoded_block[1602] ^ uncoded_block[1606];
  wire _7903 = _3934 ^ _7902;
  wire _7904 = _7901 ^ _7903;
  wire _7905 = _7900 ^ _7904;
  wire _7906 = uncoded_block[1609] ^ uncoded_block[1611];
  wire _7907 = _2396 ^ _7906;
  wire _7908 = uncoded_block[1612] ^ uncoded_block[1613];
  wire _7909 = _7908 ^ _7297;
  wire _7910 = _7907 ^ _7909;
  wire _7911 = uncoded_block[1619] ^ uncoded_block[1620];
  wire _7912 = uncoded_block[1621] ^ uncoded_block[1622];
  wire _7913 = _7911 ^ _7912;
  wire _7914 = uncoded_block[1633] ^ uncoded_block[1634];
  wire _7915 = _3942 ^ _7914;
  wire _7916 = _7913 ^ _7915;
  wire _7917 = _7910 ^ _7916;
  wire _7918 = _7905 ^ _7917;
  wire _7919 = _7896 ^ _7918;
  wire _7920 = _1642 ^ _7309;
  wire _7921 = uncoded_block[1643] ^ uncoded_block[1647];
  wire _7922 = uncoded_block[1648] ^ uncoded_block[1654];
  wire _7923 = _7921 ^ _7922;
  wire _7924 = _7920 ^ _7923;
  wire _7925 = uncoded_block[1655] ^ uncoded_block[1657];
  wire _7926 = _7925 ^ _1653;
  wire _7927 = uncoded_block[1661] ^ uncoded_block[1664];
  wire _7928 = uncoded_block[1669] ^ uncoded_block[1670];
  wire _7929 = _7927 ^ _7928;
  wire _7930 = _7926 ^ _7929;
  wire _7931 = _7924 ^ _7930;
  wire _7932 = uncoded_block[1671] ^ uncoded_block[1679];
  wire _7933 = uncoded_block[1681] ^ uncoded_block[1685];
  wire _7934 = _7932 ^ _7933;
  wire _7935 = uncoded_block[1689] ^ uncoded_block[1691];
  wire _7936 = _1665 ^ _7935;
  wire _7937 = _7934 ^ _7936;
  wire _7938 = _3968 ^ _4700;
  wire _7939 = _3976 ^ _2435;
  wire _7940 = _7938 ^ _7939;
  wire _7941 = _7937 ^ _7940;
  wire _7942 = _7931 ^ _7941;
  wire _7943 = uncoded_block[1708] ^ uncoded_block[1713];
  wire _7944 = uncoded_block[1714] ^ uncoded_block[1716];
  wire _7945 = _7943 ^ _7944;
  wire _7946 = uncoded_block[1717] ^ uncoded_block[1720];
  wire _7947 = _7946 ^ uncoded_block[1722];
  wire _7948 = _7945 ^ _7947;
  wire _7949 = _7942 ^ _7948;
  wire _7950 = _7919 ^ _7949;
  wire _7951 = _7873 ^ _7950;
  wire _7952 = _7702 ^ _7951;
  wire _7953 = _3209 ^ _7347;
  wire _7954 = _1684 ^ _7;
  wire _7955 = _7953 ^ _7954;
  wire _7956 = uncoded_block[13] ^ uncoded_block[14];
  wire _7957 = uncoded_block[16] ^ uncoded_block[20];
  wire _7958 = _7956 ^ _7957;
  wire _7959 = uncoded_block[26] ^ uncoded_block[27];
  wire _7960 = _10 ^ _7959;
  wire _7961 = _7958 ^ _7960;
  wire _7962 = _7955 ^ _7961;
  wire _7963 = _879 ^ _18;
  wire _7964 = _876 ^ _7963;
  wire _7965 = uncoded_block[42] ^ uncoded_block[43];
  wire _7966 = uncoded_block[44] ^ uncoded_block[47];
  wire _7967 = _7965 ^ _7966;
  wire _7968 = uncoded_block[48] ^ uncoded_block[53];
  wire _7969 = uncoded_block[57] ^ uncoded_block[59];
  wire _7970 = _7968 ^ _7969;
  wire _7971 = _7967 ^ _7970;
  wire _7972 = _7964 ^ _7971;
  wire _7973 = _7962 ^ _7972;
  wire _7974 = uncoded_block[60] ^ uncoded_block[65];
  wire _7975 = _7974 ^ _6744;
  wire _7976 = uncoded_block[70] ^ uncoded_block[71];
  wire _7977 = _7976 ^ _897;
  wire _7978 = _7975 ^ _7977;
  wire _7979 = uncoded_block[77] ^ uncoded_block[80];
  wire _7980 = _4020 ^ _7979;
  wire _7981 = uncoded_block[88] ^ uncoded_block[91];
  wire _7982 = _4025 ^ _7981;
  wire _7983 = _7980 ^ _7982;
  wire _7984 = _7978 ^ _7983;
  wire _7985 = uncoded_block[92] ^ uncoded_block[98];
  wire _7986 = uncoded_block[103] ^ uncoded_block[104];
  wire _7987 = _7985 ^ _7986;
  wire _7988 = _911 ^ _4034;
  wire _7989 = _7987 ^ _7988;
  wire _7990 = uncoded_block[113] ^ uncoded_block[114];
  wire _7991 = _7990 ^ _56;
  wire _7992 = _7386 ^ _1733;
  wire _7993 = _7991 ^ _7992;
  wire _7994 = _7989 ^ _7993;
  wire _7995 = _7984 ^ _7994;
  wire _7996 = _7973 ^ _7995;
  wire _7997 = uncoded_block[134] ^ uncoded_block[138];
  wire _7998 = _2504 ^ _7997;
  wire _7999 = uncoded_block[139] ^ uncoded_block[142];
  wire _8000 = uncoded_block[148] ^ uncoded_block[151];
  wire _8001 = _7999 ^ _8000;
  wire _8002 = _7998 ^ _8001;
  wire _8003 = uncoded_block[152] ^ uncoded_block[155];
  wire _8004 = _8003 ^ _1748;
  wire _8005 = _78 ^ _4056;
  wire _8006 = _8004 ^ _8005;
  wire _8007 = _8002 ^ _8006;
  wire _8008 = _81 ^ _1756;
  wire _8009 = uncoded_block[180] ^ uncoded_block[181];
  wire _8010 = _940 ^ _8009;
  wire _8011 = _8008 ^ _8010;
  wire _8012 = _86 ^ _1759;
  wire _8013 = _945 ^ _5483;
  wire _8014 = _8012 ^ _8013;
  wire _8015 = _8011 ^ _8014;
  wire _8016 = _8007 ^ _8015;
  wire _8017 = _4776 ^ _2532;
  wire _8018 = uncoded_block[199] ^ uncoded_block[201];
  wire _8019 = _8018 ^ _3289;
  wire _8020 = _8017 ^ _8019;
  wire _8021 = uncoded_block[204] ^ uncoded_block[207];
  wire _8022 = _8021 ^ _955;
  wire _8023 = uncoded_block[215] ^ uncoded_block[220];
  wire _8024 = _3295 ^ _8023;
  wire _8025 = _8022 ^ _8024;
  wire _8026 = _8020 ^ _8025;
  wire _8027 = _4788 ^ _6168;
  wire _8028 = uncoded_block[228] ^ uncoded_block[231];
  wire _8029 = uncoded_block[232] ^ uncoded_block[235];
  wire _8030 = _8028 ^ _8029;
  wire _8031 = _8027 ^ _8030;
  wire _8032 = uncoded_block[241] ^ uncoded_block[246];
  wire _8033 = _7423 ^ _8032;
  wire _8034 = uncoded_block[250] ^ uncoded_block[253];
  wire _8035 = _8034 ^ _3311;
  wire _8036 = _8033 ^ _8035;
  wire _8037 = _8031 ^ _8036;
  wire _8038 = _8026 ^ _8037;
  wire _8039 = _8016 ^ _8038;
  wire _8040 = _7996 ^ _8039;
  wire _8041 = uncoded_block[257] ^ uncoded_block[259];
  wire _8042 = _8041 ^ _120;
  wire _8043 = _1792 ^ _130;
  wire _8044 = _8042 ^ _8043;
  wire _8045 = uncoded_block[276] ^ uncoded_block[283];
  wire _8046 = _8045 ^ _1803;
  wire _8047 = _992 ^ _3328;
  wire _8048 = _8046 ^ _8047;
  wire _8049 = _8044 ^ _8048;
  wire _8050 = _4820 ^ _1806;
  wire _8051 = uncoded_block[298] ^ uncoded_block[302];
  wire _8052 = uncoded_block[303] ^ uncoded_block[305];
  wire _8053 = _8051 ^ _8052;
  wire _8054 = _8050 ^ _8053;
  wire _8055 = uncoded_block[306] ^ uncoded_block[307];
  wire _8056 = uncoded_block[310] ^ uncoded_block[311];
  wire _8057 = _8055 ^ _8056;
  wire _8058 = uncoded_block[324] ^ uncoded_block[327];
  wire _8059 = _4830 ^ _8058;
  wire _8060 = _8057 ^ _8059;
  wire _8061 = _8054 ^ _8060;
  wire _8062 = _8049 ^ _8061;
  wire _8063 = uncoded_block[331] ^ uncoded_block[332];
  wire _8064 = _8063 ^ _5536;
  wire _8065 = uncoded_block[336] ^ uncoded_block[338];
  wire _8066 = _8065 ^ _2595;
  wire _8067 = _8064 ^ _8066;
  wire _8068 = _4844 ^ _2599;
  wire _8069 = uncoded_block[354] ^ uncoded_block[356];
  wire _8070 = _162 ^ _8069;
  wire _8071 = _8068 ^ _8070;
  wire _8072 = _8067 ^ _8071;
  wire _8073 = uncoded_block[357] ^ uncoded_block[360];
  wire _8074 = _8073 ^ _5548;
  wire _8075 = uncoded_block[365] ^ uncoded_block[368];
  wire _8076 = uncoded_block[369] ^ uncoded_block[370];
  wire _8077 = _8075 ^ _8076;
  wire _8078 = _8074 ^ _8077;
  wire _8079 = uncoded_block[375] ^ uncoded_block[376];
  wire _8080 = _6873 ^ _8079;
  wire _8081 = _2609 ^ _4149;
  wire _8082 = _8080 ^ _8081;
  wire _8083 = _8078 ^ _8082;
  wire _8084 = _8072 ^ _8083;
  wire _8085 = _8062 ^ _8084;
  wire _8086 = _3381 ^ _3384;
  wire _8087 = uncoded_block[398] ^ uncoded_block[401];
  wire _8088 = uncoded_block[403] ^ uncoded_block[407];
  wire _8089 = _8087 ^ _8088;
  wire _8090 = _8086 ^ _8089;
  wire _8091 = uncoded_block[410] ^ uncoded_block[411];
  wire _8092 = uncoded_block[414] ^ uncoded_block[417];
  wire _8093 = _8091 ^ _8092;
  wire _8094 = _4164 ^ _197;
  wire _8095 = _8093 ^ _8094;
  wire _8096 = _8090 ^ _8095;
  wire _8097 = _6894 ^ _1857;
  wire _8098 = uncoded_block[438] ^ uncoded_block[441];
  wire _8099 = _6255 ^ _8098;
  wire _8100 = _8097 ^ _8099;
  wire _8101 = _5578 ^ _6259;
  wire _8102 = _8101 ^ _6901;
  wire _8103 = _8100 ^ _8102;
  wire _8104 = _8096 ^ _8103;
  wire _8105 = uncoded_block[461] ^ uncoded_block[465];
  wire _8106 = _3415 ^ _8105;
  wire _8107 = _3416 ^ _1082;
  wire _8108 = _8106 ^ _8107;
  wire _8109 = _2657 ^ _3421;
  wire _8110 = uncoded_block[480] ^ uncoded_block[482];
  wire _8111 = uncoded_block[483] ^ uncoded_block[486];
  wire _8112 = _8110 ^ _8111;
  wire _8113 = _8109 ^ _8112;
  wire _8114 = _8108 ^ _8113;
  wire _8115 = uncoded_block[489] ^ uncoded_block[491];
  wire _8116 = _6276 ^ _8115;
  wire _8117 = uncoded_block[493] ^ uncoded_block[495];
  wire _8118 = _8117 ^ _228;
  wire _8119 = _8116 ^ _8118;
  wire _8120 = uncoded_block[501] ^ uncoded_block[504];
  wire _8121 = _8120 ^ _1892;
  wire _8122 = uncoded_block[512] ^ uncoded_block[515];
  wire _8123 = _7531 ^ _8122;
  wire _8124 = _8121 ^ _8123;
  wire _8125 = _8119 ^ _8124;
  wire _8126 = _8114 ^ _8125;
  wire _8127 = _8104 ^ _8126;
  wire _8128 = _8085 ^ _8127;
  wire _8129 = _8040 ^ _8128;
  wire _8130 = _4918 ^ _3445;
  wire _8131 = _8130 ^ _5618;
  wire _8132 = uncoded_block[541] ^ uncoded_block[542];
  wire _8133 = _8132 ^ _244;
  wire _8134 = uncoded_block[550] ^ uncoded_block[553];
  wire _8135 = _6300 ^ _8134;
  wire _8136 = _8133 ^ _8135;
  wire _8137 = _8131 ^ _8136;
  wire _8138 = _6304 ^ _1916;
  wire _8139 = uncoded_block[559] ^ uncoded_block[560];
  wire _8140 = _8139 ^ _5633;
  wire _8141 = _8138 ^ _8140;
  wire _8142 = _6942 ^ _6945;
  wire _8143 = uncoded_block[583] ^ uncoded_block[587];
  wire _8144 = _1138 ^ _8143;
  wire _8145 = _8142 ^ _8144;
  wire _8146 = _8141 ^ _8145;
  wire _8147 = _8137 ^ _8146;
  wire _8148 = uncoded_block[592] ^ uncoded_block[595];
  wire _8149 = uncoded_block[596] ^ uncoded_block[597];
  wire _8150 = _8148 ^ _8149;
  wire _8151 = _4951 ^ _8150;
  wire _8152 = uncoded_block[604] ^ uncoded_block[606];
  wire _8153 = _7558 ^ _8152;
  wire _8154 = uncoded_block[610] ^ uncoded_block[611];
  wire _8155 = uncoded_block[612] ^ uncoded_block[617];
  wire _8156 = _8154 ^ _8155;
  wire _8157 = _8153 ^ _8156;
  wire _8158 = _8151 ^ _8157;
  wire _8159 = uncoded_block[625] ^ uncoded_block[628];
  wire _8160 = _4243 ^ _8159;
  wire _8161 = uncoded_block[630] ^ uncoded_block[632];
  wire _8162 = _8161 ^ _6331;
  wire _8163 = _8160 ^ _8162;
  wire _8164 = _293 ^ _4972;
  wire _8165 = uncoded_block[647] ^ uncoded_block[650];
  wire _8166 = uncoded_block[651] ^ uncoded_block[654];
  wire _8167 = _8165 ^ _8166;
  wire _8168 = _8164 ^ _8167;
  wire _8169 = _8163 ^ _8168;
  wire _8170 = _8158 ^ _8169;
  wire _8171 = _8147 ^ _8170;
  wire _8172 = uncoded_block[659] ^ uncoded_block[661];
  wire _8173 = _2738 ^ _8172;
  wire _8174 = _4978 ^ _311;
  wire _8175 = _8173 ^ _8174;
  wire _8176 = uncoded_block[672] ^ uncoded_block[675];
  wire _8177 = uncoded_block[676] ^ uncoded_block[677];
  wire _8178 = _8176 ^ _8177;
  wire _8179 = uncoded_block[678] ^ uncoded_block[681];
  wire _8180 = uncoded_block[682] ^ uncoded_block[685];
  wire _8181 = _8179 ^ _8180;
  wire _8182 = _8178 ^ _8181;
  wire _8183 = _8175 ^ _8182;
  wire _8184 = uncoded_block[690] ^ uncoded_block[694];
  wire _8185 = _2751 ^ _8184;
  wire _8186 = uncoded_block[695] ^ uncoded_block[696];
  wire _8187 = _8186 ^ _6360;
  wire _8188 = _8185 ^ _8187;
  wire _8189 = uncoded_block[702] ^ uncoded_block[707];
  wire _8190 = uncoded_block[708] ^ uncoded_block[709];
  wire _8191 = _8189 ^ _8190;
  wire _8192 = uncoded_block[710] ^ uncoded_block[714];
  wire _8193 = uncoded_block[716] ^ uncoded_block[718];
  wire _8194 = _8192 ^ _8193;
  wire _8195 = _8191 ^ _8194;
  wire _8196 = _8188 ^ _8195;
  wire _8197 = _8183 ^ _8196;
  wire _8198 = uncoded_block[721] ^ uncoded_block[723];
  wire _8199 = _8198 ^ _1988;
  wire _8200 = uncoded_block[730] ^ uncoded_block[731];
  wire _8201 = uncoded_block[732] ^ uncoded_block[734];
  wire _8202 = _8200 ^ _8201;
  wire _8203 = _8199 ^ _8202;
  wire _8204 = uncoded_block[735] ^ uncoded_block[739];
  wire _8205 = _8204 ^ _352;
  wire _8206 = _5699 ^ _5702;
  wire _8207 = _8205 ^ _8206;
  wire _8208 = _8203 ^ _8207;
  wire _8209 = uncoded_block[747] ^ uncoded_block[750];
  wire _8210 = _8209 ^ _7013;
  wire _8211 = _5709 ^ _1218;
  wire _8212 = _8210 ^ _8211;
  wire _8213 = uncoded_block[773] ^ uncoded_block[777];
  wire _8214 = _8213 ^ _368;
  wire _8215 = uncoded_block[786] ^ uncoded_block[788];
  wire _8216 = _3568 ^ _8215;
  wire _8217 = _8214 ^ _8216;
  wire _8218 = _8212 ^ _8217;
  wire _8219 = _8208 ^ _8218;
  wire _8220 = _8197 ^ _8219;
  wire _8221 = _8171 ^ _8220;
  wire _8222 = _374 ^ _5723;
  wire _8223 = uncoded_block[797] ^ uncoded_block[798];
  wire _8224 = uncoded_block[799] ^ uncoded_block[802];
  wire _8225 = _8223 ^ _8224;
  wire _8226 = _8222 ^ _8225;
  wire _8227 = _3577 ^ _5727;
  wire _8228 = uncoded_block[809] ^ uncoded_block[811];
  wire _8229 = _8228 ^ _2026;
  wire _8230 = _8227 ^ _8229;
  wire _8231 = _8226 ^ _8230;
  wire _8232 = _4324 ^ _6398;
  wire _8233 = uncoded_block[820] ^ uncoded_block[825];
  wire _8234 = _8233 ^ _6401;
  wire _8235 = _8232 ^ _8234;
  wire _8236 = _3590 ^ _3597;
  wire _8237 = uncoded_block[853] ^ uncoded_block[854];
  wire _8238 = _3599 ^ _8237;
  wire _8239 = _8236 ^ _8238;
  wire _8240 = _8235 ^ _8239;
  wire _8241 = _8231 ^ _8240;
  wire _8242 = _408 ^ _6412;
  wire _8243 = uncoded_block[865] ^ uncoded_block[869];
  wire _8244 = uncoded_block[870] ^ uncoded_block[874];
  wire _8245 = _8243 ^ _8244;
  wire _8246 = _8242 ^ _8245;
  wire _8247 = uncoded_block[879] ^ uncoded_block[886];
  wire _8248 = uncoded_block[889] ^ uncoded_block[893];
  wire _8249 = _8247 ^ _8248;
  wire _8250 = uncoded_block[896] ^ uncoded_block[898];
  wire _8251 = _4355 ^ _8250;
  wire _8252 = _8249 ^ _8251;
  wire _8253 = _8246 ^ _8252;
  wire _8254 = uncoded_block[904] ^ uncoded_block[905];
  wire _8255 = _7066 ^ _8254;
  wire _8256 = uncoded_block[914] ^ uncoded_block[918];
  wire _8257 = _6428 ^ _8256;
  wire _8258 = _8255 ^ _8257;
  wire _8259 = uncoded_block[919] ^ uncoded_block[922];
  wire _8260 = uncoded_block[925] ^ uncoded_block[930];
  wire _8261 = _8259 ^ _8260;
  wire _8262 = uncoded_block[933] ^ uncoded_block[934];
  wire _8263 = _5096 ^ _8262;
  wire _8264 = _8261 ^ _8263;
  wire _8265 = _8258 ^ _8264;
  wire _8266 = _8253 ^ _8265;
  wire _8267 = _8241 ^ _8266;
  wire _8268 = uncoded_block[935] ^ uncoded_block[937];
  wire _8269 = uncoded_block[938] ^ uncoded_block[943];
  wire _8270 = _8268 ^ _8269;
  wire _8271 = uncoded_block[944] ^ uncoded_block[945];
  wire _8272 = _8271 ^ _5777;
  wire _8273 = _8270 ^ _8272;
  wire _8274 = uncoded_block[950] ^ uncoded_block[952];
  wire _8275 = uncoded_block[953] ^ uncoded_block[954];
  wire _8276 = _8274 ^ _8275;
  wire _8277 = uncoded_block[957] ^ uncoded_block[959];
  wire _8278 = _4384 ^ _8277;
  wire _8279 = _8276 ^ _8278;
  wire _8280 = _8273 ^ _8279;
  wire _8281 = _4385 ^ _2872;
  wire _8282 = uncoded_block[966] ^ uncoded_block[971];
  wire _8283 = uncoded_block[972] ^ uncoded_block[975];
  wire _8284 = _8282 ^ _8283;
  wire _8285 = _8281 ^ _8284;
  wire _8286 = uncoded_block[976] ^ uncoded_block[979];
  wire _8287 = uncoded_block[984] ^ uncoded_block[986];
  wire _8288 = _8286 ^ _8287;
  wire _8289 = _1318 ^ _1323;
  wire _8290 = _8288 ^ _8289;
  wire _8291 = _8285 ^ _8290;
  wire _8292 = _8280 ^ _8291;
  wire _8293 = uncoded_block[994] ^ uncoded_block[997];
  wire _8294 = _8293 ^ _5798;
  wire _8295 = uncoded_block[1004] ^ uncoded_block[1009];
  wire _8296 = uncoded_block[1012] ^ uncoded_block[1013];
  wire _8297 = _8295 ^ _8296;
  wire _8298 = _8294 ^ _8297;
  wire _8299 = uncoded_block[1021] ^ uncoded_block[1023];
  wire _8300 = _5134 ^ _8299;
  wire _8301 = uncoded_block[1024] ^ uncoded_block[1025];
  wire _8302 = _8301 ^ _498;
  wire _8303 = _8300 ^ _8302;
  wire _8304 = _8298 ^ _8303;
  wire _8305 = _3675 ^ _4418;
  wire _8306 = uncoded_block[1040] ^ uncoded_block[1043];
  wire _8307 = _502 ^ _8306;
  wire _8308 = _8305 ^ _8307;
  wire _8309 = uncoded_block[1045] ^ uncoded_block[1047];
  wire _8310 = _8309 ^ _2134;
  wire _8311 = uncoded_block[1055] ^ uncoded_block[1056];
  wire _8312 = _7714 ^ _8311;
  wire _8313 = _8310 ^ _8312;
  wire _8314 = _8308 ^ _8313;
  wire _8315 = _8304 ^ _8314;
  wire _8316 = _8292 ^ _8315;
  wire _8317 = _8267 ^ _8316;
  wire _8318 = _8221 ^ _8317;
  wire _8319 = _8129 ^ _8318;
  wire _8320 = _1363 ^ _4433;
  wire _8321 = _2142 ^ _5828;
  wire _8322 = _8320 ^ _8321;
  wire _8323 = _527 ^ _5831;
  wire _8324 = _5832 ^ _5834;
  wire _8325 = _8323 ^ _8324;
  wire _8326 = _8322 ^ _8325;
  wire _8327 = _7724 ^ _4438;
  wire _8328 = _1374 ^ _2930;
  wire _8329 = _8327 ^ _8328;
  wire _8330 = uncoded_block[1096] ^ uncoded_block[1099];
  wire _8331 = _3698 ^ _8330;
  wire _8332 = _545 ^ _3707;
  wire _8333 = _8331 ^ _8332;
  wire _8334 = _8329 ^ _8333;
  wire _8335 = _8326 ^ _8334;
  wire _8336 = uncoded_block[1106] ^ uncoded_block[1108];
  wire _8337 = uncoded_block[1112] ^ uncoded_block[1117];
  wire _8338 = _8336 ^ _8337;
  wire _8339 = uncoded_block[1118] ^ uncoded_block[1120];
  wire _8340 = _8339 ^ _4455;
  wire _8341 = _8338 ^ _8340;
  wire _8342 = uncoded_block[1123] ^ uncoded_block[1126];
  wire _8343 = uncoded_block[1129] ^ uncoded_block[1130];
  wire _8344 = _8342 ^ _8343;
  wire _8345 = uncoded_block[1133] ^ uncoded_block[1136];
  wire _8346 = uncoded_block[1137] ^ uncoded_block[1139];
  wire _8347 = _8345 ^ _8346;
  wire _8348 = _8344 ^ _8347;
  wire _8349 = _8341 ^ _8348;
  wire _8350 = _567 ^ _2953;
  wire _8351 = uncoded_block[1151] ^ uncoded_block[1153];
  wire _8352 = _5862 ^ _8351;
  wire _8353 = _8350 ^ _8352;
  wire _8354 = uncoded_block[1155] ^ uncoded_block[1156];
  wire _8355 = _8354 ^ _578;
  wire _8356 = uncoded_block[1161] ^ uncoded_block[1163];
  wire _8357 = _8356 ^ _4476;
  wire _8358 = _8355 ^ _8357;
  wire _8359 = _8353 ^ _8358;
  wire _8360 = _8349 ^ _8359;
  wire _8361 = _8335 ^ _8360;
  wire _8362 = uncoded_block[1171] ^ uncoded_block[1173];
  wire _8363 = _1408 ^ _8362;
  wire _8364 = _2967 ^ _590;
  wire _8365 = _8363 ^ _8364;
  wire _8366 = _2196 ^ _5203;
  wire _8367 = _6525 ^ _7160;
  wire _8368 = _8366 ^ _8367;
  wire _8369 = _8365 ^ _8368;
  wire _8370 = uncoded_block[1200] ^ uncoded_block[1202];
  wire _8371 = uncoded_block[1203] ^ uncoded_block[1206];
  wire _8372 = _8370 ^ _8371;
  wire _8373 = uncoded_block[1211] ^ uncoded_block[1218];
  wire _8374 = _2217 ^ _8373;
  wire _8375 = _8372 ^ _8374;
  wire _8376 = _5215 ^ _5891;
  wire _8377 = uncoded_block[1227] ^ uncoded_block[1229];
  wire _8378 = _8377 ^ _1442;
  wire _8379 = _8376 ^ _8378;
  wire _8380 = _8375 ^ _8379;
  wire _8381 = _8369 ^ _8380;
  wire _8382 = uncoded_block[1239] ^ uncoded_block[1243];
  wire _8383 = _2989 ^ _8382;
  wire _8384 = uncoded_block[1244] ^ uncoded_block[1248];
  wire _8385 = uncoded_block[1250] ^ uncoded_block[1251];
  wire _8386 = _8384 ^ _8385;
  wire _8387 = _8383 ^ _8386;
  wire _8388 = uncoded_block[1252] ^ uncoded_block[1254];
  wire _8389 = uncoded_block[1255] ^ uncoded_block[1259];
  wire _8390 = _8388 ^ _8389;
  wire _8391 = uncoded_block[1263] ^ uncoded_block[1267];
  wire _8392 = _2238 ^ _8391;
  wire _8393 = _8390 ^ _8392;
  wire _8394 = _8387 ^ _8393;
  wire _8395 = _7179 ^ _3010;
  wire _8396 = uncoded_block[1285] ^ uncoded_block[1290];
  wire _8397 = _5241 ^ _8396;
  wire _8398 = _8395 ^ _8397;
  wire _8399 = uncoded_block[1291] ^ uncoded_block[1293];
  wire _8400 = _8399 ^ _3015;
  wire _8401 = _4532 ^ _2255;
  wire _8402 = _8400 ^ _8401;
  wire _8403 = _8398 ^ _8402;
  wire _8404 = _8394 ^ _8403;
  wire _8405 = _8381 ^ _8404;
  wire _8406 = _8361 ^ _8405;
  wire _8407 = uncoded_block[1310] ^ uncoded_block[1312];
  wire _8408 = _3807 ^ _8407;
  wire _8409 = _3026 ^ _5254;
  wire _8410 = _8408 ^ _8409;
  wire _8411 = uncoded_block[1324] ^ uncoded_block[1325];
  wire _8412 = _8411 ^ _1490;
  wire _8413 = uncoded_block[1333] ^ uncoded_block[1334];
  wire _8414 = _8413 ^ _1497;
  wire _8415 = _8412 ^ _8414;
  wire _8416 = _8410 ^ _8415;
  wire _8417 = uncoded_block[1344] ^ uncoded_block[1348];
  wire _8418 = uncoded_block[1350] ^ uncoded_block[1353];
  wire _8419 = _8417 ^ _8418;
  wire _8420 = _6587 ^ _5273;
  wire _8421 = _8419 ^ _8420;
  wire _8422 = _2283 ^ _3052;
  wire _8423 = uncoded_block[1371] ^ uncoded_block[1372];
  wire _8424 = _8423 ^ _2289;
  wire _8425 = _8422 ^ _8424;
  wire _8426 = _8421 ^ _8425;
  wire _8427 = _8416 ^ _8426;
  wire _8428 = _3834 ^ _7222;
  wire _8429 = _5286 ^ _8428;
  wire _8430 = uncoded_block[1393] ^ uncoded_block[1397];
  wire _8431 = _691 ^ _8430;
  wire _8432 = _4572 ^ _2297;
  wire _8433 = _8431 ^ _8432;
  wire _8434 = _8429 ^ _8433;
  wire _8435 = uncoded_block[1404] ^ uncoded_block[1407];
  wire _8436 = uncoded_block[1409] ^ uncoded_block[1410];
  wire _8437 = _8435 ^ _8436;
  wire _8438 = uncoded_block[1415] ^ uncoded_block[1416];
  wire _8439 = _8438 ^ _705;
  wire _8440 = _8437 ^ _8439;
  wire _8441 = uncoded_block[1419] ^ uncoded_block[1424];
  wire _8442 = _8441 ^ _3075;
  wire _8443 = uncoded_block[1433] ^ uncoded_block[1436];
  wire _8444 = _1531 ^ _8443;
  wire _8445 = _8442 ^ _8444;
  wire _8446 = _8440 ^ _8445;
  wire _8447 = _8434 ^ _8446;
  wire _8448 = _8427 ^ _8447;
  wire _8449 = uncoded_block[1440] ^ uncoded_block[1445];
  wire _8450 = uncoded_block[1446] ^ uncoded_block[1448];
  wire _8451 = _8449 ^ _8450;
  wire _8452 = uncoded_block[1459] ^ uncoded_block[1462];
  wire _8453 = _5978 ^ _8452;
  wire _8454 = _8451 ^ _8453;
  wire _8455 = uncoded_block[1463] ^ uncoded_block[1464];
  wire _8456 = uncoded_block[1465] ^ uncoded_block[1471];
  wire _8457 = _8455 ^ _8456;
  wire _8458 = _3881 ^ _3884;
  wire _8459 = _8457 ^ _8458;
  wire _8460 = _8454 ^ _8459;
  wire _8461 = uncoded_block[1484] ^ uncoded_block[1489];
  wire _8462 = uncoded_block[1491] ^ uncoded_block[1495];
  wire _8463 = _8461 ^ _8462;
  wire _8464 = _743 ^ _747;
  wire _8465 = _8463 ^ _8464;
  wire _8466 = _4614 ^ _7259;
  wire _8467 = uncoded_block[1509] ^ uncoded_block[1515];
  wire _8468 = _3112 ^ _8467;
  wire _8469 = _8466 ^ _8468;
  wire _8470 = _8465 ^ _8469;
  wire _8471 = _8460 ^ _8470;
  wire _8472 = _5337 ^ _7269;
  wire _8473 = uncoded_block[1524] ^ uncoded_block[1525];
  wire _8474 = uncoded_block[1529] ^ uncoded_block[1530];
  wire _8475 = _8473 ^ _8474;
  wire _8476 = _8472 ^ _8475;
  wire _8477 = _5347 ^ _3906;
  wire _8478 = uncoded_block[1538] ^ uncoded_block[1541];
  wire _8479 = _8478 ^ _1590;
  wire _8480 = _8477 ^ _8479;
  wire _8481 = _8476 ^ _8480;
  wire _8482 = uncoded_block[1548] ^ uncoded_block[1549];
  wire _8483 = _2367 ^ _8482;
  wire _8484 = uncoded_block[1555] ^ uncoded_block[1560];
  wire _8485 = _7277 ^ _8484;
  wire _8486 = _8483 ^ _8485;
  wire _8487 = _774 ^ _5361;
  wire _8488 = _7891 ^ _6028;
  wire _8489 = _8487 ^ _8488;
  wire _8490 = _8486 ^ _8489;
  wire _8491 = _8481 ^ _8490;
  wire _8492 = _8471 ^ _8491;
  wire _8493 = _8448 ^ _8492;
  wire _8494 = _8406 ^ _8493;
  wire _8495 = _784 ^ _2386;
  wire _8496 = uncoded_block[1589] ^ uncoded_block[1593];
  wire _8497 = _8496 ^ _4654;
  wire _8498 = _8495 ^ _8497;
  wire _8499 = uncoded_block[1596] ^ uncoded_block[1598];
  wire _8500 = uncoded_block[1599] ^ uncoded_block[1602];
  wire _8501 = _8499 ^ _8500;
  wire _8502 = uncoded_block[1603] ^ uncoded_block[1604];
  wire _8503 = _8502 ^ _1625;
  wire _8504 = _8501 ^ _8503;
  wire _8505 = _8498 ^ _8504;
  wire _8506 = _1627 ^ _3937;
  wire _8507 = _8506 ^ _6681;
  wire _8508 = _6684 ^ _6046;
  wire _8509 = uncoded_block[1627] ^ uncoded_block[1631];
  wire _8510 = _8509 ^ _6049;
  wire _8511 = _8508 ^ _8510;
  wire _8512 = _8507 ^ _8511;
  wire _8513 = _8505 ^ _8512;
  wire _8514 = _3951 ^ _816;
  wire _8515 = uncoded_block[1653] ^ uncoded_block[1656];
  wire _8516 = _819 ^ _8515;
  wire _8517 = _8514 ^ _8516;
  wire _8518 = _4681 ^ _4686;
  wire _8519 = _8517 ^ _8518;
  wire _8520 = _4687 ^ _7928;
  wire _8521 = uncoded_block[1671] ^ uncoded_block[1672];
  wire _8522 = uncoded_block[1673] ^ uncoded_block[1675];
  wire _8523 = _8521 ^ _8522;
  wire _8524 = _8520 ^ _8523;
  wire _8525 = _833 ^ _3187;
  wire _8526 = uncoded_block[1687] ^ uncoded_block[1692];
  wire _8527 = uncoded_block[1693] ^ uncoded_block[1696];
  wire _8528 = _8526 ^ _8527;
  wire _8529 = _8525 ^ _8528;
  wire _8530 = _8524 ^ _8529;
  wire _8531 = _8519 ^ _8530;
  wire _8532 = _8513 ^ _8531;
  wire _8533 = uncoded_block[1699] ^ uncoded_block[1701];
  wire _8534 = _5409 ^ _8533;
  wire _8535 = uncoded_block[1703] ^ uncoded_block[1704];
  wire _8536 = uncoded_block[1706] ^ uncoded_block[1708];
  wire _8537 = _8535 ^ _8536;
  wire _8538 = _8534 ^ _8537;
  wire _8539 = _2441 ^ uncoded_block[1721];
  wire _8540 = _8538 ^ _8539;
  wire _8541 = _8532 ^ _8540;
  wire _8542 = _8494 ^ _8541;
  wire _8543 = _8319 ^ _8542;
  wire _8544 = _4712 ^ _6083;
  wire _8545 = uncoded_block[15] ^ uncoded_block[17];
  wire _8546 = _4713 ^ _8545;
  wire _8547 = _8544 ^ _8546;
  wire _8548 = uncoded_block[30] ^ uncoded_block[35];
  wire _8549 = uncoded_block[36] ^ uncoded_block[37];
  wire _8550 = _8548 ^ _8549;
  wire _8551 = _19 ^ _22;
  wire _8552 = _8550 ^ _8551;
  wire _8553 = _8547 ^ _8552;
  wire _8554 = uncoded_block[46] ^ uncoded_block[47];
  wire _8555 = _8554 ^ _3232;
  wire _8556 = uncoded_block[51] ^ uncoded_block[54];
  wire _8557 = _8556 ^ _7969;
  wire _8558 = _8555 ^ _8557;
  wire _8559 = uncoded_block[63] ^ uncoded_block[67];
  wire _8560 = _31 ^ _8559;
  wire _8561 = _7367 ^ _5442;
  wire _8562 = _8560 ^ _8561;
  wire _8563 = _8558 ^ _8562;
  wire _8564 = _8553 ^ _8563;
  wire _8565 = _1714 ^ _6754;
  wire _8566 = uncoded_block[89] ^ uncoded_block[91];
  wire _8567 = uncoded_block[93] ^ uncoded_block[95];
  wire _8568 = _8566 ^ _8567;
  wire _8569 = _8565 ^ _8568;
  wire _8570 = uncoded_block[100] ^ uncoded_block[106];
  wire _8571 = _7375 ^ _8570;
  wire _8572 = uncoded_block[107] ^ uncoded_block[109];
  wire _8573 = _8572 ^ _1726;
  wire _8574 = _8571 ^ _8573;
  wire _8575 = _8569 ^ _8574;
  wire _8576 = _2495 ^ _2497;
  wire _8577 = _3255 ^ _2502;
  wire _8578 = _8576 ^ _8577;
  wire _8579 = uncoded_block[129] ^ uncoded_block[131];
  wire _8580 = _4753 ^ _8579;
  wire _8581 = uncoded_block[135] ^ uncoded_block[136];
  wire _8582 = _8581 ^ _66;
  wire _8583 = _8580 ^ _8582;
  wire _8584 = _8578 ^ _8583;
  wire _8585 = _8575 ^ _8584;
  wire _8586 = _8564 ^ _8585;
  wire _8587 = _1744 ^ _3269;
  wire _8588 = _8587 ^ _2515;
  wire _8589 = uncoded_block[165] ^ uncoded_block[166];
  wire _8590 = _1749 ^ _8589;
  wire _8591 = uncoded_block[170] ^ uncoded_block[171];
  wire _8592 = _8591 ^ _938;
  wire _8593 = _8590 ^ _8592;
  wire _8594 = _8588 ^ _8593;
  wire _8595 = uncoded_block[175] ^ uncoded_block[178];
  wire _8596 = _8595 ^ _2528;
  wire _8597 = uncoded_block[188] ^ uncoded_block[194];
  wire _8598 = _8597 ^ _3289;
  wire _8599 = _8596 ^ _8598;
  wire _8600 = uncoded_block[207] ^ uncoded_block[208];
  wire _8601 = _4070 ^ _8600;
  wire _8602 = _7415 ^ _2540;
  wire _8603 = _8601 ^ _8602;
  wire _8604 = _8599 ^ _8603;
  wire _8605 = _8594 ^ _8604;
  wire _8606 = uncoded_block[216] ^ uncoded_block[218];
  wire _8607 = _8606 ^ _102;
  wire _8608 = uncoded_block[224] ^ uncoded_block[227];
  wire _8609 = _5497 ^ _8608;
  wire _8610 = _8607 ^ _8609;
  wire _8611 = _6169 ^ _1775;
  wire _8612 = uncoded_block[239] ^ uncoded_block[243];
  wire _8613 = _3305 ^ _8612;
  wire _8614 = _8611 ^ _8613;
  wire _8615 = _8610 ^ _8614;
  wire _8616 = uncoded_block[245] ^ uncoded_block[246];
  wire _8617 = uncoded_block[247] ^ uncoded_block[248];
  wire _8618 = _8616 ^ _8617;
  wire _8619 = uncoded_block[249] ^ uncoded_block[254];
  wire _8620 = uncoded_block[256] ^ uncoded_block[259];
  wire _8621 = _8619 ^ _8620;
  wire _8622 = _8618 ^ _8621;
  wire _8623 = uncoded_block[263] ^ uncoded_block[268];
  wire _8624 = _6185 ^ _8623;
  wire _8625 = _3320 ^ _4813;
  wire _8626 = _8624 ^ _8625;
  wire _8627 = _8622 ^ _8626;
  wire _8628 = _8615 ^ _8627;
  wire _8629 = _8605 ^ _8628;
  wire _8630 = _8586 ^ _8629;
  wire _8631 = _6834 ^ _7446;
  wire _8632 = uncoded_block[285] ^ uncoded_block[286];
  wire _8633 = uncoded_block[292] ^ uncoded_block[294];
  wire _8634 = _8632 ^ _8633;
  wire _8635 = _8631 ^ _8634;
  wire _8636 = uncoded_block[299] ^ uncoded_block[300];
  wire _8637 = uncoded_block[301] ^ uncoded_block[305];
  wire _8638 = _8636 ^ _8637;
  wire _8639 = _8055 ^ _6206;
  wire _8640 = _8638 ^ _8639;
  wire _8641 = _8635 ^ _8640;
  wire _8642 = uncoded_block[323] ^ uncoded_block[325];
  wire _8643 = _1818 ^ _8642;
  wire _8644 = _4831 ^ _8643;
  wire _8645 = _1014 ^ _6853;
  wire _8646 = uncoded_block[335] ^ uncoded_block[337];
  wire _8647 = _8646 ^ _2593;
  wire _8648 = _8645 ^ _8647;
  wire _8649 = _8644 ^ _8648;
  wire _8650 = _8641 ^ _8649;
  wire _8651 = _1021 ^ _6218;
  wire _8652 = uncoded_block[346] ^ uncoded_block[348];
  wire _8653 = _8652 ^ _2601;
  wire _8654 = _8651 ^ _8653;
  wire _8655 = uncoded_block[366] ^ uncoded_block[369];
  wire _8656 = _8655 ^ _6873;
  wire _8657 = _3367 ^ _8656;
  wire _8658 = _8654 ^ _8657;
  wire _8659 = uncoded_block[379] ^ uncoded_block[383];
  wire _8660 = _4853 ^ _8659;
  wire _8661 = uncoded_block[393] ^ uncoded_block[396];
  wire _8662 = _4149 ^ _8661;
  wire _8663 = _8660 ^ _8662;
  wire _8664 = _2629 ^ _3394;
  wire _8665 = uncoded_block[418] ^ uncoded_block[422];
  wire _8666 = _1055 ^ _8665;
  wire _8667 = _8664 ^ _8666;
  wire _8668 = _8663 ^ _8667;
  wire _8669 = _8658 ^ _8668;
  wire _8670 = _8650 ^ _8669;
  wire _8671 = uncoded_block[423] ^ uncoded_block[424];
  wire _8672 = uncoded_block[425] ^ uncoded_block[426];
  wire _8673 = _8671 ^ _8672;
  wire _8674 = uncoded_block[428] ^ uncoded_block[433];
  wire _8675 = _8674 ^ _6255;
  wire _8676 = _8673 ^ _8675;
  wire _8677 = _1863 ^ _5578;
  wire _8678 = _1864 ^ _1866;
  wire _8679 = _8677 ^ _8678;
  wire _8680 = _8676 ^ _8679;
  wire _8681 = uncoded_block[459] ^ uncoded_block[460];
  wire _8682 = _1867 ^ _8681;
  wire _8683 = uncoded_block[465] ^ uncoded_block[466];
  wire _8684 = _4181 ^ _8683;
  wire _8685 = _8682 ^ _8684;
  wire _8686 = uncoded_block[470] ^ uncoded_block[472];
  wire _8687 = _1878 ^ _8686;
  wire _8688 = uncoded_block[476] ^ uncoded_block[478];
  wire _8689 = _1083 ^ _8688;
  wire _8690 = _8687 ^ _8689;
  wire _8691 = _8685 ^ _8690;
  wire _8692 = _8680 ^ _8691;
  wire _8693 = uncoded_block[479] ^ uncoded_block[482];
  wire _8694 = uncoded_block[484] ^ uncoded_block[486];
  wire _8695 = _8693 ^ _8694;
  wire _8696 = _4194 ^ _4902;
  wire _8697 = _8695 ^ _8696;
  wire _8698 = uncoded_block[497] ^ uncoded_block[500];
  wire _8699 = _5603 ^ _8698;
  wire _8700 = uncoded_block[501] ^ uncoded_block[505];
  wire _8701 = uncoded_block[507] ^ uncoded_block[510];
  wire _8702 = _8700 ^ _8701;
  wire _8703 = _8699 ^ _8702;
  wire _8704 = _8697 ^ _8703;
  wire _8705 = uncoded_block[511] ^ uncoded_block[513];
  wire _8706 = uncoded_block[515] ^ uncoded_block[516];
  wire _8707 = _8705 ^ _8706;
  wire _8708 = uncoded_block[519] ^ uncoded_block[522];
  wire _8709 = _8708 ^ _6289;
  wire _8710 = _8707 ^ _8709;
  wire _8711 = _4214 ^ _6932;
  wire _8712 = _4923 ^ _8711;
  wire _8713 = _8710 ^ _8712;
  wire _8714 = _8704 ^ _8713;
  wire _8715 = _8692 ^ _8714;
  wire _8716 = _8670 ^ _8715;
  wire _8717 = _8630 ^ _8716;
  wire _8718 = uncoded_block[539] ^ uncoded_block[542];
  wire _8719 = _8718 ^ _244;
  wire _8720 = uncoded_block[549] ^ uncoded_block[552];
  wire _8721 = uncoded_block[553] ^ uncoded_block[554];
  wire _8722 = _8720 ^ _8721;
  wire _8723 = _8719 ^ _8722;
  wire _8724 = uncoded_block[555] ^ uncoded_block[556];
  wire _8725 = uncoded_block[559] ^ uncoded_block[564];
  wire _8726 = _8724 ^ _8725;
  wire _8727 = uncoded_block[568] ^ uncoded_block[571];
  wire _8728 = _5635 ^ _8727;
  wire _8729 = _8726 ^ _8728;
  wire _8730 = _8723 ^ _8729;
  wire _8731 = uncoded_block[574] ^ uncoded_block[576];
  wire _8732 = _8731 ^ _263;
  wire _8733 = uncoded_block[584] ^ uncoded_block[586];
  wire _8734 = _265 ^ _8733;
  wire _8735 = _8732 ^ _8734;
  wire _8736 = uncoded_block[598] ^ uncoded_block[601];
  wire _8737 = _1939 ^ _8736;
  wire _8738 = uncoded_block[603] ^ uncoded_block[605];
  wire _8739 = uncoded_block[607] ^ uncoded_block[611];
  wire _8740 = _8738 ^ _8739;
  wire _8741 = _8737 ^ _8740;
  wire _8742 = _8735 ^ _8741;
  wire _8743 = _8730 ^ _8742;
  wire _8744 = uncoded_block[613] ^ uncoded_block[615];
  wire _8745 = uncoded_block[616] ^ uncoded_block[619];
  wire _8746 = _8744 ^ _8745;
  wire _8747 = _1946 ^ _1948;
  wire _8748 = _8746 ^ _8747;
  wire _8749 = uncoded_block[628] ^ uncoded_block[633];
  wire _8750 = _8749 ^ _7577;
  wire _8751 = uncoded_block[642] ^ uncoded_block[644];
  wire _8752 = _1163 ^ _8751;
  wire _8753 = _8750 ^ _8752;
  wire _8754 = _8748 ^ _8753;
  wire _8755 = uncoded_block[655] ^ uncoded_block[659];
  wire _8756 = _296 ^ _8755;
  wire _8757 = _3514 ^ _4978;
  wire _8758 = _8756 ^ _8757;
  wire _8759 = _309 ^ _4982;
  wire _8760 = uncoded_block[674] ^ uncoded_block[676];
  wire _8761 = uncoded_block[677] ^ uncoded_block[680];
  wire _8762 = _8760 ^ _8761;
  wire _8763 = _8759 ^ _8762;
  wire _8764 = _8758 ^ _8763;
  wire _8765 = _8754 ^ _8764;
  wire _8766 = _8743 ^ _8765;
  wire _8767 = uncoded_block[691] ^ uncoded_block[696];
  wire _8768 = _6353 ^ _8767;
  wire _8769 = _6992 ^ _3533;
  wire _8770 = _8768 ^ _8769;
  wire _8771 = _4996 ^ _5002;
  wire _8772 = _5690 ^ _4283;
  wire _8773 = _8771 ^ _8772;
  wire _8774 = _8770 ^ _8773;
  wire _8775 = uncoded_block[736] ^ uncoded_block[739];
  wire _8776 = _8775 ^ _352;
  wire _8777 = _3548 ^ _8776;
  wire _8778 = uncoded_block[747] ^ uncoded_block[751];
  wire _8779 = uncoded_block[752] ^ uncoded_block[755];
  wire _8780 = _8778 ^ _8779;
  wire _8781 = uncoded_block[761] ^ uncoded_block[762];
  wire _8782 = _3556 ^ _8781;
  wire _8783 = _8780 ^ _8782;
  wire _8784 = _8777 ^ _8783;
  wire _8785 = _8774 ^ _8784;
  wire _8786 = _365 ^ _5027;
  wire _8787 = uncoded_block[772] ^ uncoded_block[776];
  wire _8788 = _8787 ^ _3568;
  wire _8789 = _8786 ^ _8788;
  wire _8790 = uncoded_block[787] ^ uncoded_block[789];
  wire _8791 = uncoded_block[791] ^ uncoded_block[794];
  wire _8792 = _8790 ^ _8791;
  wire _8793 = uncoded_block[804] ^ uncoded_block[806];
  wire _8794 = _4317 ^ _8793;
  wire _8795 = _8792 ^ _8794;
  wire _8796 = _8789 ^ _8795;
  wire _8797 = _5043 ^ _5047;
  wire _8798 = uncoded_block[821] ^ uncoded_block[826];
  wire _8799 = _1242 ^ _8798;
  wire _8800 = uncoded_block[828] ^ uncoded_block[831];
  wire _8801 = _8800 ^ _4331;
  wire _8802 = _8799 ^ _8801;
  wire _8803 = _8797 ^ _8802;
  wire _8804 = _8796 ^ _8803;
  wire _8805 = _8785 ^ _8804;
  wire _8806 = _8766 ^ _8805;
  wire _8807 = _4336 ^ _7043;
  wire _8808 = uncoded_block[843] ^ uncoded_block[845];
  wire _8809 = uncoded_block[850] ^ uncoded_block[852];
  wire _8810 = _8808 ^ _8809;
  wire _8811 = _8807 ^ _8810;
  wire _8812 = uncoded_block[856] ^ uncoded_block[857];
  wire _8813 = _8237 ^ _8812;
  wire _8814 = _408 ^ _413;
  wire _8815 = _8813 ^ _8814;
  wire _8816 = _8811 ^ _8815;
  wire _8817 = uncoded_block[864] ^ uncoded_block[869];
  wire _8818 = _8817 ^ _8244;
  wire _8819 = _8818 ^ _3609;
  wire _8820 = uncoded_block[882] ^ uncoded_block[884];
  wire _8821 = _8820 ^ _5082;
  wire _8822 = _4354 ^ _1277;
  wire _8823 = _8821 ^ _8822;
  wire _8824 = _8819 ^ _8823;
  wire _8825 = _8816 ^ _8824;
  wire _8826 = uncoded_block[897] ^ uncoded_block[899];
  wire _8827 = uncoded_block[901] ^ uncoded_block[905];
  wire _8828 = _8826 ^ _8827;
  wire _8829 = uncoded_block[906] ^ uncoded_block[911];
  wire _8830 = _8829 ^ _5762;
  wire _8831 = _8828 ^ _8830;
  wire _8832 = uncoded_block[918] ^ uncoded_block[924];
  wire _8833 = _3628 ^ _8832;
  wire _8834 = uncoded_block[926] ^ uncoded_block[928];
  wire _8835 = uncoded_block[929] ^ uncoded_block[931];
  wire _8836 = _8834 ^ _8835;
  wire _8837 = _8833 ^ _8836;
  wire _8838 = _8831 ^ _8837;
  wire _8839 = uncoded_block[937] ^ uncoded_block[940];
  wire _8840 = _1299 ^ _8839;
  wire _8841 = uncoded_block[943] ^ uncoded_block[948];
  wire _8842 = uncoded_block[950] ^ uncoded_block[953];
  wire _8843 = _8841 ^ _8842;
  wire _8844 = _8840 ^ _8843;
  wire _8845 = uncoded_block[957] ^ uncoded_block[963];
  wire _8846 = _8845 ^ _2092;
  wire _8847 = uncoded_block[970] ^ uncoded_block[972];
  wire _8848 = _5785 ^ _8847;
  wire _8849 = _8846 ^ _8848;
  wire _8850 = _8844 ^ _8849;
  wire _8851 = _8838 ^ _8850;
  wire _8852 = _8825 ^ _8851;
  wire _8853 = uncoded_block[979] ^ uncoded_block[981];
  wire _8854 = _5114 ^ _8853;
  wire _8855 = uncoded_block[982] ^ uncoded_block[984];
  wire _8856 = uncoded_block[987] ^ uncoded_block[988];
  wire _8857 = _8855 ^ _8856;
  wire _8858 = _8854 ^ _8857;
  wire _8859 = uncoded_block[989] ^ uncoded_block[991];
  wire _8860 = uncoded_block[993] ^ uncoded_block[995];
  wire _8861 = _8859 ^ _8860;
  wire _8862 = uncoded_block[996] ^ uncoded_block[1000];
  wire _8863 = _8862 ^ _483;
  wire _8864 = _8861 ^ _8863;
  wire _8865 = _8858 ^ _8864;
  wire _8866 = uncoded_block[1004] ^ uncoded_block[1006];
  wire _8867 = _8866 ^ _5129;
  wire _8868 = uncoded_block[1013] ^ uncoded_block[1017];
  wire _8869 = _4410 ^ _8868;
  wire _8870 = _8867 ^ _8869;
  wire _8871 = uncoded_block[1018] ^ uncoded_block[1019];
  wire _8872 = uncoded_block[1022] ^ uncoded_block[1025];
  wire _8873 = _8871 ^ _8872;
  wire _8874 = uncoded_block[1026] ^ uncoded_block[1027];
  wire _8875 = uncoded_block[1028] ^ uncoded_block[1029];
  wire _8876 = _8874 ^ _8875;
  wire _8877 = _8873 ^ _8876;
  wire _8878 = _8870 ^ _8877;
  wire _8879 = _8865 ^ _8878;
  wire _8880 = _499 ^ _2127;
  wire _8881 = _1342 ^ _1345;
  wire _8882 = _8880 ^ _8881;
  wire _8883 = _6478 ^ _2910;
  wire _8884 = uncoded_block[1053] ^ uncoded_block[1056];
  wire _8885 = _2134 ^ _8884;
  wire _8886 = _8883 ^ _8885;
  wire _8887 = _8882 ^ _8886;
  wire _8888 = uncoded_block[1064] ^ uncoded_block[1065];
  wire _8889 = uncoded_block[1066] ^ uncoded_block[1067];
  wire _8890 = _8888 ^ _8889;
  wire _8891 = _2141 ^ _8890;
  wire _8892 = uncoded_block[1070] ^ uncoded_block[1071];
  wire _8893 = uncoded_block[1073] ^ uncoded_block[1075];
  wire _8894 = _8892 ^ _8893;
  wire _8895 = uncoded_block[1077] ^ uncoded_block[1078];
  wire _8896 = _8895 ^ _5834;
  wire _8897 = _8894 ^ _8896;
  wire _8898 = _8891 ^ _8897;
  wire _8899 = _8887 ^ _8898;
  wire _8900 = _8879 ^ _8899;
  wire _8901 = _8852 ^ _8900;
  wire _8902 = _8806 ^ _8901;
  wire _8903 = _8717 ^ _8902;
  wire _8904 = uncoded_block[1081] ^ uncoded_block[1083];
  wire _8905 = _8904 ^ _4438;
  wire _8906 = uncoded_block[1089] ^ uncoded_block[1091];
  wire _8907 = _2149 ^ _8906;
  wire _8908 = _8905 ^ _8907;
  wire _8909 = _3698 ^ _3704;
  wire _8910 = uncoded_block[1101] ^ uncoded_block[1102];
  wire _8911 = _5169 ^ _8910;
  wire _8912 = _8909 ^ _8911;
  wire _8913 = _8908 ^ _8912;
  wire _8914 = uncoded_block[1104] ^ uncoded_block[1106];
  wire _8915 = uncoded_block[1107] ^ uncoded_block[1109];
  wire _8916 = _8914 ^ _8915;
  wire _8917 = uncoded_block[1112] ^ uncoded_block[1113];
  wire _8918 = _7132 ^ _8917;
  wire _8919 = _8916 ^ _8918;
  wire _8920 = uncoded_block[1118] ^ uncoded_block[1119];
  wire _8921 = _8920 ^ _7736;
  wire _8922 = _3718 ^ _4459;
  wire _8923 = _8921 ^ _8922;
  wire _8924 = _8919 ^ _8923;
  wire _8925 = _8913 ^ _8924;
  wire _8926 = _6499 ^ _560;
  wire _8927 = _561 ^ _5856;
  wire _8928 = _8926 ^ _8927;
  wire _8929 = uncoded_block[1136] ^ uncoded_block[1137];
  wire _8930 = uncoded_block[1139] ^ uncoded_block[1142];
  wire _8931 = _8929 ^ _8930;
  wire _8932 = uncoded_block[1145] ^ uncoded_block[1146];
  wire _8933 = uncoded_block[1149] ^ uncoded_block[1152];
  wire _8934 = _8932 ^ _8933;
  wire _8935 = _8931 ^ _8934;
  wire _8936 = _8928 ^ _8935;
  wire _8937 = uncoded_block[1153] ^ uncoded_block[1154];
  wire _8938 = uncoded_block[1155] ^ uncoded_block[1160];
  wire _8939 = _8937 ^ _8938;
  wire _8940 = uncoded_block[1161] ^ uncoded_block[1170];
  wire _8941 = _8940 ^ _7154;
  wire _8942 = _8939 ^ _8941;
  wire _8943 = _5195 ^ _3742;
  wire _8944 = uncoded_block[1181] ^ uncoded_block[1184];
  wire _8945 = _8944 ^ _2200;
  wire _8946 = _8943 ^ _8945;
  wire _8947 = _8942 ^ _8946;
  wire _8948 = _8936 ^ _8947;
  wire _8949 = _8925 ^ _8948;
  wire _8950 = _1420 ^ _6525;
  wire _8951 = uncoded_block[1197] ^ uncoded_block[1198];
  wire _8952 = _8951 ^ _7162;
  wire _8953 = _8950 ^ _8952;
  wire _8954 = _8371 ^ _2216;
  wire _8955 = _8954 ^ _2983;
  wire _8956 = _8953 ^ _8955;
  wire _8957 = _605 ^ _608;
  wire _8958 = uncoded_block[1223] ^ uncoded_block[1225];
  wire _8959 = _8958 ^ _1439;
  wire _8960 = _8957 ^ _8959;
  wire _8961 = _5219 ^ _7174;
  wire _8962 = uncoded_block[1239] ^ uncoded_block[1241];
  wire _8963 = uncoded_block[1243] ^ uncoded_block[1246];
  wire _8964 = _8962 ^ _8963;
  wire _8965 = _8961 ^ _8964;
  wire _8966 = _8960 ^ _8965;
  wire _8967 = _8956 ^ _8966;
  wire _8968 = uncoded_block[1251] ^ uncoded_block[1256];
  wire _8969 = _1451 ^ _8968;
  wire _8970 = uncoded_block[1259] ^ uncoded_block[1262];
  wire _8971 = _8970 ^ _6550;
  wire _8972 = _8969 ^ _8971;
  wire _8973 = _2239 ^ _2244;
  wire _8974 = uncoded_block[1272] ^ uncoded_block[1277];
  wire _8975 = _2245 ^ _8974;
  wire _8976 = _8973 ^ _8975;
  wire _8977 = _8972 ^ _8976;
  wire _8978 = uncoded_block[1280] ^ uncoded_block[1285];
  wire _8979 = _3793 ^ _8978;
  wire _8980 = uncoded_block[1288] ^ uncoded_block[1290];
  wire _8981 = uncoded_block[1291] ^ uncoded_block[1296];
  wire _8982 = _8980 ^ _8981;
  wire _8983 = _8979 ^ _8982;
  wire _8984 = uncoded_block[1300] ^ uncoded_block[1301];
  wire _8985 = _3017 ^ _8984;
  wire _8986 = _8985 ^ _2256;
  wire _8987 = _8983 ^ _8986;
  wire _8988 = _8977 ^ _8987;
  wire _8989 = _8967 ^ _8988;
  wire _8990 = _8949 ^ _8989;
  wire _8991 = uncoded_block[1306] ^ uncoded_block[1307];
  wire _8992 = uncoded_block[1308] ^ uncoded_block[1310];
  wire _8993 = _8991 ^ _8992;
  wire _8994 = uncoded_block[1324] ^ uncoded_block[1327];
  wire _8995 = _3028 ^ _8994;
  wire _8996 = _8993 ^ _8995;
  wire _8997 = uncoded_block[1328] ^ uncoded_block[1330];
  wire _8998 = uncoded_block[1331] ^ uncoded_block[1332];
  wire _8999 = _8997 ^ _8998;
  wire _9000 = _8413 ^ _661;
  wire _9001 = _8999 ^ _9000;
  wire _9002 = _8996 ^ _9001;
  wire _9003 = uncoded_block[1344] ^ uncoded_block[1346];
  wire _9004 = _1497 ^ _9003;
  wire _9005 = _5268 ^ _3041;
  wire _9006 = _9004 ^ _9005;
  wire _9007 = _3045 ^ _7211;
  wire _9008 = _674 ^ _9007;
  wire _9009 = _9006 ^ _9008;
  wire _9010 = _9002 ^ _9009;
  wire _9011 = _3047 ^ _680;
  wire _9012 = uncoded_block[1376] ^ uncoded_block[1383];
  wire _9013 = _7823 ^ _9012;
  wire _9014 = _9011 ^ _9013;
  wire _9015 = _4569 ^ _4571;
  wire _9016 = uncoded_block[1401] ^ uncoded_block[1403];
  wire _9017 = _9016 ^ _4578;
  wire _9018 = _9015 ^ _9017;
  wire _9019 = _9014 ^ _9018;
  wire _9020 = _8436 ^ _704;
  wire _9021 = uncoded_block[1419] ^ uncoded_block[1421];
  wire _9022 = uncoded_block[1422] ^ uncoded_block[1424];
  wire _9023 = _9021 ^ _9022;
  wire _9024 = _9020 ^ _9023;
  wire _9025 = uncoded_block[1426] ^ uncoded_block[1430];
  wire _9026 = _9025 ^ _1533;
  wire _9027 = uncoded_block[1434] ^ uncoded_block[1439];
  wire _9028 = _9027 ^ _2319;
  wire _9029 = _9026 ^ _9028;
  wire _9030 = _9024 ^ _9029;
  wire _9031 = _9019 ^ _9030;
  wire _9032 = _9010 ^ _9031;
  wire _9033 = uncoded_block[1445] ^ uncoded_block[1447];
  wire _9034 = _2321 ^ _9033;
  wire _9035 = _2325 ^ _1544;
  wire _9036 = _9034 ^ _9035;
  wire _9037 = uncoded_block[1455] ^ uncoded_block[1459];
  wire _9038 = _9037 ^ _7243;
  wire _9039 = _1550 ^ _4603;
  wire _9040 = _9038 ^ _9039;
  wire _9041 = _9036 ^ _9040;
  wire _9042 = uncoded_block[1481] ^ uncoded_block[1484];
  wire _9043 = _4604 ^ _9042;
  wire _9044 = uncoded_block[1491] ^ uncoded_block[1494];
  wire _9045 = _1563 ^ _9044;
  wire _9046 = _9043 ^ _9045;
  wire _9047 = _743 ^ _3109;
  wire _9048 = uncoded_block[1504] ^ uncoded_block[1507];
  wire _9049 = _9048 ^ _5333;
  wire _9050 = _9047 ^ _9049;
  wire _9051 = _9046 ^ _9050;
  wire _9052 = _9041 ^ _9051;
  wire _9053 = uncoded_block[1512] ^ uncoded_block[1513];
  wire _9054 = _5334 ^ _9053;
  wire _9055 = uncoded_block[1514] ^ uncoded_block[1515];
  wire _9056 = _9055 ^ _5337;
  wire _9057 = _9054 ^ _9056;
  wire _9058 = uncoded_block[1518] ^ uncoded_block[1519];
  wire _9059 = uncoded_block[1522] ^ uncoded_block[1523];
  wire _9060 = _9058 ^ _9059;
  wire _9061 = _8473 ^ _4624;
  wire _9062 = _9060 ^ _9061;
  wire _9063 = _9057 ^ _9062;
  wire _9064 = uncoded_block[1533] ^ uncoded_block[1535];
  wire _9065 = _9064 ^ _6650;
  wire _9066 = uncoded_block[1540] ^ uncoded_block[1548];
  wire _9067 = uncoded_block[1549] ^ uncoded_block[1551];
  wire _9068 = _9066 ^ _9067;
  wire _9069 = _9065 ^ _9068;
  wire _9070 = uncoded_block[1554] ^ uncoded_block[1555];
  wire _9071 = _9070 ^ _1596;
  wire _9072 = uncoded_block[1567] ^ uncoded_block[1571];
  wire _9073 = _6019 ^ _9072;
  wire _9074 = _9071 ^ _9073;
  wire _9075 = _9069 ^ _9074;
  wire _9076 = _9063 ^ _9075;
  wire _9077 = _9052 ^ _9076;
  wire _9078 = _9032 ^ _9077;
  wire _9079 = _8990 ^ _9078;
  wire _9080 = uncoded_block[1572] ^ uncoded_block[1573];
  wire _9081 = _9080 ^ _781;
  wire _9082 = uncoded_block[1577] ^ uncoded_block[1586];
  wire _9083 = uncoded_block[1588] ^ uncoded_block[1592];
  wire _9084 = _9082 ^ _9083;
  wire _9085 = _9081 ^ _9084;
  wire _9086 = uncoded_block[1595] ^ uncoded_block[1602];
  wire _9087 = _6673 ^ _9086;
  wire _9088 = uncoded_block[1604] ^ uncoded_block[1606];
  wire _9089 = uncoded_block[1607] ^ uncoded_block[1610];
  wire _9090 = _9088 ^ _9089;
  wire _9091 = _9087 ^ _9090;
  wire _9092 = _9085 ^ _9091;
  wire _9093 = _7908 ^ _6679;
  wire _9094 = uncoded_block[1617] ^ uncoded_block[1619];
  wire _9095 = uncoded_block[1620] ^ uncoded_block[1621];
  wire _9096 = _9094 ^ _9095;
  wire _9097 = _9093 ^ _9096;
  wire _9098 = _7300 ^ _1636;
  wire _9099 = uncoded_block[1633] ^ uncoded_block[1637];
  wire _9100 = _1639 ^ _9099;
  wire _9101 = _9098 ^ _9100;
  wire _9102 = _9097 ^ _9101;
  wire _9103 = _9092 ^ _9102;
  wire _9104 = _7308 ^ _6689;
  wire _9105 = uncoded_block[1645] ^ uncoded_block[1650];
  wire _9106 = uncoded_block[1652] ^ uncoded_block[1654];
  wire _9107 = _9105 ^ _9106;
  wire _9108 = _9104 ^ _9107;
  wire _9109 = _3174 ^ _3958;
  wire _9110 = _7319 ^ _2422;
  wire _9111 = _9109 ^ _9110;
  wire _9112 = _9108 ^ _9111;
  wire _9113 = uncoded_block[1680] ^ uncoded_block[1682];
  wire _9114 = _7325 ^ _9113;
  wire _9115 = uncoded_block[1690] ^ uncoded_block[1692];
  wire _9116 = _3965 ^ _9115;
  wire _9117 = _9114 ^ _9116;
  wire _9118 = uncoded_block[1695] ^ uncoded_block[1698];
  wire _9119 = _6066 ^ _9118;
  wire _9120 = uncoded_block[1699] ^ uncoded_block[1702];
  wire _9121 = _9120 ^ _847;
  wire _9122 = _9119 ^ _9121;
  wire _9123 = _9117 ^ _9122;
  wire _9124 = _9112 ^ _9123;
  wire _9125 = _9103 ^ _9124;
  wire _9126 = uncoded_block[1712] ^ uncoded_block[1714];
  wire _9127 = _848 ^ _9126;
  wire _9128 = _1677 ^ _860;
  wire _9129 = _9127 ^ _9128;
  wire _9130 = _9129 ^ uncoded_block[1722];
  wire _9131 = _9125 ^ _9130;
  wire _9132 = _9079 ^ _9131;
  wire _9133 = _8903 ^ _9132;
  wire _9134 = _3209 ^ _6080;
  wire _9135 = uncoded_block[8] ^ uncoded_block[11];
  wire _9136 = _9135 ^ _7956;
  wire _9137 = _9134 ^ _9136;
  wire _9138 = _5423 ^ _3217;
  wire _9139 = uncoded_block[21] ^ uncoded_block[25];
  wire _9140 = _9139 ^ _7959;
  wire _9141 = _9138 ^ _9140;
  wire _9142 = _9137 ^ _9141;
  wire _9143 = uncoded_block[28] ^ uncoded_block[29];
  wire _9144 = uncoded_block[30] ^ uncoded_block[33];
  wire _9145 = _9143 ^ _9144;
  wire _9146 = _3227 ^ _19;
  wire _9147 = _9145 ^ _9146;
  wire _9148 = uncoded_block[41] ^ uncoded_block[45];
  wire _9149 = _9148 ^ _8554;
  wire _9150 = uncoded_block[48] ^ uncoded_block[50];
  wire _9151 = _9150 ^ _8556;
  wire _9152 = _9149 ^ _9151;
  wire _9153 = _9147 ^ _9152;
  wire _9154 = _9142 ^ _9153;
  wire _9155 = uncoded_block[55] ^ uncoded_block[58];
  wire _9156 = uncoded_block[62] ^ uncoded_block[67];
  wire _9157 = _9155 ^ _9156;
  wire _9158 = _7367 ^ _4733;
  wire _9159 = _9157 ^ _9158;
  wire _9160 = _1712 ^ _6750;
  wire _9161 = uncoded_block[83] ^ uncoded_block[85];
  wire _9162 = _9161 ^ _42;
  wire _9163 = _9160 ^ _9162;
  wire _9164 = _9159 ^ _9163;
  wire _9165 = _6115 ^ _46;
  wire _9166 = uncoded_block[104] ^ uncoded_block[107];
  wire _9167 = _910 ^ _9166;
  wire _9168 = _9165 ^ _9167;
  wire _9169 = _2491 ^ _5453;
  wire _9170 = _6763 ^ _2495;
  wire _9171 = _9169 ^ _9170;
  wire _9172 = _9168 ^ _9171;
  wire _9173 = _9164 ^ _9172;
  wire _9174 = _9154 ^ _9173;
  wire _9175 = uncoded_block[125] ^ uncoded_block[127];
  wire _9176 = _4750 ^ _9175;
  wire _9177 = uncoded_block[133] ^ uncoded_block[134];
  wire _9178 = _8579 ^ _9177;
  wire _9179 = _9176 ^ _9178;
  wire _9180 = uncoded_block[137] ^ uncoded_block[141];
  wire _9181 = _8581 ^ _9180;
  wire _9182 = uncoded_block[145] ^ uncoded_block[148];
  wire _9183 = _9182 ^ _70;
  wire _9184 = _9181 ^ _9183;
  wire _9185 = _9179 ^ _9184;
  wire _9186 = uncoded_block[153] ^ uncoded_block[155];
  wire _9187 = _9186 ^ _1748;
  wire _9188 = uncoded_block[158] ^ uncoded_block[160];
  wire _9189 = _9188 ^ _6785;
  wire _9190 = _9187 ^ _9189;
  wire _9191 = _6147 ^ _6149;
  wire _9192 = _6789 ^ _9191;
  wire _9193 = _9190 ^ _9192;
  wire _9194 = _9185 ^ _9193;
  wire _9195 = uncoded_block[178] ^ uncoded_block[181];
  wire _9196 = uncoded_block[185] ^ uncoded_block[190];
  wire _9197 = _9195 ^ _9196;
  wire _9198 = _1763 ^ _94;
  wire _9199 = _9197 ^ _9198;
  wire _9200 = uncoded_block[198] ^ uncoded_block[202];
  wire _9201 = _9200 ^ _955;
  wire _9202 = uncoded_block[213] ^ uncoded_block[218];
  wire _9203 = _9202 ^ _102;
  wire _9204 = _9201 ^ _9203;
  wire _9205 = _9199 ^ _9204;
  wire _9206 = uncoded_block[222] ^ uncoded_block[225];
  wire _9207 = _9206 ^ _6168;
  wire _9208 = uncoded_block[235] ^ uncoded_block[237];
  wire _9209 = _8028 ^ _9208;
  wire _9210 = _9207 ^ _9209;
  wire _9211 = uncoded_block[240] ^ uncoded_block[244];
  wire _9212 = uncoded_block[246] ^ uncoded_block[249];
  wire _9213 = _9211 ^ _9212;
  wire _9214 = uncoded_block[254] ^ uncoded_block[260];
  wire _9215 = _7434 ^ _9214;
  wire _9216 = _9213 ^ _9215;
  wire _9217 = _9210 ^ _9216;
  wire _9218 = _9205 ^ _9217;
  wire _9219 = _9194 ^ _9218;
  wire _9220 = _9174 ^ _9219;
  wire _9221 = _120 ^ _1792;
  wire _9222 = uncoded_block[273] ^ uncoded_block[277];
  wire _9223 = _2566 ^ _9222;
  wire _9224 = _9221 ^ _9223;
  wire _9225 = uncoded_block[279] ^ uncoded_block[287];
  wire _9226 = uncoded_block[289] ^ uncoded_block[290];
  wire _9227 = _9225 ^ _9226;
  wire _9228 = _4819 ^ _1806;
  wire _9229 = _9227 ^ _9228;
  wire _9230 = _9224 ^ _9229;
  wire _9231 = _142 ^ _6845;
  wire _9232 = _9231 ^ _7455;
  wire _9233 = uncoded_block[313] ^ uncoded_block[317];
  wire _9234 = _9233 ^ _4832;
  wire _9235 = uncoded_block[329] ^ uncoded_block[330];
  wire _9236 = _2583 ^ _9235;
  wire _9237 = _9234 ^ _9236;
  wire _9238 = _9232 ^ _9237;
  wire _9239 = _9230 ^ _9238;
  wire _9240 = uncoded_block[331] ^ uncoded_block[333];
  wire _9241 = _9240 ^ _5536;
  wire _9242 = uncoded_block[339] ^ uncoded_block[340];
  wire _9243 = _8065 ^ _9242;
  wire _9244 = _9241 ^ _9243;
  wire _9245 = _3355 ^ _3359;
  wire _9246 = _4132 ^ _1028;
  wire _9247 = _9245 ^ _9246;
  wire _9248 = _9244 ^ _9247;
  wire _9249 = uncoded_block[355] ^ uncoded_block[358];
  wire _9250 = uncoded_block[364] ^ uncoded_block[365];
  wire _9251 = _9249 ^ _9250;
  wire _9252 = uncoded_block[369] ^ uncoded_block[375];
  wire _9253 = _9252 ^ _4854;
  wire _9254 = _9251 ^ _9253;
  wire _9255 = uncoded_block[384] ^ uncoded_block[388];
  wire _9256 = _9255 ^ _2615;
  wire _9257 = _7477 ^ _9256;
  wire _9258 = _9254 ^ _9257;
  wire _9259 = _9248 ^ _9258;
  wire _9260 = _9239 ^ _9259;
  wire _9261 = uncoded_block[394] ^ uncoded_block[398];
  wire _9262 = _3383 ^ _9261;
  wire _9263 = _4155 ^ _184;
  wire _9264 = _9262 ^ _9263;
  wire _9265 = uncoded_block[408] ^ uncoded_block[412];
  wire _9266 = uncoded_block[413] ^ uncoded_block[414];
  wire _9267 = _9265 ^ _9266;
  wire _9268 = _3396 ^ _6249;
  wire _9269 = _9267 ^ _9268;
  wire _9270 = _9264 ^ _9269;
  wire _9271 = uncoded_block[433] ^ uncoded_block[434];
  wire _9272 = _7495 ^ _9271;
  wire _9273 = _4875 ^ _9272;
  wire _9274 = _4169 ^ _5574;
  wire _9275 = uncoded_block[445] ^ uncoded_block[446];
  wire _9276 = _9275 ^ _1866;
  wire _9277 = _9274 ^ _9276;
  wire _9278 = _9273 ^ _9277;
  wire _9279 = _9270 ^ _9278;
  wire _9280 = uncoded_block[456] ^ uncoded_block[461];
  wire _9281 = uncoded_block[462] ^ uncoded_block[465];
  wire _9282 = _9280 ^ _9281;
  wire _9283 = uncoded_block[467] ^ uncoded_block[468];
  wire _9284 = _9283 ^ _4186;
  wire _9285 = _9282 ^ _9284;
  wire _9286 = _1083 ^ _2657;
  wire _9287 = uncoded_block[477] ^ uncoded_block[483];
  wire _9288 = _9287 ^ _4897;
  wire _9289 = _9286 ^ _9288;
  wire _9290 = _9285 ^ _9289;
  wire _9291 = uncoded_block[488] ^ uncoded_block[492];
  wire _9292 = uncoded_block[497] ^ uncoded_block[501];
  wire _9293 = _9291 ^ _9292;
  wire _9294 = uncoded_block[507] ^ uncoded_block[509];
  wire _9295 = uncoded_block[511] ^ uncoded_block[512];
  wire _9296 = _9294 ^ _9295;
  wire _9297 = _9293 ^ _9296;
  wire _9298 = uncoded_block[513] ^ uncoded_block[516];
  wire _9299 = uncoded_block[518] ^ uncoded_block[521];
  wire _9300 = _9298 ^ _9299;
  wire _9301 = uncoded_block[525] ^ uncoded_block[527];
  wire _9302 = _6289 ^ _9301;
  wire _9303 = _9300 ^ _9302;
  wire _9304 = _9297 ^ _9303;
  wire _9305 = _9290 ^ _9304;
  wire _9306 = _9279 ^ _9305;
  wire _9307 = _9260 ^ _9306;
  wire _9308 = _9220 ^ _9307;
  wire _9309 = uncoded_block[532] ^ uncoded_block[533];
  wire _9310 = _3447 ^ _9309;
  wire _9311 = uncoded_block[538] ^ uncoded_block[541];
  wire _9312 = _6932 ^ _9311;
  wire _9313 = _9310 ^ _9312;
  wire _9314 = uncoded_block[542] ^ uncoded_block[548];
  wire _9315 = _9314 ^ _4933;
  wire _9316 = _1122 ^ _256;
  wire _9317 = _9315 ^ _9316;
  wire _9318 = _9313 ^ _9317;
  wire _9319 = uncoded_block[561] ^ uncoded_block[562];
  wire _9320 = uncoded_block[563] ^ uncoded_block[564];
  wire _9321 = _9319 ^ _9320;
  wire _9322 = _1927 ^ _4224;
  wire _9323 = _9321 ^ _9322;
  wire _9324 = _4941 ^ _4229;
  wire _9325 = uncoded_block[582] ^ uncoded_block[583];
  wire _9326 = _9325 ^ _270;
  wire _9327 = _9324 ^ _9326;
  wire _9328 = _9323 ^ _9327;
  wire _9329 = _9318 ^ _9328;
  wire _9330 = uncoded_block[590] ^ uncoded_block[592];
  wire _9331 = _9330 ^ _2701;
  wire _9332 = uncoded_block[599] ^ uncoded_block[601];
  wire _9333 = _9332 ^ _2709;
  wire _9334 = _9331 ^ _9333;
  wire _9335 = _2710 ^ _277;
  wire _9336 = _2713 ^ _8744;
  wire _9337 = _9335 ^ _9336;
  wire _9338 = _9334 ^ _9337;
  wire _9339 = _4243 ^ _7568;
  wire _9340 = uncoded_block[624] ^ uncoded_block[629];
  wire _9341 = _9340 ^ _5661;
  wire _9342 = _9339 ^ _9341;
  wire _9343 = uncoded_block[640] ^ uncoded_block[642];
  wire _9344 = _1161 ^ _9343;
  wire _9345 = _4256 ^ _6338;
  wire _9346 = _9344 ^ _9345;
  wire _9347 = _9342 ^ _9346;
  wire _9348 = _9338 ^ _9347;
  wire _9349 = _9329 ^ _9348;
  wire _9350 = uncoded_block[649] ^ uncoded_block[651];
  wire _9351 = _9350 ^ _4975;
  wire _9352 = uncoded_block[659] ^ uncoded_block[664];
  wire _9353 = _2738 ^ _9352;
  wire _9354 = _9351 ^ _9353;
  wire _9355 = uncoded_block[665] ^ uncoded_block[668];
  wire _9356 = _9355 ^ _312;
  wire _9357 = _2748 ^ _8177;
  wire _9358 = _9356 ^ _9357;
  wire _9359 = _9354 ^ _9358;
  wire _9360 = _1971 ^ _321;
  wire _9361 = uncoded_block[686] ^ uncoded_block[691];
  wire _9362 = _9361 ^ _2755;
  wire _9363 = _9360 ^ _9362;
  wire _9364 = _4990 ^ _6364;
  wire _9365 = _2762 ^ _6366;
  wire _9366 = _9364 ^ _9365;
  wire _9367 = _9363 ^ _9366;
  wire _9368 = _9359 ^ _9367;
  wire _9369 = uncoded_block[721] ^ uncoded_block[722];
  wire _9370 = _1984 ^ _9369;
  wire _9371 = _9370 ^ _3545;
  wire _9372 = _7001 ^ _5005;
  wire _9373 = _7006 ^ _1209;
  wire _9374 = _9372 ^ _9373;
  wire _9375 = _9371 ^ _9374;
  wire _9376 = _5704 ^ _7013;
  wire _9377 = uncoded_block[756] ^ uncoded_block[760];
  wire _9378 = uncoded_block[762] ^ uncoded_block[765];
  wire _9379 = _9377 ^ _9378;
  wire _9380 = _9376 ^ _9379;
  wire _9381 = uncoded_block[767] ^ uncoded_block[771];
  wire _9382 = uncoded_block[777] ^ uncoded_block[778];
  wire _9383 = _9381 ^ _9382;
  wire _9384 = uncoded_block[779] ^ uncoded_block[782];
  wire _9385 = _9384 ^ _4309;
  wire _9386 = _9383 ^ _9385;
  wire _9387 = _9380 ^ _9386;
  wire _9388 = _9375 ^ _9387;
  wire _9389 = _9368 ^ _9388;
  wire _9390 = _9349 ^ _9389;
  wire _9391 = _371 ^ _5033;
  wire _9392 = _375 ^ _8223;
  wire _9393 = _9391 ^ _9392;
  wire _9394 = uncoded_block[803] ^ uncoded_block[806];
  wire _9395 = _4317 ^ _9394;
  wire _9396 = uncoded_block[808] ^ uncoded_block[813];
  wire _9397 = uncoded_block[814] ^ uncoded_block[817];
  wire _9398 = _9396 ^ _9397;
  wire _9399 = _9395 ^ _9398;
  wire _9400 = _9393 ^ _9399;
  wire _9401 = _7634 ^ _2032;
  wire _9402 = uncoded_block[833] ^ uncoded_block[835];
  wire _9403 = _9402 ^ _4337;
  wire _9404 = _9401 ^ _9403;
  wire _9405 = uncoded_block[842] ^ uncoded_block[847];
  wire _9406 = _5057 ^ _9405;
  wire _9407 = _2044 ^ _5742;
  wire _9408 = _9406 ^ _9407;
  wire _9409 = _9404 ^ _9408;
  wire _9410 = _9400 ^ _9409;
  wire _9411 = _5747 ^ _5069;
  wire _9412 = uncoded_block[871] ^ uncoded_block[875];
  wire _9413 = _1266 ^ _9412;
  wire _9414 = _9411 ^ _9413;
  wire _9415 = _420 ^ _7062;
  wire _9416 = uncoded_block[888] ^ uncoded_block[889];
  wire _9417 = _2058 ^ _9416;
  wire _9418 = _9415 ^ _9417;
  wire _9419 = _9414 ^ _9418;
  wire _9420 = _4355 ^ _5759;
  wire _9421 = uncoded_block[907] ^ uncoded_block[909];
  wire _9422 = _3622 ^ _9421;
  wire _9423 = _9420 ^ _9422;
  wire _9424 = uncoded_block[910] ^ uncoded_block[913];
  wire _9425 = _9424 ^ _3628;
  wire _9426 = _2076 ^ _8834;
  wire _9427 = _9425 ^ _9426;
  wire _9428 = _9423 ^ _9427;
  wire _9429 = _9419 ^ _9428;
  wire _9430 = _9410 ^ _9429;
  wire _9431 = uncoded_block[931] ^ uncoded_block[935];
  wire _9432 = _1296 ^ _9431;
  wire _9433 = uncoded_block[944] ^ uncoded_block[947];
  wire _9434 = _5101 ^ _9433;
  wire _9435 = _9432 ^ _9434;
  wire _9436 = _460 ^ _1303;
  wire _9437 = uncoded_block[954] ^ uncoded_block[957];
  wire _9438 = uncoded_block[959] ^ uncoded_block[962];
  wire _9439 = _9437 ^ _9438;
  wire _9440 = _9436 ^ _9439;
  wire _9441 = _9435 ^ _9440;
  wire _9442 = _5790 ^ _5792;
  wire _9443 = _3658 ^ _9442;
  wire _9444 = _8856 ^ _2882;
  wire _9445 = _8860 ^ _480;
  wire _9446 = _9444 ^ _9445;
  wire _9447 = _9443 ^ _9446;
  wire _9448 = _9441 ^ _9447;
  wire _9449 = uncoded_block[1000] ^ uncoded_block[1002];
  wire _9450 = _9449 ^ _2112;
  wire _9451 = uncoded_block[1011] ^ uncoded_block[1015];
  wire _9452 = _5129 ^ _9451;
  wire _9453 = _9450 ^ _9452;
  wire _9454 = uncoded_block[1022] ^ uncoded_block[1024];
  wire _9455 = uncoded_block[1025] ^ uncoded_block[1027];
  wire _9456 = _9454 ^ _9455;
  wire _9457 = _5136 ^ _9456;
  wire _9458 = _9453 ^ _9457;
  wire _9459 = uncoded_block[1029] ^ uncoded_block[1032];
  wire _9460 = _9459 ^ _2127;
  wire _9461 = uncoded_block[1035] ^ uncoded_block[1039];
  wire _9462 = _9461 ^ _6478;
  wire _9463 = _9460 ^ _9462;
  wire _9464 = uncoded_block[1050] ^ uncoded_block[1052];
  wire _9465 = uncoded_block[1054] ^ uncoded_block[1056];
  wire _9466 = _9464 ^ _9465;
  wire _9467 = _8310 ^ _9466;
  wire _9468 = _9463 ^ _9467;
  wire _9469 = _9458 ^ _9468;
  wire _9470 = _9448 ^ _9469;
  wire _9471 = _9430 ^ _9470;
  wire _9472 = _9390 ^ _9471;
  wire _9473 = _9308 ^ _9472;
  wire _9474 = _4431 ^ _4433;
  wire _9475 = uncoded_block[1066] ^ uncoded_block[1068];
  wire _9476 = _8888 ^ _9475;
  wire _9477 = _9474 ^ _9476;
  wire _9478 = uncoded_block[1075] ^ uncoded_block[1077];
  wire _9479 = _7722 ^ _9478;
  wire _9480 = uncoded_block[1082] ^ uncoded_block[1086];
  wire _9481 = _9480 ^ _1374;
  wire _9482 = _9479 ^ _9481;
  wire _9483 = _9477 ^ _9482;
  wire _9484 = uncoded_block[1104] ^ uncoded_block[1108];
  wire _9485 = _8910 ^ _9484;
  wire _9486 = _1379 ^ _9485;
  wire _9487 = uncoded_block[1113] ^ uncoded_block[1118];
  wire _9488 = _4450 ^ _9487;
  wire _9489 = uncoded_block[1119] ^ uncoded_block[1124];
  wire _9490 = _9489 ^ _5854;
  wire _9491 = _9488 ^ _9490;
  wire _9492 = _9486 ^ _9491;
  wire _9493 = _9483 ^ _9492;
  wire _9494 = uncoded_block[1130] ^ uncoded_block[1133];
  wire _9495 = _6499 ^ _9494;
  wire _9496 = uncoded_block[1136] ^ uncoded_block[1140];
  wire _9497 = _9496 ^ _568;
  wire _9498 = _9495 ^ _9497;
  wire _9499 = uncoded_block[1144] ^ uncoded_block[1148];
  wire _9500 = uncoded_block[1155] ^ uncoded_block[1157];
  wire _9501 = _9499 ^ _9500;
  wire _9502 = uncoded_block[1158] ^ uncoded_block[1164];
  wire _9503 = _9502 ^ _5193;
  wire _9504 = _9501 ^ _9503;
  wire _9505 = _9498 ^ _9504;
  wire _9506 = uncoded_block[1170] ^ uncoded_block[1172];
  wire _9507 = _9506 ^ _2967;
  wire _9508 = uncoded_block[1186] ^ uncoded_block[1188];
  wire _9509 = _2195 ^ _9508;
  wire _9510 = _9507 ^ _9509;
  wire _9511 = _2201 ^ _1420;
  wire _9512 = _6525 ^ _1421;
  wire _9513 = _9511 ^ _9512;
  wire _9514 = _9510 ^ _9513;
  wire _9515 = _9505 ^ _9514;
  wire _9516 = _9493 ^ _9515;
  wire _9517 = uncoded_block[1202] ^ uncoded_block[1208];
  wire _9518 = _9517 ^ _7765;
  wire _9519 = uncoded_block[1215] ^ uncoded_block[1222];
  wire _9520 = _3762 ^ _9519;
  wire _9521 = _9518 ^ _9520;
  wire _9522 = uncoded_block[1223] ^ uncoded_block[1228];
  wire _9523 = _9522 ^ _5218;
  wire _9524 = _2226 ^ _3772;
  wire _9525 = _9523 ^ _9524;
  wire _9526 = _9521 ^ _9525;
  wire _9527 = _6536 ^ _4509;
  wire _9528 = _4511 ^ _7778;
  wire _9529 = _9527 ^ _9528;
  wire _9530 = uncoded_block[1262] ^ uncoded_block[1265];
  wire _9531 = _1456 ^ _9530;
  wire _9532 = uncoded_block[1266] ^ uncoded_block[1268];
  wire _9533 = uncoded_block[1269] ^ uncoded_block[1271];
  wire _9534 = _9532 ^ _9533;
  wire _9535 = _9531 ^ _9534;
  wire _9536 = _9529 ^ _9535;
  wire _9537 = _9526 ^ _9536;
  wire _9538 = uncoded_block[1272] ^ uncoded_block[1273];
  wire _9539 = uncoded_block[1274] ^ uncoded_block[1277];
  wire _9540 = _9538 ^ _9539;
  wire _9541 = uncoded_block[1281] ^ uncoded_block[1283];
  wire _9542 = _631 ^ _9541;
  wire _9543 = _9540 ^ _9542;
  wire _9544 = uncoded_block[1284] ^ uncoded_block[1289];
  wire _9545 = uncoded_block[1290] ^ uncoded_block[1292];
  wire _9546 = _9544 ^ _9545;
  wire _9547 = uncoded_block[1294] ^ uncoded_block[1296];
  wire _9548 = _9547 ^ _7799;
  wire _9549 = _9546 ^ _9548;
  wire _9550 = _9543 ^ _9549;
  wire _9551 = _8984 ^ _1479;
  wire _9552 = uncoded_block[1315] ^ uncoded_block[1317];
  wire _9553 = _2261 ^ _9552;
  wire _9554 = _9551 ^ _9553;
  wire _9555 = uncoded_block[1320] ^ uncoded_block[1321];
  wire _9556 = _9555 ^ _1489;
  wire _9557 = _2268 ^ _5931;
  wire _9558 = _9556 ^ _9557;
  wire _9559 = _9554 ^ _9558;
  wire _9560 = _9550 ^ _9559;
  wire _9561 = _9537 ^ _9560;
  wire _9562 = _9516 ^ _9561;
  wire _9563 = uncoded_block[1337] ^ uncoded_block[1338];
  wire _9564 = uncoded_block[1340] ^ uncoded_block[1343];
  wire _9565 = _9563 ^ _9564;
  wire _9566 = _8417 ^ _5269;
  wire _9567 = _9565 ^ _9566;
  wire _9568 = _670 ^ _4559;
  wire _9569 = _2284 ^ _3052;
  wire _9570 = _9568 ^ _9569;
  wire _9571 = _9567 ^ _9570;
  wire _9572 = uncoded_block[1373] ^ uncoded_block[1374];
  wire _9573 = uncoded_block[1375] ^ uncoded_block[1377];
  wire _9574 = _9572 ^ _9573;
  wire _9575 = uncoded_block[1380] ^ uncoded_block[1385];
  wire _9576 = _2290 ^ _9575;
  wire _9577 = _9574 ^ _9576;
  wire _9578 = uncoded_block[1387] ^ uncoded_block[1390];
  wire _9579 = uncoded_block[1394] ^ uncoded_block[1400];
  wire _9580 = _9578 ^ _9579;
  wire _9581 = _5293 ^ _4578;
  wire _9582 = _9580 ^ _9581;
  wire _9583 = _9577 ^ _9582;
  wire _9584 = _9571 ^ _9583;
  wire _9585 = uncoded_block[1407] ^ uncoded_block[1408];
  wire _9586 = _9585 ^ _8436;
  wire _9587 = _9586 ^ _5965;
  wire _9588 = uncoded_block[1422] ^ uncoded_block[1423];
  wire _9589 = _9588 ^ _5967;
  wire _9590 = uncoded_block[1428] ^ uncoded_block[1430];
  wire _9591 = uncoded_block[1431] ^ uncoded_block[1432];
  wire _9592 = _9590 ^ _9591;
  wire _9593 = _9589 ^ _9592;
  wire _9594 = _9587 ^ _9593;
  wire _9595 = uncoded_block[1435] ^ uncoded_block[1438];
  wire _9596 = _9595 ^ _3861;
  wire _9597 = uncoded_block[1445] ^ uncoded_block[1448];
  wire _9598 = _9597 ^ _2326;
  wire _9599 = _9596 ^ _9598;
  wire _9600 = uncoded_block[1454] ^ uncoded_block[1459];
  wire _9601 = _9600 ^ _3870;
  wire _9602 = uncoded_block[1464] ^ uncoded_block[1467];
  wire _9603 = _9602 ^ _2338;
  wire _9604 = _9601 ^ _9603;
  wire _9605 = _9599 ^ _9604;
  wire _9606 = _9594 ^ _9605;
  wire _9607 = _9584 ^ _9606;
  wire _9608 = uncoded_block[1471] ^ uncoded_block[1472];
  wire _9609 = _9608 ^ _4603;
  wire _9610 = uncoded_block[1476] ^ uncoded_block[1479];
  wire _9611 = _9610 ^ _5320;
  wire _9612 = _9609 ^ _9611;
  wire _9613 = _5321 ^ _3103;
  wire _9614 = uncoded_block[1492] ^ uncoded_block[1494];
  wire _9615 = _9614 ^ _2352;
  wire _9616 = _9613 ^ _9615;
  wire _9617 = _9612 ^ _9616;
  wire _9618 = uncoded_block[1500] ^ uncoded_block[1504];
  wire _9619 = _9618 ^ _3894;
  wire _9620 = uncoded_block[1510] ^ uncoded_block[1513];
  wire _9621 = uncoded_block[1515] ^ uncoded_block[1516];
  wire _9622 = _9620 ^ _9621;
  wire _9623 = _9619 ^ _9622;
  wire _9624 = uncoded_block[1517] ^ uncoded_block[1520];
  wire _9625 = _9624 ^ _9059;
  wire _9626 = uncoded_block[1525] ^ uncoded_block[1527];
  wire _9627 = _9626 ^ _2360;
  wire _9628 = _9625 ^ _9627;
  wire _9629 = _9623 ^ _9628;
  wire _9630 = _9617 ^ _9629;
  wire _9631 = uncoded_block[1531] ^ uncoded_block[1532];
  wire _9632 = uncoded_block[1534] ^ uncoded_block[1539];
  wire _9633 = _9631 ^ _9632;
  wire _9634 = uncoded_block[1540] ^ uncoded_block[1550];
  wire _9635 = _9634 ^ _1596;
  wire _9636 = _9633 ^ _9635;
  wire _9637 = _5361 ^ _4644;
  wire _9638 = _9080 ^ _6663;
  wire _9639 = _9637 ^ _9638;
  wire _9640 = _9636 ^ _9639;
  wire _9641 = _5368 ^ _5371;
  wire _9642 = uncoded_block[1596] ^ uncoded_block[1601];
  wire _9643 = _6673 ^ _9642;
  wire _9644 = _9641 ^ _9643;
  wire _9645 = _6039 ^ _1625;
  wire _9646 = uncoded_block[1607] ^ uncoded_block[1613];
  wire _9647 = uncoded_block[1615] ^ uncoded_block[1620];
  wire _9648 = _9646 ^ _9647;
  wire _9649 = _9645 ^ _9648;
  wire _9650 = _9644 ^ _9649;
  wire _9651 = _9640 ^ _9650;
  wire _9652 = _9630 ^ _9651;
  wire _9653 = _9607 ^ _9652;
  wire _9654 = _9562 ^ _9653;
  wire _9655 = _7300 ^ _6046;
  wire _9656 = uncoded_block[1626] ^ uncoded_block[1629];
  wire _9657 = _9656 ^ _1639;
  wire _9658 = _9655 ^ _9657;
  wire _9659 = uncoded_block[1635] ^ uncoded_block[1637];
  wire _9660 = _9659 ^ _7921;
  wire _9661 = uncoded_block[1648] ^ uncoded_block[1650];
  wire _9662 = uncoded_block[1652] ^ uncoded_block[1656];
  wire _9663 = _9661 ^ _9662;
  wire _9664 = _9660 ^ _9663;
  wire _9665 = _9658 ^ _9664;
  wire _9666 = uncoded_block[1666] ^ uncoded_block[1668];
  wire _9667 = _1654 ^ _9666;
  wire _9668 = _4681 ^ _9667;
  wire _9669 = uncoded_block[1681] ^ uncoded_block[1686];
  wire _9670 = _8521 ^ _9669;
  wire _9671 = _837 ^ _7331;
  wire _9672 = _9670 ^ _9671;
  wire _9673 = _9668 ^ _9672;
  wire _9674 = _9665 ^ _9673;
  wire _9675 = uncoded_block[1692] ^ uncoded_block[1693];
  wire _9676 = _9675 ^ _840;
  wire _9677 = uncoded_block[1696] ^ uncoded_block[1697];
  wire _9678 = _9677 ^ _4700;
  wire _9679 = _9676 ^ _9678;
  wire _9680 = _2435 ^ _2437;
  wire _9681 = _9126 ^ _855;
  wire _9682 = _9680 ^ _9681;
  wire _9683 = _9679 ^ _9682;
  wire _9684 = _9683 ^ uncoded_block[1719];
  wire _9685 = _9674 ^ _9684;
  wire _9686 = _9654 ^ _9685;
  wire _9687 = _9473 ^ _9686;
  wire _9688 = uncoded_block[3] ^ uncoded_block[8];
  wire _9689 = _3209 ^ _9688;
  wire _9690 = _4 ^ _4713;
  wire _9691 = _9689 ^ _9690;
  wire _9692 = uncoded_block[16] ^ uncoded_block[18];
  wire _9693 = _9692 ^ _3217;
  wire _9694 = uncoded_block[25] ^ uncoded_block[26];
  wire _9695 = _10 ^ _9694;
  wire _9696 = _9693 ^ _9695;
  wire _9697 = _9691 ^ _9696;
  wire _9698 = _9143 ^ _875;
  wire _9699 = _9698 ^ _7963;
  wire _9700 = _882 ^ _22;
  wire _9701 = _9700 ^ _8555;
  wire _9702 = _9699 ^ _9701;
  wire _9703 = _9697 ^ _9702;
  wire _9704 = _4726 ^ _7969;
  wire _9705 = uncoded_block[65] ^ uncoded_block[66];
  wire _9706 = _9705 ^ _35;
  wire _9707 = _9704 ^ _9706;
  wire _9708 = _7976 ^ _4020;
  wire _9709 = _39 ^ _6749;
  wire _9710 = _9708 ^ _9709;
  wire _9711 = _9707 ^ _9710;
  wire _9712 = uncoded_block[82] ^ uncoded_block[87];
  wire _9713 = uncoded_block[88] ^ uncoded_block[89];
  wire _9714 = _9712 ^ _9713;
  wire _9715 = uncoded_block[92] ^ uncoded_block[94];
  wire _9716 = _903 ^ _9715;
  wire _9717 = _9714 ^ _9716;
  wire _9718 = uncoded_block[98] ^ uncoded_block[99];
  wire _9719 = _9718 ^ _4031;
  wire _9720 = uncoded_block[108] ^ uncoded_block[111];
  wire _9721 = uncoded_block[118] ^ uncoded_block[120];
  wire _9722 = _9720 ^ _9721;
  wire _9723 = _9719 ^ _9722;
  wire _9724 = _9717 ^ _9723;
  wire _9725 = _9711 ^ _9724;
  wire _9726 = _9703 ^ _9725;
  wire _9727 = uncoded_block[123] ^ uncoded_block[127];
  wire _9728 = _9727 ^ _9177;
  wire _9729 = uncoded_block[137] ^ uncoded_block[139];
  wire _9730 = uncoded_block[140] ^ uncoded_block[142];
  wire _9731 = _9729 ^ _9730;
  wire _9732 = _9728 ^ _9731;
  wire _9733 = _67 ^ _1745;
  wire _9734 = _4764 ^ _4054;
  wire _9735 = _9733 ^ _9734;
  wire _9736 = _9732 ^ _9735;
  wire _9737 = _1751 ^ _5473;
  wire _9738 = uncoded_block[174] ^ uncoded_block[179];
  wire _9739 = _938 ^ _9738;
  wire _9740 = _9737 ^ _9739;
  wire _9741 = _5480 ^ _1761;
  wire _9742 = _9740 ^ _9741;
  wire _9743 = _9736 ^ _9742;
  wire _9744 = uncoded_block[193] ^ uncoded_block[196];
  wire _9745 = uncoded_block[199] ^ uncoded_block[200];
  wire _9746 = _9744 ^ _9745;
  wire _9747 = uncoded_block[204] ^ uncoded_block[208];
  wire _9748 = _6805 ^ _9747;
  wire _9749 = _9746 ^ _9748;
  wire _9750 = uncoded_block[214] ^ uncoded_block[215];
  wire _9751 = _7415 ^ _9750;
  wire _9752 = _6812 ^ _2545;
  wire _9753 = _9751 ^ _9752;
  wire _9754 = _9749 ^ _9753;
  wire _9755 = _109 ^ _2549;
  wire _9756 = uncoded_block[240] ^ uncoded_block[241];
  wire _9757 = _9208 ^ _9756;
  wire _9758 = _9755 ^ _9757;
  wire _9759 = uncoded_block[245] ^ uncoded_block[251];
  wire _9760 = _9759 ^ _4803;
  wire _9761 = uncoded_block[254] ^ uncoded_block[255];
  wire _9762 = _9761 ^ _8041;
  wire _9763 = _9760 ^ _9762;
  wire _9764 = _9758 ^ _9763;
  wire _9765 = _9754 ^ _9764;
  wire _9766 = _9743 ^ _9765;
  wire _9767 = _9726 ^ _9766;
  wire _9768 = _977 ^ _984;
  wire _9769 = _2566 ^ _6833;
  wire _9770 = _9768 ^ _9769;
  wire _9771 = _4814 ^ _7446;
  wire _9772 = uncoded_block[287] ^ uncoded_block[289];
  wire _9773 = _8632 ^ _9772;
  wire _9774 = _9771 ^ _9773;
  wire _9775 = _9770 ^ _9774;
  wire _9776 = uncoded_block[298] ^ uncoded_block[303];
  wire _9777 = _1806 ^ _9776;
  wire _9778 = _996 ^ _9777;
  wire _9779 = uncoded_block[305] ^ uncoded_block[323];
  wire _9780 = uncoded_block[324] ^ uncoded_block[326];
  wire _9781 = _9779 ^ _9780;
  wire _9782 = uncoded_block[327] ^ uncoded_block[330];
  wire _9783 = _9782 ^ _8063;
  wire _9784 = _9781 ^ _9783;
  wire _9785 = _9778 ^ _9784;
  wire _9786 = _9775 ^ _9785;
  wire _9787 = _5536 ^ _8065;
  wire _9788 = _2595 ^ _4131;
  wire _9789 = _9787 ^ _9788;
  wire _9790 = uncoded_block[348] ^ uncoded_block[350];
  wire _9791 = _9790 ^ _1024;
  wire _9792 = _1028 ^ _8073;
  wire _9793 = _9791 ^ _9792;
  wire _9794 = _9789 ^ _9793;
  wire _9795 = _5548 ^ _8075;
  wire _9796 = _8076 ^ _6873;
  wire _9797 = _9795 ^ _9796;
  wire _9798 = uncoded_block[375] ^ uncoded_block[378];
  wire _9799 = uncoded_block[381] ^ uncoded_block[384];
  wire _9800 = _9798 ^ _9799;
  wire _9801 = _3380 ^ _2613;
  wire _9802 = _9800 ^ _9801;
  wire _9803 = _9797 ^ _9802;
  wire _9804 = _9794 ^ _9803;
  wire _9805 = _9786 ^ _9804;
  wire _9806 = uncoded_block[393] ^ uncoded_block[398];
  wire _9807 = _6239 ^ _9806;
  wire _9808 = _5559 ^ _7487;
  wire _9809 = _9807 ^ _9808;
  wire _9810 = uncoded_block[405] ^ uncoded_block[408];
  wire _9811 = _9810 ^ _4868;
  wire _9812 = uncoded_block[414] ^ uncoded_block[422];
  wire _9813 = _9812 ^ _8671;
  wire _9814 = _9811 ^ _9813;
  wire _9815 = _9809 ^ _9814;
  wire _9816 = uncoded_block[427] ^ uncoded_block[428];
  wire _9817 = _8672 ^ _9816;
  wire _9818 = _1063 ^ _6255;
  wire _9819 = _9817 ^ _9818;
  wire _9820 = uncoded_block[437] ^ uncoded_block[438];
  wire _9821 = _9820 ^ _1863;
  wire _9822 = uncoded_block[443] ^ uncoded_block[451];
  wire _9823 = _9822 ^ _1075;
  wire _9824 = _9821 ^ _9823;
  wire _9825 = _9819 ^ _9824;
  wire _9826 = _9815 ^ _9825;
  wire _9827 = uncoded_block[462] ^ uncoded_block[464];
  wire _9828 = _3415 ^ _9827;
  wire _9829 = _7509 ^ _8688;
  wire _9830 = _9828 ^ _9829;
  wire _9831 = _1086 ^ _1090;
  wire _9832 = uncoded_block[489] ^ uncoded_block[490];
  wire _9833 = _6276 ^ _9832;
  wire _9834 = _9831 ^ _9833;
  wire _9835 = _9830 ^ _9834;
  wire _9836 = _2664 ^ _8117;
  wire _9837 = uncoded_block[496] ^ uncoded_block[499];
  wire _9838 = _9837 ^ _8120;
  wire _9839 = _9836 ^ _9838;
  wire _9840 = uncoded_block[515] ^ uncoded_block[517];
  wire _9841 = uncoded_block[519] ^ uncoded_block[521];
  wire _9842 = _9840 ^ _9841;
  wire _9843 = _5612 ^ _9842;
  wire _9844 = _9839 ^ _9843;
  wire _9845 = _9835 ^ _9844;
  wire _9846 = _9826 ^ _9845;
  wire _9847 = _9805 ^ _9846;
  wire _9848 = _9767 ^ _9847;
  wire _9849 = _1898 ^ _1900;
  wire _9850 = uncoded_block[532] ^ uncoded_block[534];
  wire _9851 = _3447 ^ _9850;
  wire _9852 = _9849 ^ _9851;
  wire _9853 = uncoded_block[536] ^ uncoded_block[540];
  wire _9854 = uncoded_block[542] ^ uncoded_block[543];
  wire _9855 = _9853 ^ _9854;
  wire _9856 = _2687 ^ _3459;
  wire _9857 = _9855 ^ _9856;
  wire _9858 = _9852 ^ _9857;
  wire _9859 = _259 ^ _6945;
  wire _9860 = _4229 ^ _9325;
  wire _9861 = _9859 ^ _9860;
  wire _9862 = _8141 ^ _9861;
  wire _9863 = _9858 ^ _9862;
  wire _9864 = uncoded_block[587] ^ uncoded_block[590];
  wire _9865 = _1139 ^ _9864;
  wire _9866 = _2700 ^ _1939;
  wire _9867 = _9865 ^ _9866;
  wire _9868 = uncoded_block[602] ^ uncoded_block[604];
  wire _9869 = _1142 ^ _9868;
  wire _9870 = uncoded_block[605] ^ uncoded_block[608];
  wire _9871 = _9870 ^ _8154;
  wire _9872 = _9869 ^ _9871;
  wire _9873 = _9867 ^ _9872;
  wire _9874 = uncoded_block[618] ^ uncoded_block[625];
  wire _9875 = _9874 ^ _6966;
  wire _9876 = _6326 ^ _9875;
  wire _9877 = _289 ^ _6331;
  wire _9878 = _4255 ^ _4972;
  wire _9879 = _9877 ^ _9878;
  wire _9880 = _9876 ^ _9879;
  wire _9881 = _9873 ^ _9880;
  wire _9882 = _9863 ^ _9881;
  wire _9883 = _1957 ^ _4975;
  wire _9884 = _9883 ^ _2740;
  wire _9885 = uncoded_block[664] ^ uncoded_block[667];
  wire _9886 = uncoded_block[669] ^ uncoded_block[671];
  wire _9887 = _9885 ^ _9886;
  wire _9888 = _1178 ^ _2748;
  wire _9889 = _9887 ^ _9888;
  wire _9890 = _9884 ^ _9889;
  wire _9891 = uncoded_block[682] ^ uncoded_block[686];
  wire _9892 = _8761 ^ _9891;
  wire _9893 = _4271 ^ _325;
  wire _9894 = _9892 ^ _9893;
  wire _9895 = uncoded_block[692] ^ uncoded_block[695];
  wire _9896 = uncoded_block[696] ^ uncoded_block[700];
  wire _9897 = _9895 ^ _9896;
  wire _9898 = _334 ^ _8190;
  wire _9899 = _9897 ^ _9898;
  wire _9900 = _9894 ^ _9899;
  wire _9901 = _9890 ^ _9900;
  wire _9902 = uncoded_block[718] ^ uncoded_block[721];
  wire _9903 = _4999 ^ _9902;
  wire _9904 = uncoded_block[723] ^ uncoded_block[725];
  wire _9905 = uncoded_block[726] ^ uncoded_block[730];
  wire _9906 = _9904 ^ _9905;
  wire _9907 = _9903 ^ _9906;
  wire _9908 = uncoded_block[737] ^ uncoded_block[741];
  wire _9909 = _1203 ^ _9908;
  wire _9910 = _5702 ^ _4293;
  wire _9911 = _9909 ^ _9910;
  wire _9912 = _9907 ^ _9911;
  wire _9913 = _7013 ^ _2778;
  wire _9914 = uncoded_block[760] ^ uncoded_block[761];
  wire _9915 = _9914 ^ _9378;
  wire _9916 = _9913 ^ _9915;
  wire _9917 = uncoded_block[768] ^ uncoded_block[771];
  wire _9918 = _365 ^ _9917;
  wire _9919 = _7620 ^ _9382;
  wire _9920 = _9918 ^ _9919;
  wire _9921 = _9916 ^ _9920;
  wire _9922 = _9912 ^ _9921;
  wire _9923 = _9901 ^ _9922;
  wire _9924 = _9882 ^ _9923;
  wire _9925 = _3568 ^ _4309;
  wire _9926 = _5032 ^ _7626;
  wire _9927 = _9925 ^ _9926;
  wire _9928 = uncoded_block[798] ^ uncoded_block[802];
  wire _9929 = _382 ^ _9928;
  wire _9930 = _3577 ^ _390;
  wire _9931 = _9929 ^ _9930;
  wire _9932 = _9927 ^ _9931;
  wire _9933 = _2026 ^ _5046;
  wire _9934 = _1242 ^ _3588;
  wire _9935 = _9933 ^ _9934;
  wire _9936 = uncoded_block[831] ^ uncoded_block[835];
  wire _9937 = _5734 ^ _9936;
  wire _9938 = uncoded_block[837] ^ uncoded_block[839];
  wire _9939 = _9938 ^ _5737;
  wire _9940 = _9937 ^ _9939;
  wire _9941 = _9935 ^ _9940;
  wire _9942 = _9932 ^ _9941;
  wire _9943 = uncoded_block[845] ^ uncoded_block[851];
  wire _9944 = _1256 ^ _9943;
  wire _9945 = uncoded_block[853] ^ uncoded_block[856];
  wire _9946 = _9945 ^ _408;
  wire _9947 = _9944 ^ _9946;
  wire _9948 = uncoded_block[861] ^ uncoded_block[862];
  wire _9949 = uncoded_block[863] ^ uncoded_block[864];
  wire _9950 = _9948 ^ _9949;
  wire _9951 = _9950 ^ _5750;
  wire _9952 = _9947 ^ _9951;
  wire _9953 = uncoded_block[871] ^ uncoded_block[874];
  wire _9954 = uncoded_block[875] ^ uncoded_block[879];
  wire _9955 = _9953 ^ _9954;
  wire _9956 = uncoded_block[886] ^ uncoded_block[893];
  wire _9957 = _9956 ^ _4355;
  wire _9958 = _9955 ^ _9957;
  wire _9959 = _8250 ^ _2843;
  wire _9960 = uncoded_block[902] ^ uncoded_block[903];
  wire _9961 = uncoded_block[904] ^ uncoded_block[908];
  wire _9962 = _9960 ^ _9961;
  wire _9963 = _9959 ^ _9962;
  wire _9964 = _9958 ^ _9963;
  wire _9965 = _9952 ^ _9964;
  wire _9966 = _9942 ^ _9965;
  wire _9967 = _1287 ^ _3629;
  wire _9968 = uncoded_block[927] ^ uncoded_block[930];
  wire _9969 = _4368 ^ _9968;
  wire _9970 = _9967 ^ _9969;
  wire _9971 = uncoded_block[939] ^ uncoded_block[941];
  wire _9972 = _452 ^ _9971;
  wire _9973 = _2080 ^ _9972;
  wire _9974 = _9970 ^ _9973;
  wire _9975 = uncoded_block[947] ^ uncoded_block[948];
  wire _9976 = _455 ^ _9975;
  wire _9977 = _1303 ^ _8275;
  wire _9978 = _9976 ^ _9977;
  wire _9979 = uncoded_block[957] ^ uncoded_block[960];
  wire _9980 = _4384 ^ _9979;
  wire _9981 = uncoded_block[966] ^ uncoded_block[967];
  wire _9982 = _2872 ^ _9981;
  wire _9983 = _9980 ^ _9982;
  wire _9984 = _9978 ^ _9983;
  wire _9985 = _9974 ^ _9984;
  wire _9986 = _3657 ^ _8853;
  wire _9987 = _5113 ^ _9986;
  wire _9988 = _4397 ^ _1318;
  wire _9989 = _9988 ^ _9445;
  wire _9990 = _9987 ^ _9989;
  wire _9991 = uncoded_block[999] ^ uncoded_block[1005];
  wire _9992 = _9991 ^ _4405;
  wire _9993 = uncoded_block[1009] ^ uncoded_block[1012];
  wire _9994 = _9993 ^ _2117;
  wire _9995 = _9992 ^ _9994;
  wire _9996 = uncoded_block[1015] ^ uncoded_block[1016];
  wire _9997 = _9996 ^ _1333;
  wire _9998 = uncoded_block[1021] ^ uncoded_block[1024];
  wire _9999 = _9998 ^ _495;
  wire _10000 = _9997 ^ _9999;
  wire _10001 = _9995 ^ _10000;
  wire _10002 = _9990 ^ _10001;
  wire _10003 = _9985 ^ _10002;
  wire _10004 = _9966 ^ _10003;
  wire _10005 = _9924 ^ _10004;
  wire _10006 = _9848 ^ _10005;
  wire _10007 = _498 ^ _3675;
  wire _10008 = uncoded_block[1036] ^ uncoded_block[1041];
  wire _10009 = _10008 ^ _8309;
  wire _10010 = _10007 ^ _10009;
  wire _10011 = uncoded_block[1048] ^ uncoded_block[1053];
  wire _10012 = _10011 ^ _519;
  wire _10013 = uncoded_block[1060] ^ uncoded_block[1065];
  wire _10014 = _1363 ^ _10013;
  wire _10015 = _10012 ^ _10014;
  wire _10016 = _10010 ^ _10015;
  wire _10017 = _5158 ^ _2146;
  wire _10018 = _5162 ^ _7724;
  wire _10019 = _10017 ^ _10018;
  wire _10020 = _2928 ^ _1374;
  wire _10021 = uncoded_block[1090] ^ uncoded_block[1091];
  wire _10022 = _10021 ^ _1377;
  wire _10023 = _10020 ^ _10022;
  wire _10024 = _10019 ^ _10023;
  wire _10025 = _10016 ^ _10024;
  wire _10026 = uncoded_block[1095] ^ uncoded_block[1097];
  wire _10027 = _10026 ^ _3705;
  wire _10028 = _3707 ^ _8336;
  wire _10029 = _10027 ^ _10028;
  wire _10030 = _2165 ^ _2938;
  wire _10031 = _6496 ^ _8342;
  wire _10032 = _10030 ^ _10031;
  wire _10033 = _10029 ^ _10032;
  wire _10034 = _8343 ^ _561;
  wire _10035 = _8929 ^ _565;
  wire _10036 = _10034 ^ _10035;
  wire _10037 = _568 ^ _2953;
  wire _10038 = _5184 ^ _4466;
  wire _10039 = _10037 ^ _10038;
  wire _10040 = _10036 ^ _10039;
  wire _10041 = _10033 ^ _10040;
  wire _10042 = _10025 ^ _10041;
  wire _10043 = uncoded_block[1158] ^ uncoded_block[1161];
  wire _10044 = _8354 ^ _10043;
  wire _10045 = uncoded_block[1164] ^ uncoded_block[1167];
  wire _10046 = uncoded_block[1168] ^ uncoded_block[1170];
  wire _10047 = _10045 ^ _10046;
  wire _10048 = _10044 ^ _10047;
  wire _10049 = _8362 ^ _2967;
  wire _10050 = _2193 ^ _2195;
  wire _10051 = _10049 ^ _10050;
  wire _10052 = _10048 ^ _10051;
  wire _10053 = uncoded_block[1184] ^ uncoded_block[1187];
  wire _10054 = uncoded_block[1188] ^ uncoded_block[1197];
  wire _10055 = _10053 ^ _10054;
  wire _10056 = _2206 ^ _1425;
  wire _10057 = _10055 ^ _10056;
  wire _10058 = uncoded_block[1210] ^ uncoded_block[1215];
  wire _10059 = uncoded_block[1219] ^ uncoded_block[1221];
  wire _10060 = _10058 ^ _10059;
  wire _10061 = uncoded_block[1224] ^ uncoded_block[1227];
  wire _10062 = _7168 ^ _10061;
  wire _10063 = _10060 ^ _10062;
  wire _10064 = _10057 ^ _10063;
  wire _10065 = _10052 ^ _10064;
  wire _10066 = _1439 ^ _3771;
  wire _10067 = uncoded_block[1238] ^ uncoded_block[1241];
  wire _10068 = _10067 ^ _8963;
  wire _10069 = _10066 ^ _10068;
  wire _10070 = _2232 ^ _8385;
  wire _10071 = uncoded_block[1261] ^ uncoded_block[1266];
  wire _10072 = _8388 ^ _10071;
  wire _10073 = _10070 ^ _10072;
  wire _10074 = _10069 ^ _10073;
  wire _10075 = uncoded_block[1271] ^ uncoded_block[1274];
  wire _10076 = _10075 ^ _630;
  wire _10077 = uncoded_block[1282] ^ uncoded_block[1285];
  wire _10078 = _7183 ^ _10077;
  wire _10079 = _10076 ^ _10078;
  wire _10080 = _3798 ^ _642;
  wire _10081 = uncoded_block[1301] ^ uncoded_block[1304];
  wire _10082 = _4532 ^ _10081;
  wire _10083 = _10080 ^ _10082;
  wire _10084 = _10079 ^ _10083;
  wire _10085 = _10074 ^ _10084;
  wire _10086 = _10065 ^ _10085;
  wire _10087 = _10042 ^ _10086;
  wire _10088 = _1479 ^ _3808;
  wire _10089 = _3811 ^ _5254;
  wire _10090 = _10088 ^ _10089;
  wire _10091 = _2266 ^ _4550;
  wire _10092 = uncoded_block[1340] ^ uncoded_block[1342];
  wire _10093 = _4551 ^ _10092;
  wire _10094 = _10091 ^ _10093;
  wire _10095 = _10090 ^ _10094;
  wire _10096 = _1498 ^ _5268;
  wire _10097 = uncoded_block[1355] ^ uncoded_block[1357];
  wire _10098 = _8418 ^ _10097;
  wire _10099 = _10096 ^ _10098;
  wire _10100 = uncoded_block[1358] ^ uncoded_block[1363];
  wire _10101 = uncoded_block[1366] ^ uncoded_block[1369];
  wire _10102 = _10100 ^ _10101;
  wire _10103 = uncoded_block[1372] ^ uncoded_block[1374];
  wire _10104 = _10103 ^ _9573;
  wire _10105 = _10102 ^ _10104;
  wire _10106 = _10099 ^ _10105;
  wire _10107 = _10095 ^ _10106;
  wire _10108 = uncoded_block[1383] ^ uncoded_block[1384];
  wire _10109 = _7219 ^ _10108;
  wire _10110 = _7222 ^ _692;
  wire _10111 = _10109 ^ _10110;
  wire _10112 = _3065 ^ _6600;
  wire _10113 = uncoded_block[1407] ^ uncoded_block[1409];
  wire _10114 = _3846 ^ _10113;
  wire _10115 = _10112 ^ _10114;
  wire _10116 = _10111 ^ _10115;
  wire _10117 = uncoded_block[1410] ^ uncoded_block[1415];
  wire _10118 = uncoded_block[1416] ^ uncoded_block[1418];
  wire _10119 = _10117 ^ _10118;
  wire _10120 = uncoded_block[1419] ^ uncoded_block[1420];
  wire _10121 = _10120 ^ _7842;
  wire _10122 = _10119 ^ _10121;
  wire _10123 = _7844 ^ _9590;
  wire _10124 = uncoded_block[1433] ^ uncoded_block[1435];
  wire _10125 = _9591 ^ _10124;
  wire _10126 = _10123 ^ _10125;
  wire _10127 = _10122 ^ _10126;
  wire _10128 = _10116 ^ _10127;
  wire _10129 = _10107 ^ _10128;
  wire _10130 = uncoded_block[1440] ^ uncoded_block[1443];
  wire _10131 = _1540 ^ _10130;
  wire _10132 = uncoded_block[1452] ^ uncoded_block[1458];
  wire _10133 = _3084 ^ _10132;
  wire _10134 = _10131 ^ _10133;
  wire _10135 = _724 ^ _2336;
  wire _10136 = uncoded_block[1465] ^ uncoded_block[1467];
  wire _10137 = _10136 ^ _5983;
  wire _10138 = _10135 ^ _10137;
  wire _10139 = _10134 ^ _10138;
  wire _10140 = _5316 ^ _3884;
  wire _10141 = uncoded_block[1485] ^ uncoded_block[1495];
  wire _10142 = _9042 ^ _10141;
  wire _10143 = _10140 ^ _10142;
  wire _10144 = _7258 ^ _1572;
  wire _10145 = _7257 ^ _10144;
  wire _10146 = _10143 ^ _10145;
  wire _10147 = _10139 ^ _10146;
  wire _10148 = uncoded_block[1507] ^ uncoded_block[1514];
  wire _10149 = _10148 ^ _9621;
  wire _10150 = _9058 ^ _7269;
  wire _10151 = _10149 ^ _10150;
  wire _10152 = uncoded_block[1530] ^ uncoded_block[1534];
  wire _10153 = _9626 ^ _10152;
  wire _10154 = _6648 ^ _3908;
  wire _10155 = _10153 ^ _10154;
  wire _10156 = _10151 ^ _10155;
  wire _10157 = uncoded_block[1548] ^ uncoded_block[1552];
  wire _10158 = _10157 ^ _9070;
  wire _10159 = _3130 ^ _10158;
  wire _10160 = uncoded_block[1558] ^ uncoded_block[1561];
  wire _10161 = uncoded_block[1564] ^ uncoded_block[1567];
  wire _10162 = _10160 ^ _10161;
  wire _10163 = uncoded_block[1573] ^ uncoded_block[1578];
  wire _10164 = _7891 ^ _10163;
  wire _10165 = _10162 ^ _10164;
  wire _10166 = _10159 ^ _10165;
  wire _10167 = _10156 ^ _10166;
  wire _10168 = _10147 ^ _10167;
  wire _10169 = _10129 ^ _10168;
  wire _10170 = _10087 ^ _10169;
  wire _10171 = uncoded_block[1581] ^ uncoded_block[1585];
  wire _10172 = uncoded_block[1586] ^ uncoded_block[1589];
  wire _10173 = _10171 ^ _10172;
  wire _10174 = _4653 ^ _6673;
  wire _10175 = _10173 ^ _10174;
  wire _10176 = uncoded_block[1598] ^ uncoded_block[1604];
  wire _10177 = _10176 ^ _1625;
  wire _10178 = _5380 ^ _801;
  wire _10179 = _10177 ^ _10178;
  wire _10180 = _10175 ^ _10179;
  wire _10181 = uncoded_block[1615] ^ uncoded_block[1616];
  wire _10182 = _6042 ^ _10181;
  wire _10183 = _804 ^ _9095;
  wire _10184 = _10182 ^ _10183;
  wire _10185 = uncoded_block[1624] ^ uncoded_block[1626];
  wire _10186 = _7300 ^ _10185;
  wire _10187 = _3161 ^ _1639;
  wire _10188 = _10186 ^ _10187;
  wire _10189 = _10184 ^ _10188;
  wire _10190 = _10180 ^ _10189;
  wire _10191 = _2405 ^ _3951;
  wire _10192 = _816 ^ _1649;
  wire _10193 = _10191 ^ _10192;
  wire _10194 = uncoded_block[1651] ^ uncoded_block[1656];
  wire _10195 = _10194 ^ _1653;
  wire _10196 = uncoded_block[1660] ^ uncoded_block[1662];
  wire _10197 = _10196 ^ _3179;
  wire _10198 = _10195 ^ _10197;
  wire _10199 = _10193 ^ _10198;
  wire _10200 = uncoded_block[1666] ^ uncoded_block[1670];
  wire _10201 = _10200 ^ _2423;
  wire _10202 = uncoded_block[1679] ^ uncoded_block[1683];
  wire _10203 = _3183 ^ _10202;
  wire _10204 = _10201 ^ _10203;
  wire _10205 = uncoded_block[1687] ^ uncoded_block[1690];
  wire _10206 = _3187 ^ _10205;
  wire _10207 = _9675 ^ _3972;
  wire _10208 = _10206 ^ _10207;
  wire _10209 = _10204 ^ _10208;
  wire _10210 = _10199 ^ _10209;
  wire _10211 = _10190 ^ _10210;
  wire _10212 = uncoded_block[1697] ^ uncoded_block[1699];
  wire _10213 = _10212 ^ _3975;
  wire _10214 = uncoded_block[1707] ^ uncoded_block[1709];
  wire _10215 = _847 ^ _10214;
  wire _10216 = _10213 ^ _10215;
  wire _10217 = _2444 ^ uncoded_block[1722];
  wire _10218 = _856 ^ _10217;
  wire _10219 = _10216 ^ _10218;
  wire _10220 = _10211 ^ _10219;
  wire _10221 = _10170 ^ _10220;
  wire _10222 = _10006 ^ _10221;
  wire _10223 = uncoded_block[1] ^ uncoded_block[5];
  wire _10224 = uncoded_block[6] ^ uncoded_block[11];
  wire _10225 = _10223 ^ _10224;
  wire _10226 = uncoded_block[18] ^ uncoded_block[19];
  wire _10227 = _7956 ^ _10226;
  wire _10228 = _10225 ^ _10227;
  wire _10229 = uncoded_block[23] ^ uncoded_block[29];
  wire _10230 = _10229 ^ _3225;
  wire _10231 = _3227 ^ _882;
  wire _10232 = _10230 ^ _10231;
  wire _10233 = _10228 ^ _10232;
  wire _10234 = uncoded_block[45] ^ uncoded_block[48];
  wire _10235 = _22 ^ _10234;
  wire _10236 = _1699 ^ _4014;
  wire _10237 = _10235 ^ _10236;
  wire _10238 = uncoded_block[54] ^ uncoded_block[56];
  wire _10239 = _10238 ^ _2472;
  wire _10240 = _894 ^ _6744;
  wire _10241 = _10239 ^ _10240;
  wire _10242 = _10237 ^ _10241;
  wire _10243 = _10233 ^ _10242;
  wire _10244 = uncoded_block[73] ^ uncoded_block[75];
  wire _10245 = _3241 ^ _10244;
  wire _10246 = uncoded_block[78] ^ uncoded_block[83];
  wire _10247 = _39 ^ _10246;
  wire _10248 = _10245 ^ _10247;
  wire _10249 = uncoded_block[84] ^ uncoded_block[88];
  wire _10250 = _10249 ^ _6757;
  wire _10251 = uncoded_block[97] ^ uncoded_block[101];
  wire _10252 = uncoded_block[105] ^ uncoded_block[114];
  wire _10253 = _10251 ^ _10252;
  wire _10254 = _10250 ^ _10253;
  wire _10255 = _10248 ^ _10254;
  wire _10256 = uncoded_block[121] ^ uncoded_block[124];
  wire _10257 = _2497 ^ _10256;
  wire _10258 = _4753 ^ _4042;
  wire _10259 = _10257 ^ _10258;
  wire _10260 = _926 ^ _4760;
  wire _10261 = uncoded_block[141] ^ uncoded_block[149];
  wire _10262 = uncoded_block[150] ^ uncoded_block[152];
  wire _10263 = _10261 ^ _10262;
  wire _10264 = _10260 ^ _10263;
  wire _10265 = _10259 ^ _10264;
  wire _10266 = _10255 ^ _10265;
  wire _10267 = _10243 ^ _10266;
  wire _10268 = _4050 ^ _4055;
  wire _10269 = uncoded_block[166] ^ uncoded_block[170];
  wire _10270 = uncoded_block[172] ^ uncoded_block[176];
  wire _10271 = _10269 ^ _10270;
  wire _10272 = _940 ^ _2525;
  wire _10273 = _10271 ^ _10272;
  wire _10274 = _10268 ^ _10273;
  wire _10275 = uncoded_block[184] ^ uncoded_block[188];
  wire _10276 = _10275 ^ _6798;
  wire _10277 = uncoded_block[195] ^ uncoded_block[196];
  wire _10278 = uncoded_block[202] ^ uncoded_block[204];
  wire _10279 = _10277 ^ _10278;
  wire _10280 = _10276 ^ _10279;
  wire _10281 = _8600 ^ _7415;
  wire _10282 = uncoded_block[217] ^ uncoded_block[223];
  wire _10283 = _3296 ^ _10282;
  wire _10284 = _10281 ^ _10283;
  wire _10285 = _10280 ^ _10284;
  wire _10286 = _10274 ^ _10285;
  wire _10287 = uncoded_block[227] ^ uncoded_block[230];
  wire _10288 = _105 ^ _10287;
  wire _10289 = uncoded_block[235] ^ uncoded_block[236];
  wire _10290 = _967 ^ _10289;
  wire _10291 = _10288 ^ _10290;
  wire _10292 = uncoded_block[239] ^ uncoded_block[240];
  wire _10293 = _970 ^ _10292;
  wire _10294 = _4799 ^ _7434;
  wire _10295 = _10293 ^ _10294;
  wire _10296 = _10291 ^ _10295;
  wire _10297 = uncoded_block[259] ^ uncoded_block[262];
  wire _10298 = _2559 ^ _10297;
  wire _10299 = uncoded_block[263] ^ uncoded_block[273];
  wire _10300 = uncoded_block[274] ^ uncoded_block[276];
  wire _10301 = _10299 ^ _10300;
  wire _10302 = _10298 ^ _10301;
  wire _10303 = uncoded_block[277] ^ uncoded_block[278];
  wire _10304 = uncoded_block[280] ^ uncoded_block[282];
  wire _10305 = _10303 ^ _10304;
  wire _10306 = _6197 ^ _9226;
  wire _10307 = _10305 ^ _10306;
  wire _10308 = _10302 ^ _10307;
  wire _10309 = _10296 ^ _10308;
  wire _10310 = _10286 ^ _10309;
  wire _10311 = _10267 ^ _10310;
  wire _10312 = uncoded_block[297] ^ uncoded_block[298];
  wire _10313 = _3328 ^ _10312;
  wire _10314 = _1000 ^ _8055;
  wire _10315 = _10313 ^ _10314;
  wire _10316 = _4115 ^ _146;
  wire _10317 = _4118 ^ _1009;
  wire _10318 = _10316 ^ _10317;
  wire _10319 = _10315 ^ _10318;
  wire _10320 = _1014 ^ _2584;
  wire _10321 = _1821 ^ _6857;
  wire _10322 = _10320 ^ _10321;
  wire _10323 = uncoded_block[337] ^ uncoded_block[339];
  wire _10324 = _10323 ^ _6217;
  wire _10325 = _6859 ^ _3359;
  wire _10326 = _10324 ^ _10325;
  wire _10327 = _10322 ^ _10326;
  wire _10328 = _10319 ^ _10327;
  wire _10329 = uncoded_block[351] ^ uncoded_block[357];
  wire _10330 = _10329 ^ _6227;
  wire _10331 = uncoded_block[361] ^ uncoded_block[365];
  wire _10332 = _10331 ^ _1835;
  wire _10333 = _10330 ^ _10332;
  wire _10334 = uncoded_block[372] ^ uncoded_block[374];
  wire _10335 = uncoded_block[375] ^ uncoded_block[381];
  wire _10336 = _10334 ^ _10335;
  wire _10337 = _3377 ^ _3380;
  wire _10338 = _10336 ^ _10337;
  wire _10339 = _10333 ^ _10338;
  wire _10340 = uncoded_block[395] ^ uncoded_block[398];
  wire _10341 = uncoded_block[400] ^ uncoded_block[402];
  wire _10342 = _10340 ^ _10341;
  wire _10343 = _4153 ^ _10342;
  wire _10344 = uncoded_block[408] ^ uncoded_block[411];
  wire _10345 = _6244 ^ _10344;
  wire _10346 = _1055 ^ _6249;
  wire _10347 = _10345 ^ _10346;
  wire _10348 = _10343 ^ _10347;
  wire _10349 = _10339 ^ _10348;
  wire _10350 = _10328 ^ _10349;
  wire _10351 = _4874 ^ _4167;
  wire _10352 = uncoded_block[433] ^ uncoded_block[435];
  wire _10353 = _2638 ^ _10352;
  wire _10354 = _10351 ^ _10353;
  wire _10355 = _3405 ^ _3408;
  wire _10356 = uncoded_block[446] ^ uncoded_block[447];
  wire _10357 = _10356 ^ _4177;
  wire _10358 = _10355 ^ _10357;
  wire _10359 = _10354 ^ _10358;
  wire _10360 = _8681 ^ _4181;
  wire _10361 = _1077 ^ _10360;
  wire _10362 = uncoded_block[463] ^ uncoded_block[467];
  wire _10363 = _10362 ^ _8686;
  wire _10364 = _4189 ^ _7513;
  wire _10365 = _10363 ^ _10364;
  wire _10366 = _10361 ^ _10365;
  wire _10367 = _10359 ^ _10366;
  wire _10368 = uncoded_block[482] ^ uncoded_block[485];
  wire _10369 = _10368 ^ _224;
  wire _10370 = uncoded_block[490] ^ uncoded_block[491];
  wire _10371 = _10370 ^ _3432;
  wire _10372 = _10369 ^ _10371;
  wire _10373 = uncoded_block[498] ^ uncoded_block[502];
  wire _10374 = _6919 ^ _10373;
  wire _10375 = uncoded_block[505] ^ uncoded_block[507];
  wire _10376 = uncoded_block[508] ^ uncoded_block[509];
  wire _10377 = _10375 ^ _10376;
  wire _10378 = _10374 ^ _10377;
  wire _10379 = _10372 ^ _10378;
  wire _10380 = _8705 ^ _232;
  wire _10381 = uncoded_block[523] ^ uncoded_block[529];
  wire _10382 = _3445 ^ _10381;
  wire _10383 = _10380 ^ _10382;
  wire _10384 = uncoded_block[531] ^ uncoded_block[532];
  wire _10385 = uncoded_block[536] ^ uncoded_block[541];
  wire _10386 = _10384 ^ _10385;
  wire _10387 = _1117 ^ _8720;
  wire _10388 = _10386 ^ _10387;
  wire _10389 = _10383 ^ _10388;
  wire _10390 = _10379 ^ _10389;
  wire _10391 = _10367 ^ _10390;
  wire _10392 = _10350 ^ _10391;
  wire _10393 = _10311 ^ _10392;
  wire _10394 = _1915 ^ _6940;
  wire _10395 = uncoded_block[560] ^ uncoded_block[563];
  wire _10396 = _10395 ^ _7550;
  wire _10397 = _10394 ^ _10396;
  wire _10398 = _6942 ^ _262;
  wire _10399 = uncoded_block[575] ^ uncoded_block[577];
  wire _10400 = uncoded_block[578] ^ uncoded_block[580];
  wire _10401 = _10399 ^ _10400;
  wire _10402 = _10398 ^ _10401;
  wire _10403 = _10397 ^ _10402;
  wire _10404 = uncoded_block[581] ^ uncoded_block[585];
  wire _10405 = _10404 ^ _4233;
  wire _10406 = _9330 ^ _6316;
  wire _10407 = _10405 ^ _10406;
  wire _10408 = uncoded_block[597] ^ uncoded_block[600];
  wire _10409 = _1939 ^ _10408;
  wire _10410 = _3487 ^ _3489;
  wire _10411 = _10409 ^ _10410;
  wire _10412 = _10407 ^ _10411;
  wire _10413 = _10403 ^ _10412;
  wire _10414 = _4240 ^ _6957;
  wire _10415 = uncoded_block[617] ^ uncoded_block[623];
  wire _10416 = _8744 ^ _10415;
  wire _10417 = _10414 ^ _10416;
  wire _10418 = uncoded_block[624] ^ uncoded_block[625];
  wire _10419 = _10418 ^ _287;
  wire _10420 = uncoded_block[632] ^ uncoded_block[634];
  wire _10421 = _10420 ^ _1161;
  wire _10422 = _10419 ^ _10421;
  wire _10423 = _10417 ^ _10422;
  wire _10424 = uncoded_block[640] ^ uncoded_block[644];
  wire _10425 = uncoded_block[646] ^ uncoded_block[648];
  wire _10426 = _10424 ^ _10425;
  wire _10427 = uncoded_block[650] ^ uncoded_block[652];
  wire _10428 = _10427 ^ _304;
  wire _10429 = _10426 ^ _10428;
  wire _10430 = uncoded_block[657] ^ uncoded_block[662];
  wire _10431 = uncoded_block[665] ^ uncoded_block[669];
  wire _10432 = _10430 ^ _10431;
  wire _10433 = uncoded_block[670] ^ uncoded_block[673];
  wire _10434 = uncoded_block[675] ^ uncoded_block[676];
  wire _10435 = _10433 ^ _10434;
  wire _10436 = _10432 ^ _10435;
  wire _10437 = _10429 ^ _10436;
  wire _10438 = _10423 ^ _10437;
  wire _10439 = _10413 ^ _10438;
  wire _10440 = uncoded_block[678] ^ uncoded_block[680];
  wire _10441 = _10440 ^ _6353;
  wire _10442 = uncoded_block[685] ^ uncoded_block[688];
  wire _10443 = _10442 ^ _325;
  wire _10444 = _10441 ^ _10443;
  wire _10445 = uncoded_block[698] ^ uncoded_block[703];
  wire _10446 = _328 ^ _10445;
  wire _10447 = uncoded_block[704] ^ uncoded_block[705];
  wire _10448 = uncoded_block[707] ^ uncoded_block[708];
  wire _10449 = _10447 ^ _10448;
  wire _10450 = _10446 ^ _10449;
  wire _10451 = _10444 ^ _10450;
  wire _10452 = uncoded_block[713] ^ uncoded_block[714];
  wire _10453 = _4996 ^ _10452;
  wire _10454 = _4999 ^ _1984;
  wire _10455 = _10453 ^ _10454;
  wire _10456 = _6374 ^ _1988;
  wire _10457 = uncoded_block[727] ^ uncoded_block[728];
  wire _10458 = _10457 ^ _7603;
  wire _10459 = _10456 ^ _10458;
  wire _10460 = _10455 ^ _10459;
  wire _10461 = _10451 ^ _10460;
  wire _10462 = uncoded_block[737] ^ uncoded_block[744];
  wire _10463 = _8201 ^ _10462;
  wire _10464 = uncoded_block[745] ^ uncoded_block[748];
  wire _10465 = _10464 ^ _1210;
  wire _10466 = _10463 ^ _10465;
  wire _10467 = _5016 ^ _3556;
  wire _10468 = _10467 ^ _3560;
  wire _10469 = _10466 ^ _10468;
  wire _10470 = uncoded_block[767] ^ uncoded_block[768];
  wire _10471 = _10470 ^ _6382;
  wire _10472 = uncoded_block[780] ^ uncoded_block[786];
  wire _10473 = _2012 ^ _10472;
  wire _10474 = _10471 ^ _10473;
  wire _10475 = uncoded_block[789] ^ uncoded_block[792];
  wire _10476 = _5032 ^ _10475;
  wire _10477 = _2021 ^ _3577;
  wire _10478 = _10476 ^ _10477;
  wire _10479 = _10474 ^ _10478;
  wire _10480 = _10469 ^ _10479;
  wire _10481 = _10461 ^ _10480;
  wire _10482 = _10439 ^ _10481;
  wire _10483 = uncoded_block[811] ^ uncoded_block[812];
  wire _10484 = _5727 ^ _10483;
  wire _10485 = uncoded_block[813] ^ uncoded_block[814];
  wire _10486 = uncoded_block[816] ^ uncoded_block[820];
  wire _10487 = _10485 ^ _10486;
  wire _10488 = _10484 ^ _10487;
  wire _10489 = _7037 ^ _1246;
  wire _10490 = uncoded_block[830] ^ uncoded_block[832];
  wire _10491 = _2812 ^ _10490;
  wire _10492 = _10489 ^ _10491;
  wire _10493 = _10488 ^ _10492;
  wire _10494 = _1250 ^ _3596;
  wire _10495 = uncoded_block[842] ^ uncoded_block[845];
  wire _10496 = _5057 ^ _10495;
  wire _10497 = _10494 ^ _10496;
  wire _10498 = uncoded_block[847] ^ uncoded_block[852];
  wire _10499 = _10498 ^ _5742;
  wire _10500 = _5069 ^ _5071;
  wire _10501 = _10499 ^ _10500;
  wire _10502 = _10497 ^ _10501;
  wire _10503 = _10493 ^ _10502;
  wire _10504 = _2835 ^ _7062;
  wire _10505 = _7653 ^ _10504;
  wire _10506 = uncoded_block[889] ^ uncoded_block[892];
  wire _10507 = _5082 ^ _10506;
  wire _10508 = uncoded_block[901] ^ uncoded_block[903];
  wire _10509 = _1277 ^ _10508;
  wire _10510 = _10507 ^ _10509;
  wire _10511 = _10505 ^ _10510;
  wire _10512 = _8254 ^ _2071;
  wire _10513 = uncoded_block[916] ^ uncoded_block[919];
  wire _10514 = _10513 ^ _3632;
  wire _10515 = _10512 ^ _10514;
  wire _10516 = _8834 ^ _5096;
  wire _10517 = uncoded_block[934] ^ uncoded_block[936];
  wire _10518 = _10517 ^ _7673;
  wire _10519 = _10516 ^ _10518;
  wire _10520 = _10515 ^ _10519;
  wire _10521 = _10511 ^ _10520;
  wire _10522 = _10503 ^ _10521;
  wire _10523 = uncoded_block[941] ^ uncoded_block[944];
  wire _10524 = _10523 ^ _4381;
  wire _10525 = uncoded_block[955] ^ uncoded_block[957];
  wire _10526 = _8275 ^ _10525;
  wire _10527 = _10524 ^ _10526;
  wire _10528 = uncoded_block[958] ^ uncoded_block[960];
  wire _10529 = uncoded_block[961] ^ uncoded_block[962];
  wire _10530 = _10528 ^ _10529;
  wire _10531 = uncoded_block[964] ^ uncoded_block[966];
  wire _10532 = _10531 ^ _2093;
  wire _10533 = _10530 ^ _10532;
  wire _10534 = _10527 ^ _10533;
  wire _10535 = _5789 ^ _2100;
  wire _10536 = _3658 ^ _10535;
  wire _10537 = uncoded_block[981] ^ uncoded_block[983];
  wire _10538 = _10537 ^ _7093;
  wire _10539 = _1317 ^ _2882;
  wire _10540 = _10538 ^ _10539;
  wire _10541 = _10536 ^ _10540;
  wire _10542 = _10534 ^ _10541;
  wire _10543 = uncoded_block[993] ^ uncoded_block[994];
  wire _10544 = _10543 ^ _6457;
  wire _10545 = _9449 ^ _3666;
  wire _10546 = _10544 ^ _10545;
  wire _10547 = uncoded_block[1014] ^ uncoded_block[1018];
  wire _10548 = _2890 ^ _10547;
  wire _10549 = _2894 ^ _1334;
  wire _10550 = _10548 ^ _10549;
  wire _10551 = _10546 ^ _10550;
  wire _10552 = _8301 ^ _8874;
  wire _10553 = _2898 ^ _2907;
  wire _10554 = _10552 ^ _10553;
  wire _10555 = _7707 ^ _2129;
  wire _10556 = _5812 ^ _8309;
  wire _10557 = _10555 ^ _10556;
  wire _10558 = _10554 ^ _10557;
  wire _10559 = _10551 ^ _10558;
  wire _10560 = _10542 ^ _10559;
  wire _10561 = _10522 ^ _10560;
  wire _10562 = _10482 ^ _10561;
  wire _10563 = _10393 ^ _10562;
  wire _10564 = uncoded_block[1050] ^ uncoded_block[1054];
  wire _10565 = _2134 ^ _10564;
  wire _10566 = uncoded_block[1058] ^ uncoded_block[1060];
  wire _10567 = _519 ^ _10566;
  wire _10568 = _10565 ^ _10567;
  wire _10569 = uncoded_block[1065] ^ uncoded_block[1067];
  wire _10570 = _2917 ^ _10569;
  wire _10571 = uncoded_block[1073] ^ uncoded_block[1078];
  wire _10572 = _5156 ^ _10571;
  wire _10573 = _10570 ^ _10572;
  wire _10574 = _10568 ^ _10573;
  wire _10575 = uncoded_block[1082] ^ uncoded_block[1083];
  wire _10576 = _5834 ^ _10575;
  wire _10577 = uncoded_block[1084] ^ uncoded_block[1089];
  wire _10578 = _10577 ^ _1377;
  wire _10579 = _10576 ^ _10578;
  wire _10580 = _3698 ^ _1380;
  wire _10581 = _8910 ^ _2160;
  wire _10582 = _10580 ^ _10581;
  wire _10583 = _10579 ^ _10582;
  wire _10584 = _10574 ^ _10583;
  wire _10585 = uncoded_block[1111] ^ uncoded_block[1115];
  wire _10586 = _8915 ^ _10585;
  wire _10587 = uncoded_block[1120] ^ uncoded_block[1122];
  wire _10588 = _8920 ^ _10587;
  wire _10589 = _10586 ^ _10588;
  wire _10590 = uncoded_block[1130] ^ uncoded_block[1132];
  wire _10591 = uncoded_block[1133] ^ uncoded_block[1135];
  wire _10592 = _10590 ^ _10591;
  wire _10593 = uncoded_block[1137] ^ uncoded_block[1138];
  wire _10594 = _10593 ^ _3721;
  wire _10595 = _10592 ^ _10594;
  wire _10596 = _10589 ^ _10595;
  wire _10597 = uncoded_block[1146] ^ uncoded_block[1147];
  wire _10598 = _568 ^ _10597;
  wire _10599 = _5866 ^ _8354;
  wire _10600 = _10598 ^ _10599;
  wire _10601 = _3734 ^ _3736;
  wire _10602 = uncoded_block[1170] ^ uncoded_block[1173];
  wire _10603 = _4476 ^ _10602;
  wire _10604 = _10601 ^ _10603;
  wire _10605 = _10600 ^ _10604;
  wire _10606 = _10596 ^ _10605;
  wire _10607 = _10584 ^ _10606;
  wire _10608 = uncoded_block[1179] ^ uncoded_block[1181];
  wire _10609 = _10608 ^ _592;
  wire _10610 = _2968 ^ _10609;
  wire _10611 = _4486 ^ _3747;
  wire _10612 = uncoded_block[1191] ^ uncoded_block[1193];
  wire _10613 = _10612 ^ _6525;
  wire _10614 = _10611 ^ _10613;
  wire _10615 = _10610 ^ _10614;
  wire _10616 = _597 ^ _8370;
  wire _10617 = uncoded_block[1210] ^ uncoded_block[1212];
  wire _10618 = _2978 ^ _10617;
  wire _10619 = _10616 ^ _10618;
  wire _10620 = uncoded_block[1216] ^ uncoded_block[1218];
  wire _10621 = _3762 ^ _10620;
  wire _10622 = _608 ^ _2986;
  wire _10623 = _10621 ^ _10622;
  wire _10624 = _10619 ^ _10623;
  wire _10625 = _10615 ^ _10624;
  wire _10626 = _7169 ^ _2989;
  wire _10627 = uncoded_block[1241] ^ uncoded_block[1242];
  wire _10628 = _5221 ^ _10627;
  wire _10629 = _10626 ^ _10628;
  wire _10630 = uncoded_block[1245] ^ uncoded_block[1251];
  wire _10631 = _2995 ^ _10630;
  wire _10632 = _5231 ^ _7780;
  wire _10633 = _10631 ^ _10632;
  wire _10634 = _10629 ^ _10633;
  wire _10635 = _2239 ^ _7179;
  wire _10636 = _3005 ^ _10635;
  wire _10637 = _5905 ^ _5907;
  wire _10638 = uncoded_block[1277] ^ uncoded_block[1280];
  wire _10639 = _10638 ^ _638;
  wire _10640 = _10637 ^ _10639;
  wire _10641 = _10636 ^ _10640;
  wire _10642 = _10634 ^ _10641;
  wire _10643 = _10625 ^ _10642;
  wire _10644 = _10607 ^ _10643;
  wire _10645 = _639 ^ _9545;
  wire _10646 = uncoded_block[1293] ^ uncoded_block[1294];
  wire _10647 = uncoded_block[1295] ^ uncoded_block[1299];
  wire _10648 = _10646 ^ _10647;
  wire _10649 = _10645 ^ _10648;
  wire _10650 = uncoded_block[1300] ^ uncoded_block[1304];
  wire _10651 = _10650 ^ _3807;
  wire _10652 = _1482 ^ _3026;
  wire _10653 = _10651 ^ _10652;
  wire _10654 = _10649 ^ _10653;
  wire _10655 = uncoded_block[1327] ^ uncoded_block[1329];
  wire _10656 = _656 ^ _10655;
  wire _10657 = _7200 ^ _10656;
  wire _10658 = _8998 ^ _7815;
  wire _10659 = uncoded_block[1346] ^ uncoded_block[1349];
  wire _10660 = _1498 ^ _10659;
  wire _10661 = _10658 ^ _10660;
  wire _10662 = _10657 ^ _10661;
  wire _10663 = _10654 ^ _10662;
  wire _10664 = _8418 ^ _3045;
  wire _10665 = uncoded_block[1365] ^ uncoded_block[1366];
  wire _10666 = _1504 ^ _10665;
  wire _10667 = _10664 ^ _10666;
  wire _10668 = uncoded_block[1368] ^ uncoded_block[1369];
  wire _10669 = uncoded_block[1372] ^ uncoded_block[1376];
  wire _10670 = _10668 ^ _10669;
  wire _10671 = uncoded_block[1377] ^ uncoded_block[1383];
  wire _10672 = _10671 ^ _6596;
  wire _10673 = _10670 ^ _10672;
  wire _10674 = _10667 ^ _10673;
  wire _10675 = uncoded_block[1387] ^ uncoded_block[1395];
  wire _10676 = uncoded_block[1396] ^ uncoded_block[1399];
  wire _10677 = _10675 ^ _10676;
  wire _10678 = uncoded_block[1403] ^ uncoded_block[1408];
  wire _10679 = _10678 ^ _7229;
  wire _10680 = _10677 ^ _10679;
  wire _10681 = uncoded_block[1413] ^ uncoded_block[1416];
  wire _10682 = _10681 ^ _5964;
  wire _10683 = uncoded_block[1422] ^ uncoded_block[1425];
  wire _10684 = uncoded_block[1428] ^ uncoded_block[1429];
  wire _10685 = _10683 ^ _10684;
  wire _10686 = _10682 ^ _10685;
  wire _10687 = _10680 ^ _10686;
  wire _10688 = _10674 ^ _10687;
  wire _10689 = _10663 ^ _10688;
  wire _10690 = uncoded_block[1433] ^ uncoded_block[1437];
  wire _10691 = _1531 ^ _10690;
  wire _10692 = _2318 ^ _8449;
  wire _10693 = _10691 ^ _10692;
  wire _10694 = uncoded_block[1446] ^ uncoded_block[1450];
  wire _10695 = _10694 ^ _2326;
  wire _10696 = _6622 ^ _3088;
  wire _10697 = _10695 ^ _10696;
  wire _10698 = _10693 ^ _10697;
  wire _10699 = uncoded_block[1463] ^ uncoded_block[1465];
  wire _10700 = _726 ^ _10699;
  wire _10701 = uncoded_block[1472] ^ uncoded_block[1476];
  wire _10702 = _732 ^ _10701;
  wire _10703 = _10700 ^ _10702;
  wire _10704 = uncoded_block[1477] ^ uncoded_block[1480];
  wire _10705 = _10704 ^ _9042;
  wire _10706 = uncoded_block[1485] ^ uncoded_block[1486];
  wire _10707 = uncoded_block[1487] ^ uncoded_block[1491];
  wire _10708 = _10706 ^ _10707;
  wire _10709 = _10705 ^ _10708;
  wire _10710 = _10703 ^ _10709;
  wire _10711 = _10698 ^ _10710;
  wire _10712 = uncoded_block[1496] ^ uncoded_block[1499];
  wire _10713 = _10712 ^ _1571;
  wire _10714 = _10713 ^ _3895;
  wire _10715 = uncoded_block[1508] ^ uncoded_block[1513];
  wire _10716 = _10715 ^ _6643;
  wire _10717 = _2357 ^ _9059;
  wire _10718 = _10716 ^ _10717;
  wire _10719 = _10714 ^ _10718;
  wire _10720 = _8473 ^ _5343;
  wire _10721 = _9631 ^ _5347;
  wire _10722 = _10720 ^ _10721;
  wire _10723 = _3906 ^ _3129;
  wire _10724 = uncoded_block[1549] ^ uncoded_block[1554];
  wire _10725 = _2367 ^ _10724;
  wire _10726 = _10723 ^ _10725;
  wire _10727 = _10722 ^ _10726;
  wire _10728 = _10719 ^ _10727;
  wire _10729 = _10711 ^ _10728;
  wire _10730 = _10689 ^ _10729;
  wire _10731 = _10644 ^ _10730;
  wire _10732 = uncoded_block[1555] ^ uncoded_block[1559];
  wire _10733 = _10732 ^ _1605;
  wire _10734 = uncoded_block[1575] ^ uncoded_block[1579];
  wire _10735 = _4645 ^ _10734;
  wire _10736 = _10733 ^ _10735;
  wire _10737 = uncoded_block[1586] ^ uncoded_block[1600];
  wire _10738 = _6031 ^ _10737;
  wire _10739 = _3151 ^ _8502;
  wire _10740 = _10738 ^ _10739;
  wire _10741 = _10736 ^ _10740;
  wire _10742 = uncoded_block[1605] ^ uncoded_block[1607];
  wire _10743 = uncoded_block[1608] ^ uncoded_block[1614];
  wire _10744 = _10742 ^ _10743;
  wire _10745 = uncoded_block[1615] ^ uncoded_block[1617];
  wire _10746 = _10745 ^ _7911;
  wire _10747 = _10744 ^ _10746;
  wire _10748 = _7300 ^ _4665;
  wire _10749 = uncoded_block[1628] ^ uncoded_block[1632];
  wire _10750 = _10749 ^ _3946;
  wire _10751 = _10748 ^ _10750;
  wire _10752 = _10747 ^ _10751;
  wire _10753 = _10741 ^ _10752;
  wire _10754 = uncoded_block[1636] ^ uncoded_block[1637];
  wire _10755 = uncoded_block[1640] ^ uncoded_block[1645];
  wire _10756 = _10754 ^ _10755;
  wire _10757 = uncoded_block[1649] ^ uncoded_block[1650];
  wire _10758 = _10757 ^ _4678;
  wire _10759 = _10756 ^ _10758;
  wire _10760 = uncoded_block[1655] ^ uncoded_block[1656];
  wire _10761 = uncoded_block[1657] ^ uncoded_block[1660];
  wire _10762 = _10760 ^ _10761;
  wire _10763 = _2420 ^ _7322;
  wire _10764 = _10762 ^ _10763;
  wire _10765 = _10759 ^ _10764;
  wire _10766 = uncoded_block[1680] ^ uncoded_block[1681];
  wire _10767 = _832 ^ _10766;
  wire _10768 = uncoded_block[1687] ^ uncoded_block[1691];
  wire _10769 = _4693 ^ _10768;
  wire _10770 = _10767 ^ _10769;
  wire _10771 = uncoded_block[1694] ^ uncoded_block[1696];
  wire _10772 = _9675 ^ _10771;
  wire _10773 = _5409 ^ _6068;
  wire _10774 = _10772 ^ _10773;
  wire _10775 = _10770 ^ _10774;
  wire _10776 = _10765 ^ _10775;
  wire _10777 = _10753 ^ _10776;
  wire _10778 = uncoded_block[1709] ^ uncoded_block[1711];
  wire _10779 = _3976 ^ _10778;
  wire _10780 = _852 ^ _854;
  wire _10781 = _10779 ^ _10780;
  wire _10782 = _9128 ^ uncoded_block[1721];
  wire _10783 = _10781 ^ _10782;
  wire _10784 = _10777 ^ _10783;
  wire _10785 = _10731 ^ _10784;
  wire _10786 = _10563 ^ _10785;
  wire _10787 = uncoded_block[0] ^ uncoded_block[5];
  wire _10788 = _10787 ^ _6724;
  wire _10789 = _4 ^ _7;
  wire _10790 = _10788 ^ _10789;
  wire _10791 = uncoded_block[21] ^ uncoded_block[23];
  wire _10792 = uncoded_block[24] ^ uncoded_block[33];
  wire _10793 = _10791 ^ _10792;
  wire _10794 = _9693 ^ _10793;
  wire _10795 = _10790 ^ _10794;
  wire _10796 = uncoded_block[37] ^ uncoded_block[40];
  wire _10797 = _3227 ^ _10796;
  wire _10798 = _4008 ^ _23;
  wire _10799 = _10797 ^ _10798;
  wire _10800 = _1699 ^ _886;
  wire _10801 = uncoded_block[59] ^ uncoded_block[62];
  wire _10802 = _5436 ^ _10801;
  wire _10803 = _10800 ^ _10802;
  wire _10804 = _10799 ^ _10803;
  wire _10805 = _10795 ^ _10804;
  wire _10806 = uncoded_block[63] ^ uncoded_block[64];
  wire _10807 = _10806 ^ _6744;
  wire _10808 = _7367 ^ _1711;
  wire _10809 = _10807 ^ _10808;
  wire _10810 = _900 ^ _6750;
  wire _10811 = _9161 ^ _46;
  wire _10812 = _10810 ^ _10811;
  wire _10813 = _10809 ^ _10812;
  wire _10814 = uncoded_block[102] ^ uncoded_block[110];
  wire _10815 = _10251 ^ _10814;
  wire _10816 = uncoded_block[114] ^ uncoded_block[115];
  wire _10817 = _6126 ^ _10816;
  wire _10818 = _10815 ^ _10817;
  wire _10819 = uncoded_block[120] ^ uncoded_block[122];
  wire _10820 = _6128 ^ _10819;
  wire _10821 = uncoded_block[123] ^ uncoded_block[124];
  wire _10822 = uncoded_block[125] ^ uncoded_block[129];
  wire _10823 = _10821 ^ _10822;
  wire _10824 = _10820 ^ _10823;
  wire _10825 = _10818 ^ _10824;
  wire _10826 = _10813 ^ _10825;
  wire _10827 = _10805 ^ _10826;
  wire _10828 = uncoded_block[130] ^ uncoded_block[136];
  wire _10829 = _10828 ^ _4760;
  wire _10830 = uncoded_block[141] ^ uncoded_block[143];
  wire _10831 = _3265 ^ _10830;
  wire _10832 = _10829 ^ _10831;
  wire _10833 = _7392 ^ _6780;
  wire _10834 = uncoded_block[155] ^ uncoded_block[159];
  wire _10835 = _5469 ^ _10834;
  wire _10836 = _10833 ^ _10835;
  wire _10837 = _10832 ^ _10836;
  wire _10838 = _74 ^ _2516;
  wire _10839 = _79 ^ _5473;
  wire _10840 = _10838 ^ _10839;
  wire _10841 = uncoded_block[171] ^ uncoded_block[175];
  wire _10842 = _10841 ^ _940;
  wire _10843 = uncoded_block[182] ^ uncoded_block[184];
  wire _10844 = _5477 ^ _10843;
  wire _10845 = _10842 ^ _10844;
  wire _10846 = _10840 ^ _10845;
  wire _10847 = _10837 ^ _10846;
  wire _10848 = _5483 ^ _6801;
  wire _10849 = uncoded_block[200] ^ uncoded_block[201];
  wire _10850 = _10849 ^ _4070;
  wire _10851 = _10848 ^ _10850;
  wire _10852 = uncoded_block[206] ^ uncoded_block[209];
  wire _10853 = _10852 ^ _3292;
  wire _10854 = uncoded_block[220] ^ uncoded_block[224];
  wire _10855 = _101 ^ _10854;
  wire _10856 = _10853 ^ _10855;
  wire _10857 = _10851 ^ _10856;
  wire _10858 = _3299 ^ _109;
  wire _10859 = uncoded_block[231] ^ uncoded_block[239];
  wire _10860 = uncoded_block[242] ^ uncoded_block[243];
  wire _10861 = _10859 ^ _10860;
  wire _10862 = _10858 ^ _10861;
  wire _10863 = _5505 ^ _3309;
  wire _10864 = uncoded_block[256] ^ uncoded_block[261];
  wire _10865 = _10864 ^ _4096;
  wire _10866 = _10863 ^ _10865;
  wire _10867 = _10862 ^ _10866;
  wire _10868 = _10857 ^ _10867;
  wire _10869 = _10847 ^ _10868;
  wire _10870 = _10827 ^ _10869;
  wire _10871 = _985 ^ _2566;
  wire _10872 = uncoded_block[272] ^ uncoded_block[273];
  wire _10873 = _10872 ^ _6833;
  wire _10874 = _10871 ^ _10873;
  wire _10875 = _4814 ^ _4817;
  wire _10876 = uncoded_block[290] ^ uncoded_block[291];
  wire _10877 = _7448 ^ _10876;
  wire _10878 = _10875 ^ _10877;
  wire _10879 = _10874 ^ _10878;
  wire _10880 = uncoded_block[296] ^ uncoded_block[300];
  wire _10881 = _4820 ^ _10880;
  wire _10882 = _142 ^ _8052;
  wire _10883 = _10881 ^ _10882;
  wire _10884 = _8057 ^ _4831;
  wire _10885 = _10883 ^ _10884;
  wire _10886 = _10879 ^ _10885;
  wire _10887 = uncoded_block[325] ^ uncoded_block[330];
  wire _10888 = _5530 ^ _10887;
  wire _10889 = _8063 ^ _8646;
  wire _10890 = _10888 ^ _10889;
  wire _10891 = _2593 ^ _4844;
  wire _10892 = _3359 ^ _162;
  wire _10893 = _10891 ^ _10892;
  wire _10894 = _10890 ^ _10893;
  wire _10895 = uncoded_block[373] ^ uncoded_block[374];
  wire _10896 = _1838 ^ _10895;
  wire _10897 = _3363 ^ _10896;
  wire _10898 = uncoded_block[375] ^ uncoded_block[377];
  wire _10899 = uncoded_block[378] ^ uncoded_block[379];
  wire _10900 = _10898 ^ _10899;
  wire _10901 = uncoded_block[382] ^ uncoded_block[385];
  wire _10902 = _1841 ^ _10901;
  wire _10903 = _10900 ^ _10902;
  wire _10904 = _10897 ^ _10903;
  wire _10905 = _10894 ^ _10904;
  wire _10906 = _10886 ^ _10905;
  wire _10907 = uncoded_block[387] ^ uncoded_block[389];
  wire _10908 = uncoded_block[391] ^ uncoded_block[394];
  wire _10909 = _10907 ^ _10908;
  wire _10910 = uncoded_block[396] ^ uncoded_block[397];
  wire _10911 = uncoded_block[398] ^ uncoded_block[402];
  wire _10912 = _10910 ^ _10911;
  wire _10913 = _10909 ^ _10912;
  wire _10914 = uncoded_block[406] ^ uncoded_block[417];
  wire _10915 = _6244 ^ _10914;
  wire _10916 = _194 ^ _1062;
  wire _10917 = _10915 ^ _10916;
  wire _10918 = _10913 ^ _10917;
  wire _10919 = uncoded_block[434] ^ uncoded_block[436];
  wire _10920 = _2638 ^ _10919;
  wire _10921 = uncoded_block[442] ^ uncoded_block[449];
  wire _10922 = _5574 ^ _10921;
  wire _10923 = _10920 ^ _10922;
  wire _10924 = uncoded_block[452] ^ uncoded_block[458];
  wire _10925 = _4883 ^ _10924;
  wire _10926 = uncoded_block[459] ^ uncoded_block[461];
  wire _10927 = uncoded_block[463] ^ uncoded_block[468];
  wire _10928 = _10926 ^ _10927;
  wire _10929 = _10925 ^ _10928;
  wire _10930 = _10923 ^ _10929;
  wire _10931 = _10918 ^ _10930;
  wire _10932 = uncoded_block[473] ^ uncoded_block[479];
  wire _10933 = _8686 ^ _10932;
  wire _10934 = uncoded_block[483] ^ uncoded_block[487];
  wire _10935 = _5593 ^ _10934;
  wire _10936 = _10933 ^ _10935;
  wire _10937 = uncoded_block[492] ^ uncoded_block[494];
  wire _10938 = _7516 ^ _10937;
  wire _10939 = _5603 ^ _4905;
  wire _10940 = _10938 ^ _10939;
  wire _10941 = _10936 ^ _10940;
  wire _10942 = _6279 ^ _10375;
  wire _10943 = _3437 ^ _9295;
  wire _10944 = _10942 ^ _10943;
  wire _10945 = uncoded_block[513] ^ uncoded_block[515];
  wire _10946 = _10945 ^ _236;
  wire _10947 = uncoded_block[520] ^ uncoded_block[522];
  wire _10948 = uncoded_block[523] ^ uncoded_block[526];
  wire _10949 = _10947 ^ _10948;
  wire _10950 = _10946 ^ _10949;
  wire _10951 = _10944 ^ _10950;
  wire _10952 = _10941 ^ _10951;
  wire _10953 = _10931 ^ _10952;
  wire _10954 = _10906 ^ _10953;
  wire _10955 = _10870 ^ _10954;
  wire _10956 = _4922 ^ _1901;
  wire _10957 = _243 ^ _4217;
  wire _10958 = _10956 ^ _10957;
  wire _10959 = uncoded_block[544] ^ uncoded_block[547];
  wire _10960 = _8132 ^ _10959;
  wire _10961 = uncoded_block[548] ^ uncoded_block[551];
  wire _10962 = _10961 ^ _8724;
  wire _10963 = _10960 ^ _10962;
  wire _10964 = _10958 ^ _10963;
  wire _10965 = _8139 ^ _1925;
  wire _10966 = _10965 ^ _4225;
  wire _10967 = uncoded_block[576] ^ uncoded_block[580];
  wire _10968 = _10967 ^ _4946;
  wire _10969 = uncoded_block[585] ^ uncoded_block[591];
  wire _10970 = _10969 ^ _1938;
  wire _10971 = _10968 ^ _10970;
  wire _10972 = _10966 ^ _10971;
  wire _10973 = _10964 ^ _10972;
  wire _10974 = _2701 ^ _3486;
  wire _10975 = uncoded_block[600] ^ uncoded_block[607];
  wire _10976 = _10975 ^ _6323;
  wire _10977 = _10974 ^ _10976;
  wire _10978 = _2715 ^ _1946;
  wire _10979 = uncoded_block[622] ^ uncoded_block[626];
  wire _10980 = uncoded_block[627] ^ uncoded_block[633];
  wire _10981 = _10979 ^ _10980;
  wire _10982 = _10978 ^ _10981;
  wire _10983 = _10977 ^ _10982;
  wire _10984 = uncoded_block[635] ^ uncoded_block[641];
  wire _10985 = uncoded_block[642] ^ uncoded_block[648];
  wire _10986 = _10984 ^ _10985;
  wire _10987 = uncoded_block[654] ^ uncoded_block[656];
  wire _10988 = _9350 ^ _10987;
  wire _10989 = _10986 ^ _10988;
  wire _10990 = uncoded_block[667] ^ uncoded_block[668];
  wire _10991 = _1173 ^ _10990;
  wire _10992 = _3515 ^ _10991;
  wire _10993 = _10989 ^ _10992;
  wire _10994 = _10983 ^ _10993;
  wire _10995 = _10973 ^ _10994;
  wire _10996 = _10433 ^ _1180;
  wire _10997 = uncoded_block[682] ^ uncoded_block[687];
  wire _10998 = _8179 ^ _10997;
  wire _10999 = _10996 ^ _10998;
  wire _11000 = _4987 ^ _333;
  wire _11001 = _6361 ^ _4995;
  wire _11002 = _11000 ^ _11001;
  wire _11003 = _10999 ^ _11002;
  wire _11004 = uncoded_block[710] ^ uncoded_block[716];
  wire _11005 = _11004 ^ _1984;
  wire _11006 = uncoded_block[728] ^ uncoded_block[731];
  wire _11007 = _9904 ^ _11006;
  wire _11008 = _11005 ^ _11007;
  wire _11009 = uncoded_block[736] ^ uncoded_block[741];
  wire _11010 = _7002 ^ _11009;
  wire _11011 = uncoded_block[747] ^ uncoded_block[753];
  wire _11012 = uncoded_block[754] ^ uncoded_block[756];
  wire _11013 = _11011 ^ _11012;
  wire _11014 = _11010 ^ _11013;
  wire _11015 = _11008 ^ _11014;
  wire _11016 = _11003 ^ _11015;
  wire _11017 = _3559 ^ _2006;
  wire _11018 = uncoded_block[765] ^ uncoded_block[767];
  wire _11019 = uncoded_block[770] ^ uncoded_block[771];
  wire _11020 = _11018 ^ _11019;
  wire _11021 = _11017 ^ _11020;
  wire _11022 = uncoded_block[775] ^ uncoded_block[779];
  wire _11023 = _11022 ^ _1225;
  wire _11024 = uncoded_block[793] ^ uncoded_block[795];
  wire _11025 = _11024 ^ _8223;
  wire _11026 = _11023 ^ _11025;
  wire _11027 = _11021 ^ _11026;
  wire _11028 = _7029 ^ _5041;
  wire _11029 = uncoded_block[810] ^ uncoded_block[813];
  wire _11030 = uncoded_block[814] ^ uncoded_block[816];
  wire _11031 = _11029 ^ _11030;
  wire _11032 = _11028 ^ _11031;
  wire _11033 = _2028 ^ _7037;
  wire _11034 = uncoded_block[823] ^ uncoded_block[825];
  wire _11035 = _11034 ^ _6401;
  wire _11036 = _11033 ^ _11035;
  wire _11037 = _11032 ^ _11036;
  wire _11038 = _11027 ^ _11037;
  wire _11039 = _11016 ^ _11038;
  wire _11040 = _10995 ^ _11039;
  wire _11041 = _1249 ^ _4331;
  wire _11042 = uncoded_block[834] ^ uncoded_block[838];
  wire _11043 = uncoded_block[839] ^ uncoded_block[840];
  wire _11044 = _11042 ^ _11043;
  wire _11045 = _11041 ^ _11044;
  wire _11046 = uncoded_block[843] ^ uncoded_block[847];
  wire _11047 = _2036 ^ _11046;
  wire _11048 = uncoded_block[852] ^ uncoded_block[854];
  wire _11049 = _4340 ^ _11048;
  wire _11050 = _11047 ^ _11049;
  wire _11051 = _11045 ^ _11050;
  wire _11052 = uncoded_block[858] ^ uncoded_block[864];
  wire _11053 = uncoded_block[866] ^ uncoded_block[871];
  wire _11054 = _11052 ^ _11053;
  wire _11055 = uncoded_block[875] ^ uncoded_block[881];
  wire _11056 = uncoded_block[882] ^ uncoded_block[885];
  wire _11057 = _11055 ^ _11056;
  wire _11058 = _11054 ^ _11057;
  wire _11059 = uncoded_block[886] ^ uncoded_block[887];
  wire _11060 = uncoded_block[890] ^ uncoded_block[893];
  wire _11061 = _11059 ^ _11060;
  wire _11062 = uncoded_block[901] ^ uncoded_block[904];
  wire _11063 = _4358 ^ _11062;
  wire _11064 = _11061 ^ _11063;
  wire _11065 = _11058 ^ _11064;
  wire _11066 = _11051 ^ _11065;
  wire _11067 = uncoded_block[907] ^ uncoded_block[910];
  wire _11068 = _11067 ^ _1287;
  wire _11069 = _2852 ^ _3631;
  wire _11070 = _11068 ^ _11069;
  wire _11071 = uncoded_block[921] ^ uncoded_block[926];
  wire _11072 = _11071 ^ _7075;
  wire _11073 = _5096 ^ _5101;
  wire _11074 = _11072 ^ _11073;
  wire _11075 = _11070 ^ _11074;
  wire _11076 = uncoded_block[938] ^ uncoded_block[941];
  wire _11077 = _11076 ^ _2865;
  wire _11078 = _2086 ^ _9975;
  wire _11079 = _11077 ^ _11078;
  wire _11080 = _4381 ^ _5779;
  wire _11081 = _2869 ^ _7680;
  wire _11082 = _11080 ^ _11081;
  wire _11083 = _11079 ^ _11082;
  wire _11084 = _11075 ^ _11083;
  wire _11085 = _11066 ^ _11084;
  wire _11086 = uncoded_block[962] ^ uncoded_block[965];
  wire _11087 = uncoded_block[966] ^ uncoded_block[968];
  wire _11088 = _11086 ^ _11087;
  wire _11089 = _468 ^ _5112;
  wire _11090 = _11088 ^ _11089;
  wire _11091 = uncoded_block[975] ^ uncoded_block[977];
  wire _11092 = uncoded_block[978] ^ uncoded_block[979];
  wire _11093 = _11091 ^ _11092;
  wire _11094 = uncoded_block[980] ^ uncoded_block[982];
  wire _11095 = _11094 ^ _7093;
  wire _11096 = _11093 ^ _11095;
  wire _11097 = _11090 ^ _11096;
  wire _11098 = uncoded_block[986] ^ uncoded_block[989];
  wire _11099 = uncoded_block[991] ^ uncoded_block[995];
  wire _11100 = _11098 ^ _11099;
  wire _11101 = uncoded_block[997] ^ uncoded_block[998];
  wire _11102 = _11101 ^ _2107;
  wire _11103 = _11100 ^ _11102;
  wire _11104 = uncoded_block[1007] ^ uncoded_block[1013];
  wire _11105 = _1326 ^ _11104;
  wire _11106 = _7107 ^ _8871;
  wire _11107 = _11105 ^ _11106;
  wire _11108 = _11103 ^ _11107;
  wire _11109 = _11097 ^ _11108;
  wire _11110 = uncoded_block[1024] ^ uncoded_block[1032];
  wire _11111 = _5137 ^ _11110;
  wire _11112 = _6474 ^ _1345;
  wire _11113 = _11111 ^ _11112;
  wire _11114 = uncoded_block[1043] ^ uncoded_block[1047];
  wire _11115 = _6478 ^ _11114;
  wire _11116 = uncoded_block[1052] ^ uncoded_block[1054];
  wire _11117 = _11116 ^ _8311;
  wire _11118 = _11115 ^ _11117;
  wire _11119 = _11113 ^ _11118;
  wire _11120 = uncoded_block[1057] ^ uncoded_block[1060];
  wire _11121 = _11120 ^ _3685;
  wire _11122 = uncoded_block[1068] ^ uncoded_block[1069];
  wire _11123 = _11122 ^ _8892;
  wire _11124 = _11121 ^ _11123;
  wire _11125 = uncoded_block[1072] ^ uncoded_block[1076];
  wire _11126 = uncoded_block[1079] ^ uncoded_block[1081];
  wire _11127 = _11125 ^ _11126;
  wire _11128 = uncoded_block[1082] ^ uncoded_block[1089];
  wire _11129 = _11128 ^ _10021;
  wire _11130 = _11127 ^ _11129;
  wire _11131 = _11124 ^ _11130;
  wire _11132 = _11119 ^ _11131;
  wire _11133 = _11109 ^ _11132;
  wire _11134 = _11085 ^ _11133;
  wire _11135 = _11040 ^ _11134;
  wire _11136 = _10955 ^ _11135;
  wire _11137 = uncoded_block[1092] ^ uncoded_block[1094];
  wire _11138 = _11137 ^ _542;
  wire _11139 = uncoded_block[1097] ^ uncoded_block[1098];
  wire _11140 = _11139 ^ _5169;
  wire _11141 = _11138 ^ _11140;
  wire _11142 = uncoded_block[1102] ^ uncoded_block[1103];
  wire _11143 = _11142 ^ _3707;
  wire _11144 = _3708 ^ _2938;
  wire _11145 = _11143 ^ _11144;
  wire _11146 = _11141 ^ _11145;
  wire _11147 = uncoded_block[1117] ^ uncoded_block[1119];
  wire _11148 = _11147 ^ _1389;
  wire _11149 = _4459 ^ _560;
  wire _11150 = _11148 ^ _11149;
  wire _11151 = _561 ^ _565;
  wire _11152 = _567 ^ _5861;
  wire _11153 = _11151 ^ _11152;
  wire _11154 = _11150 ^ _11153;
  wire _11155 = _11146 ^ _11154;
  wire _11156 = _5862 ^ _4468;
  wire _11157 = uncoded_block[1155] ^ uncoded_block[1158];
  wire _11158 = _11157 ^ _582;
  wire _11159 = _11156 ^ _11158;
  wire _11160 = uncoded_block[1168] ^ uncoded_block[1169];
  wire _11161 = uncoded_block[1170] ^ uncoded_block[1171];
  wire _11162 = _11160 ^ _11161;
  wire _11163 = uncoded_block[1172] ^ uncoded_block[1180];
  wire _11164 = _11163 ^ _1417;
  wire _11165 = _11162 ^ _11164;
  wire _11166 = _11159 ^ _11165;
  wire _11167 = _4486 ^ _9508;
  wire _11168 = _6525 ^ _599;
  wire _11169 = _11167 ^ _11168;
  wire _11170 = _2974 ^ _2978;
  wire _11171 = uncoded_block[1207] ^ uncoded_block[1209];
  wire _11172 = _11171 ^ _2981;
  wire _11173 = _11170 ^ _11172;
  wire _11174 = _11169 ^ _11173;
  wire _11175 = _11166 ^ _11174;
  wire _11176 = _11155 ^ _11175;
  wire _11177 = uncoded_block[1225] ^ uncoded_block[1226];
  wire _11178 = _4502 ^ _11177;
  wire _11179 = _4500 ^ _11178;
  wire _11180 = uncoded_block[1228] ^ uncoded_block[1234];
  wire _11181 = uncoded_block[1235] ^ uncoded_block[1238];
  wire _11182 = _11180 ^ _11181;
  wire _11183 = _6536 ^ _5229;
  wire _11184 = _11182 ^ _11183;
  wire _11185 = _11179 ^ _11184;
  wire _11186 = _7778 ^ _2235;
  wire _11187 = _11186 ^ _7782;
  wire _11188 = uncoded_block[1267] ^ uncoded_block[1269];
  wire _11189 = _1458 ^ _11188;
  wire _11190 = _5905 ^ _9539;
  wire _11191 = _11189 ^ _11190;
  wire _11192 = _11187 ^ _11191;
  wire _11193 = _11185 ^ _11192;
  wire _11194 = _7183 ^ _6557;
  wire _11195 = uncoded_block[1287] ^ uncoded_block[1290];
  wire _11196 = _5243 ^ _11195;
  wire _11197 = _11194 ^ _11196;
  wire _11198 = _3015 ^ _3017;
  wire _11199 = _8984 ^ _2254;
  wire _11200 = _11198 ^ _11199;
  wire _11201 = _11197 ^ _11200;
  wire _11202 = uncoded_block[1304] ^ uncoded_block[1313];
  wire _11203 = _11202 ^ _6574;
  wire _11204 = _4540 ^ _5927;
  wire _11205 = _11203 ^ _11204;
  wire _11206 = _8411 ^ _4545;
  wire _11207 = uncoded_block[1330] ^ uncoded_block[1334];
  wire _11208 = _11207 ^ _3034;
  wire _11209 = _11206 ^ _11208;
  wire _11210 = _11205 ^ _11209;
  wire _11211 = _11201 ^ _11210;
  wire _11212 = _11193 ^ _11211;
  wire _11213 = _11176 ^ _11212;
  wire _11214 = _9563 ^ _4553;
  wire _11215 = uncoded_block[1343] ^ uncoded_block[1345];
  wire _11216 = _5262 ^ _11215;
  wire _11217 = _11214 ^ _11216;
  wire _11218 = uncoded_block[1348] ^ uncoded_block[1350];
  wire _11219 = _11218 ^ _670;
  wire _11220 = uncoded_block[1353] ^ uncoded_block[1357];
  wire _11221 = _11220 ^ _7821;
  wire _11222 = _11219 ^ _11221;
  wire _11223 = _11217 ^ _11222;
  wire _11224 = uncoded_block[1364] ^ uncoded_block[1366];
  wire _11225 = _1504 ^ _11224;
  wire _11226 = uncoded_block[1370] ^ uncoded_block[1371];
  wire _11227 = _11226 ^ _2289;
  wire _11228 = _11225 ^ _11227;
  wire _11229 = _7824 ^ _688;
  wire _11230 = _1513 ^ _694;
  wire _11231 = _11229 ^ _11230;
  wire _11232 = _11228 ^ _11231;
  wire _11233 = _11223 ^ _11232;
  wire _11234 = uncoded_block[1399] ^ uncoded_block[1404];
  wire _11235 = _1516 ^ _11234;
  wire _11236 = uncoded_block[1405] ^ uncoded_block[1409];
  wire _11237 = _11236 ^ _7229;
  wire _11238 = _11235 ^ _11237;
  wire _11239 = uncoded_block[1425] ^ uncoded_block[1427];
  wire _11240 = _4583 ^ _11239;
  wire _11241 = _10684 ^ _5299;
  wire _11242 = _11240 ^ _11241;
  wire _11243 = _11238 ^ _11242;
  wire _11244 = _2321 ^ _3864;
  wire _11245 = _2320 ^ _11244;
  wire _11246 = uncoded_block[1449] ^ uncoded_block[1451];
  wire _11247 = uncoded_block[1453] ^ uncoded_block[1455];
  wire _11248 = _11246 ^ _11247;
  wire _11249 = uncoded_block[1456] ^ uncoded_block[1460];
  wire _11250 = _11249 ^ _2336;
  wire _11251 = _11248 ^ _11250;
  wire _11252 = _11245 ^ _11251;
  wire _11253 = _11243 ^ _11252;
  wire _11254 = _11233 ^ _11253;
  wire _11255 = uncoded_block[1471] ^ uncoded_block[1473];
  wire _11256 = _2338 ^ _11255;
  wire _11257 = _733 ^ _2342;
  wire _11258 = _11256 ^ _11257;
  wire _11259 = _4607 ^ _5321;
  wire _11260 = uncoded_block[1497] ^ uncoded_block[1499];
  wire _11261 = _742 ^ _11260;
  wire _11262 = _11259 ^ _11261;
  wire _11263 = _11258 ^ _11262;
  wire _11264 = uncoded_block[1505] ^ uncoded_block[1507];
  wire _11265 = _3893 ^ _11264;
  wire _11266 = uncoded_block[1509] ^ uncoded_block[1513];
  wire _11267 = uncoded_block[1515] ^ uncoded_block[1518];
  wire _11268 = _11266 ^ _11267;
  wire _11269 = _11265 ^ _11268;
  wire _11270 = uncoded_block[1521] ^ uncoded_block[1524];
  wire _11271 = _11270 ^ _3122;
  wire _11272 = uncoded_block[1527] ^ uncoded_block[1530];
  wire _11273 = _11272 ^ _6650;
  wire _11274 = _11271 ^ _11273;
  wire _11275 = _11269 ^ _11274;
  wire _11276 = _11263 ^ _11275;
  wire _11277 = _3128 ^ _1593;
  wire _11278 = uncoded_block[1552] ^ uncoded_block[1556];
  wire _11279 = _9067 ^ _11278;
  wire _11280 = _11277 ^ _11279;
  wire _11281 = uncoded_block[1557] ^ uncoded_block[1558];
  wire _11282 = _11281 ^ _7888;
  wire _11283 = uncoded_block[1562] ^ uncoded_block[1565];
  wire _11284 = uncoded_block[1566] ^ uncoded_block[1567];
  wire _11285 = _11283 ^ _11284;
  wire _11286 = _11282 ^ _11285;
  wire _11287 = _11280 ^ _11286;
  wire _11288 = _4645 ^ _1608;
  wire _11289 = uncoded_block[1578] ^ uncoded_block[1584];
  wire _11290 = _11289 ^ _788;
  wire _11291 = _11288 ^ _11290;
  wire _11292 = uncoded_block[1592] ^ uncoded_block[1594];
  wire _11293 = _3145 ^ _11292;
  wire _11294 = uncoded_block[1595] ^ uncoded_block[1597];
  wire _11295 = uncoded_block[1598] ^ uncoded_block[1599];
  wire _11296 = _11294 ^ _11295;
  wire _11297 = _11293 ^ _11296;
  wire _11298 = _11291 ^ _11297;
  wire _11299 = _11287 ^ _11298;
  wire _11300 = _11276 ^ _11299;
  wire _11301 = _11254 ^ _11300;
  wire _11302 = _11213 ^ _11301;
  wire _11303 = uncoded_block[1606] ^ uncoded_block[1609];
  wire _11304 = _3936 ^ _11303;
  wire _11305 = _11304 ^ _10182;
  wire _11306 = _7298 ^ _807;
  wire _11307 = uncoded_block[1627] ^ uncoded_block[1630];
  wire _11308 = _11307 ^ _5388;
  wire _11309 = _11306 ^ _11308;
  wire _11310 = _11305 ^ _11309;
  wire _11311 = uncoded_block[1642] ^ uncoded_block[1648];
  wire _11312 = _4668 ^ _11311;
  wire _11313 = _10757 ^ _9106;
  wire _11314 = _11312 ^ _11313;
  wire _11315 = _3175 ^ _2422;
  wire _11316 = _7926 ^ _11315;
  wire _11317 = _11314 ^ _11316;
  wire _11318 = _11310 ^ _11317;
  wire _11319 = uncoded_block[1674] ^ uncoded_block[1676];
  wire _11320 = _8521 ^ _11319;
  wire _11321 = uncoded_block[1678] ^ uncoded_block[1679];
  wire _11322 = _11321 ^ _9113;
  wire _11323 = _11320 ^ _11322;
  wire _11324 = uncoded_block[1685] ^ uncoded_block[1688];
  wire _11325 = uncoded_block[1691] ^ uncoded_block[1693];
  wire _11326 = _11324 ^ _11325;
  wire _11327 = uncoded_block[1698] ^ uncoded_block[1699];
  wire _11328 = uncoded_block[1700] ^ uncoded_block[1706];
  wire _11329 = _11327 ^ _11328;
  wire _11330 = _11326 ^ _11329;
  wire _11331 = _11323 ^ _11330;
  wire _11332 = uncoded_block[1707] ^ uncoded_block[1711];
  wire _11333 = uncoded_block[1712] ^ uncoded_block[1715];
  wire _11334 = _11332 ^ _11333;
  wire _11335 = _11334 ^ uncoded_block[1718];
  wire _11336 = _11331 ^ _11335;
  wire _11337 = _11318 ^ _11336;
  wire _11338 = _11302 ^ _11337;
  wire _11339 = _11136 ^ _11338;
  wire _11340 = _0 ^ _866;
  wire _11341 = _9135 ^ _10226;
  wire _11342 = _11340 ^ _11341;
  wire _11343 = uncoded_block[23] ^ uncoded_block[25];
  wire _11344 = uncoded_block[27] ^ uncoded_block[28];
  wire _11345 = _11343 ^ _11344;
  wire _11346 = uncoded_block[29] ^ uncoded_block[34];
  wire _11347 = uncoded_block[35] ^ uncoded_block[38];
  wire _11348 = _11346 ^ _11347;
  wire _11349 = _11345 ^ _11348;
  wire _11350 = _11342 ^ _11349;
  wire _11351 = _23 ^ _5433;
  wire _11352 = uncoded_block[55] ^ uncoded_block[59];
  wire _11353 = _5435 ^ _11352;
  wire _11354 = _11351 ^ _11353;
  wire _11355 = uncoded_block[60] ^ uncoded_block[64];
  wire _11356 = _11355 ^ _9705;
  wire _11357 = uncoded_block[67] ^ uncoded_block[68];
  wire _11358 = _11357 ^ _896;
  wire _11359 = _11356 ^ _11358;
  wire _11360 = _11354 ^ _11359;
  wire _11361 = _11350 ^ _11360;
  wire _11362 = _897 ^ _39;
  wire _11363 = uncoded_block[78] ^ uncoded_block[81];
  wire _11364 = uncoded_block[83] ^ uncoded_block[84];
  wire _11365 = _11363 ^ _11364;
  wire _11366 = _11362 ^ _11365;
  wire _11367 = _1718 ^ _908;
  wire _11368 = _910 ^ _4031;
  wire _11369 = _11367 ^ _11368;
  wire _11370 = _11366 ^ _11369;
  wire _11371 = _4032 ^ _7990;
  wire _11372 = _54 ^ _9721;
  wire _11373 = _11371 ^ _11372;
  wire _11374 = uncoded_block[125] ^ uncoded_block[128];
  wire _11375 = _10821 ^ _11374;
  wire _11376 = _4042 ^ _9177;
  wire _11377 = _11375 ^ _11376;
  wire _11378 = _11373 ^ _11377;
  wire _11379 = _11370 ^ _11378;
  wire _11380 = _11361 ^ _11379;
  wire _11381 = uncoded_block[142] ^ uncoded_block[145];
  wire _11382 = _6136 ^ _11381;
  wire _11383 = uncoded_block[147] ^ uncoded_block[149];
  wire _11384 = _11383 ^ _70;
  wire _11385 = _11382 ^ _11384;
  wire _11386 = _3269 ^ _7397;
  wire _11387 = _9188 ^ _4053;
  wire _11388 = _11386 ^ _11387;
  wire _11389 = _11385 ^ _11388;
  wire _11390 = uncoded_block[167] ^ uncoded_block[169];
  wire _11391 = _2516 ^ _11390;
  wire _11392 = uncoded_block[172] ^ uncoded_block[175];
  wire _11393 = _11392 ^ _940;
  wire _11394 = _11391 ^ _11393;
  wire _11395 = uncoded_block[180] ^ uncoded_block[184];
  wire _11396 = _11395 ^ _1759;
  wire _11397 = _945 ^ _4773;
  wire _11398 = _11396 ^ _11397;
  wire _11399 = _11394 ^ _11398;
  wire _11400 = _11389 ^ _11399;
  wire _11401 = _3283 ^ _7411;
  wire _11402 = uncoded_block[197] ^ uncoded_block[199];
  wire _11403 = _11402 ^ _10849;
  wire _11404 = _11401 ^ _11403;
  wire _11405 = uncoded_block[207] ^ uncoded_block[209];
  wire _11406 = _10278 ^ _11405;
  wire _11407 = _11406 ^ _4075;
  wire _11408 = _11404 ^ _11407;
  wire _11409 = uncoded_block[218] ^ uncoded_block[222];
  wire _11410 = uncoded_block[225] ^ uncoded_block[227];
  wire _11411 = _11409 ^ _11410;
  wire _11412 = _11411 ^ _8030;
  wire _11413 = _1778 ^ _9756;
  wire _11414 = _11413 ^ _10294;
  wire _11415 = _11412 ^ _11414;
  wire _11416 = _11408 ^ _11415;
  wire _11417 = _11400 ^ _11416;
  wire _11418 = _11380 ^ _11417;
  wire _11419 = uncoded_block[253] ^ uncoded_block[254];
  wire _11420 = _11419 ^ _3311;
  wire _11421 = uncoded_block[266] ^ uncoded_block[268];
  wire _11422 = _6831 ^ _11421;
  wire _11423 = _11420 ^ _11422;
  wire _11424 = uncoded_block[282] ^ uncoded_block[283];
  wire _11425 = _5515 ^ _11424;
  wire _11426 = _8625 ^ _11425;
  wire _11427 = _11423 ^ _11426;
  wire _11428 = uncoded_block[284] ^ uncoded_block[286];
  wire _11429 = uncoded_block[287] ^ uncoded_block[291];
  wire _11430 = _11428 ^ _11429;
  wire _11431 = _11430 ^ _4821;
  wire _11432 = _1806 ^ _8051;
  wire _11433 = uncoded_block[305] ^ uncoded_block[309];
  wire _11434 = uncoded_block[310] ^ uncoded_block[315];
  wire _11435 = _11433 ^ _11434;
  wire _11436 = _11432 ^ _11435;
  wire _11437 = _11431 ^ _11436;
  wire _11438 = _11427 ^ _11437;
  wire _11439 = uncoded_block[316] ^ uncoded_block[317];
  wire _11440 = _11439 ^ _6208;
  wire _11441 = uncoded_block[322] ^ uncoded_block[323];
  wire _11442 = _11441 ^ _9780;
  wire _11443 = _11440 ^ _11442;
  wire _11444 = uncoded_block[327] ^ uncoded_block[328];
  wire _11445 = _11444 ^ _2586;
  wire _11446 = uncoded_block[333] ^ uncoded_block[336];
  wire _11447 = _11446 ^ _7463;
  wire _11448 = _11445 ^ _11447;
  wire _11449 = _11443 ^ _11448;
  wire _11450 = uncoded_block[342] ^ uncoded_block[343];
  wire _11451 = _9242 ^ _11450;
  wire _11452 = _6218 ^ _1023;
  wire _11453 = _11451 ^ _11452;
  wire _11454 = uncoded_block[349] ^ uncoded_block[352];
  wire _11455 = uncoded_block[353] ^ uncoded_block[355];
  wire _11456 = _11454 ^ _11455;
  wire _11457 = uncoded_block[358] ^ uncoded_block[361];
  wire _11458 = _2602 ^ _11457;
  wire _11459 = _11456 ^ _11458;
  wire _11460 = _11453 ^ _11459;
  wire _11461 = _11449 ^ _11460;
  wire _11462 = _11438 ^ _11461;
  wire _11463 = uncoded_block[362] ^ uncoded_block[365];
  wire _11464 = _11463 ^ _8076;
  wire _11465 = _6873 ^ _10898;
  wire _11466 = _11464 ^ _11465;
  wire _11467 = _3377 ^ _1846;
  wire _11468 = _5554 ^ _1847;
  wire _11469 = _11467 ^ _11468;
  wire _11470 = _11466 ^ _11469;
  wire _11471 = uncoded_block[400] ^ uncoded_block[404];
  wire _11472 = _1849 ^ _11471;
  wire _11473 = uncoded_block[410] ^ uncoded_block[412];
  wire _11474 = _9810 ^ _11473;
  wire _11475 = _11472 ^ _11474;
  wire _11476 = uncoded_block[416] ^ uncoded_block[419];
  wire _11477 = uncoded_block[420] ^ uncoded_block[422];
  wire _11478 = _11476 ^ _11477;
  wire _11479 = uncoded_block[424] ^ uncoded_block[426];
  wire _11480 = _11479 ^ _6894;
  wire _11481 = _11478 ^ _11480;
  wire _11482 = _11475 ^ _11481;
  wire _11483 = _11470 ^ _11482;
  wire _11484 = _8098 ^ _9275;
  wire _11485 = _6256 ^ _11484;
  wire _11486 = uncoded_block[447] ^ uncoded_block[448];
  wire _11487 = _11486 ^ _4177;
  wire _11488 = _2650 ^ _1870;
  wire _11489 = _11487 ^ _11488;
  wire _11490 = _11485 ^ _11489;
  wire _11491 = uncoded_block[463] ^ uncoded_block[465];
  wire _11492 = _2653 ^ _11491;
  wire _11493 = uncoded_block[466] ^ uncoded_block[473];
  wire _11494 = uncoded_block[474] ^ uncoded_block[475];
  wire _11495 = _11493 ^ _11494;
  wire _11496 = _11492 ^ _11495;
  wire _11497 = _5590 ^ _8693;
  wire _11498 = _8694 ^ _4194;
  wire _11499 = _11497 ^ _11498;
  wire _11500 = _11496 ^ _11499;
  wire _11501 = _11490 ^ _11500;
  wire _11502 = _11483 ^ _11501;
  wire _11503 = _11462 ^ _11502;
  wire _11504 = _11418 ^ _11503;
  wire _11505 = _2664 ^ _4903;
  wire _11506 = _3434 ^ _229;
  wire _11507 = _11505 ^ _11506;
  wire _11508 = uncoded_block[510] ^ uncoded_block[514];
  wire _11509 = _6922 ^ _11508;
  wire _11510 = _8706 ^ _9841;
  wire _11511 = _11509 ^ _11510;
  wire _11512 = _11507 ^ _11511;
  wire _11513 = uncoded_block[525] ^ uncoded_block[529];
  wire _11514 = _1108 ^ _11513;
  wire _11515 = _4926 ^ _5619;
  wire _11516 = _11514 ^ _11515;
  wire _11517 = _1908 ^ _6300;
  wire _11518 = uncoded_block[549] ^ uncoded_block[556];
  wire _11519 = _11518 ^ _4937;
  wire _11520 = _11517 ^ _11519;
  wire _11521 = _11516 ^ _11520;
  wire _11522 = _11512 ^ _11521;
  wire _11523 = uncoded_block[560] ^ uncoded_block[566];
  wire _11524 = uncoded_block[567] ^ uncoded_block[575];
  wire _11525 = _11523 ^ _11524;
  wire _11526 = uncoded_block[577] ^ uncoded_block[579];
  wire _11527 = uncoded_block[580] ^ uncoded_block[583];
  wire _11528 = _11526 ^ _11527;
  wire _11529 = _11525 ^ _11528;
  wire _11530 = uncoded_block[589] ^ uncoded_block[594];
  wire _11531 = _3478 ^ _11530;
  wire _11532 = _1939 ^ _2707;
  wire _11533 = _11531 ^ _11532;
  wire _11534 = _11529 ^ _11533;
  wire _11535 = uncoded_block[602] ^ uncoded_block[605];
  wire _11536 = _11535 ^ _2713;
  wire _11537 = _11536 ^ _5654;
  wire _11538 = _6960 ^ _3495;
  wire _11539 = _11538 ^ _10419;
  wire _11540 = _11537 ^ _11539;
  wire _11541 = _11534 ^ _11540;
  wire _11542 = _11522 ^ _11541;
  wire _11543 = uncoded_block[637] ^ uncoded_block[638];
  wire _11544 = _289 ^ _11543;
  wire _11545 = uncoded_block[642] ^ uncoded_block[647];
  wire _11546 = _4255 ^ _11545;
  wire _11547 = _11544 ^ _11546;
  wire _11548 = _305 ^ _3514;
  wire _11549 = _1961 ^ _11548;
  wire _11550 = _11547 ^ _11549;
  wire _11551 = _7582 ^ _7586;
  wire _11552 = uncoded_block[674] ^ uncoded_block[677];
  wire _11553 = _1178 ^ _11552;
  wire _11554 = _11551 ^ _11553;
  wire _11555 = _8180 ^ _6983;
  wire _11556 = uncoded_block[691] ^ uncoded_block[693];
  wire _11557 = uncoded_block[694] ^ uncoded_block[697];
  wire _11558 = _11556 ^ _11557;
  wire _11559 = _11555 ^ _11558;
  wire _11560 = _11554 ^ _11559;
  wire _11561 = _11550 ^ _11560;
  wire _11562 = uncoded_block[699] ^ uncoded_block[700];
  wire _11563 = _11562 ^ _4990;
  wire _11564 = uncoded_block[704] ^ uncoded_block[707];
  wire _11565 = uncoded_block[710] ^ uncoded_block[712];
  wire _11566 = _11564 ^ _11565;
  wire _11567 = _11563 ^ _11566;
  wire _11568 = _1194 ^ _8193;
  wire _11569 = _5690 ^ _1987;
  wire _11570 = _11568 ^ _11569;
  wire _11571 = _11567 ^ _11570;
  wire _11572 = _1988 ^ _10457;
  wire _11573 = uncoded_block[729] ^ uncoded_block[735];
  wire _11574 = _11573 ^ _350;
  wire _11575 = _11572 ^ _11574;
  wire _11576 = uncoded_block[743] ^ uncoded_block[744];
  wire _11577 = _1207 ^ _11576;
  wire _11578 = uncoded_block[745] ^ uncoded_block[754];
  wire _11579 = _11578 ^ _2778;
  wire _11580 = _11577 ^ _11579;
  wire _11581 = _11575 ^ _11580;
  wire _11582 = _11571 ^ _11581;
  wire _11583 = _11561 ^ _11582;
  wire _11584 = _11542 ^ _11583;
  wire _11585 = uncoded_block[760] ^ uncoded_block[767];
  wire _11586 = _359 ^ _11585;
  wire _11587 = _11019 ^ _7019;
  wire _11588 = _11586 ^ _11587;
  wire _11589 = uncoded_block[777] ^ uncoded_block[785];
  wire _11590 = _11589 ^ _3571;
  wire _11591 = uncoded_block[796] ^ uncoded_block[798];
  wire _11592 = _374 ^ _11591;
  wire _11593 = _11590 ^ _11592;
  wire _11594 = _11588 ^ _11593;
  wire _11595 = _9394 ^ _5041;
  wire _11596 = uncoded_block[810] ^ uncoded_block[812];
  wire _11597 = uncoded_block[815] ^ uncoded_block[817];
  wire _11598 = _11596 ^ _11597;
  wire _11599 = _11595 ^ _11598;
  wire _11600 = uncoded_block[820] ^ uncoded_block[824];
  wire _11601 = _2028 ^ _11600;
  wire _11602 = uncoded_block[825] ^ uncoded_block[830];
  wire _11603 = _11602 ^ _400;
  wire _11604 = _11601 ^ _11603;
  wire _11605 = _11599 ^ _11604;
  wire _11606 = _11594 ^ _11605;
  wire _11607 = uncoded_block[835] ^ uncoded_block[840];
  wire _11608 = _11607 ^ _5058;
  wire _11609 = uncoded_block[845] ^ uncoded_block[846];
  wire _11610 = uncoded_block[847] ^ uncoded_block[850];
  wire _11611 = _11609 ^ _11610;
  wire _11612 = _11608 ^ _11611;
  wire _11613 = _6406 ^ _9945;
  wire _11614 = uncoded_block[859] ^ uncoded_block[862];
  wire _11615 = _11614 ^ _9949;
  wire _11616 = _11613 ^ _11615;
  wire _11617 = _11612 ^ _11616;
  wire _11618 = uncoded_block[866] ^ uncoded_block[869];
  wire _11619 = _11618 ^ _8244;
  wire _11620 = uncoded_block[875] ^ uncoded_block[876];
  wire _11621 = uncoded_block[877] ^ uncoded_block[882];
  wire _11622 = _11620 ^ _11621;
  wire _11623 = _11619 ^ _11622;
  wire _11624 = uncoded_block[883] ^ uncoded_block[887];
  wire _11625 = _11624 ^ _11060;
  wire _11626 = uncoded_block[895] ^ uncoded_block[900];
  wire _11627 = uncoded_block[903] ^ uncoded_block[910];
  wire _11628 = _11626 ^ _11627;
  wire _11629 = _11625 ^ _11628;
  wire _11630 = _11623 ^ _11629;
  wire _11631 = _11617 ^ _11630;
  wire _11632 = _11606 ^ _11631;
  wire _11633 = _5092 ^ _439;
  wire _11634 = uncoded_block[922] ^ uncoded_block[926];
  wire _11635 = _11634 ^ _8835;
  wire _11636 = _11633 ^ _11635;
  wire _11637 = _452 ^ _2863;
  wire _11638 = _2080 ^ _11637;
  wire _11639 = _11636 ^ _11638;
  wire _11640 = uncoded_block[947] ^ uncoded_block[953];
  wire _11641 = _455 ^ _11640;
  wire _11642 = uncoded_block[956] ^ uncoded_block[958];
  wire _11643 = uncoded_block[959] ^ uncoded_block[963];
  wire _11644 = _11642 ^ _11643;
  wire _11645 = _11641 ^ _11644;
  wire _11646 = uncoded_block[964] ^ uncoded_block[965];
  wire _11647 = _11646 ^ _9981;
  wire _11648 = uncoded_block[968] ^ uncoded_block[969];
  wire _11649 = uncoded_block[970] ^ uncoded_block[973];
  wire _11650 = _11648 ^ _11649;
  wire _11651 = _11647 ^ _11650;
  wire _11652 = _11645 ^ _11651;
  wire _11653 = _11639 ^ _11652;
  wire _11654 = _470 ^ _5114;
  wire _11655 = _476 ^ _3659;
  wire _11656 = _11654 ^ _11655;
  wire _11657 = _8856 ^ _11101;
  wire _11658 = _483 ^ _8866;
  wire _11659 = _11657 ^ _11658;
  wire _11660 = _11656 ^ _11659;
  wire _11661 = uncoded_block[1008] ^ uncoded_block[1010];
  wire _11662 = _11661 ^ _2117;
  wire _11663 = uncoded_block[1017] ^ uncoded_block[1019];
  wire _11664 = _11663 ^ _8301;
  wire _11665 = _11662 ^ _11664;
  wire _11666 = uncoded_block[1026] ^ uncoded_block[1029];
  wire _11667 = _11666 ^ _4417;
  wire _11668 = uncoded_block[1032] ^ uncoded_block[1034];
  wire _11669 = _11668 ^ _2129;
  wire _11670 = _11667 ^ _11669;
  wire _11671 = _11665 ^ _11670;
  wire _11672 = _11660 ^ _11671;
  wire _11673 = _11653 ^ _11672;
  wire _11674 = _11632 ^ _11673;
  wire _11675 = _11584 ^ _11674;
  wire _11676 = _11504 ^ _11675;
  wire _11677 = uncoded_block[1042] ^ uncoded_block[1044];
  wire _11678 = _1346 ^ _11677;
  wire _11679 = _1356 ^ _7714;
  wire _11680 = _11678 ^ _11679;
  wire _11681 = _2140 ^ _2142;
  wire _11682 = _4432 ^ _11681;
  wire _11683 = _11680 ^ _11682;
  wire _11684 = _3689 ^ _5156;
  wire _11685 = _5831 ^ _7724;
  wire _11686 = _11684 ^ _11685;
  wire _11687 = uncoded_block[1085] ^ uncoded_block[1086];
  wire _11688 = _11687 ^ _2149;
  wire _11689 = uncoded_block[1091] ^ uncoded_block[1095];
  wire _11690 = _4440 ^ _11689;
  wire _11691 = _11688 ^ _11690;
  wire _11692 = _11686 ^ _11691;
  wire _11693 = _11683 ^ _11692;
  wire _11694 = _11139 ^ _3707;
  wire _11695 = _8336 ^ _550;
  wire _11696 = _11694 ^ _11695;
  wire _11697 = _8917 ^ _2167;
  wire _11698 = _8920 ^ _2942;
  wire _11699 = _11697 ^ _11698;
  wire _11700 = _11696 ^ _11699;
  wire _11701 = _1392 ^ _8343;
  wire _11702 = uncoded_block[1131] ^ uncoded_block[1136];
  wire _11703 = _11702 ^ _10593;
  wire _11704 = _11701 ^ _11703;
  wire _11705 = _5182 ^ _2953;
  wire _11706 = _10597 ^ _2186;
  wire _11707 = _11705 ^ _11706;
  wire _11708 = _11704 ^ _11707;
  wire _11709 = _11700 ^ _11708;
  wire _11710 = _11693 ^ _11709;
  wire _11711 = uncoded_block[1157] ^ uncoded_block[1159];
  wire _11712 = _11711 ^ _7748;
  wire _11713 = _11712 ^ _10601;
  wire _11714 = uncoded_block[1170] ^ uncoded_block[1178];
  wire _11715 = _11160 ^ _11714;
  wire _11716 = _8944 ^ _5201;
  wire _11717 = _11715 ^ _11716;
  wire _11718 = _11713 ^ _11717;
  wire _11719 = uncoded_block[1194] ^ uncoded_block[1197];
  wire _11720 = _5203 ^ _11719;
  wire _11721 = uncoded_block[1198] ^ uncoded_block[1199];
  wire _11722 = uncoded_block[1202] ^ uncoded_block[1207];
  wire _11723 = _11721 ^ _11722;
  wire _11724 = _11720 ^ _11723;
  wire _11725 = _5209 ^ _2981;
  wire _11726 = uncoded_block[1214] ^ uncoded_block[1217];
  wire _11727 = _11726 ^ _609;
  wire _11728 = _11725 ^ _11727;
  wire _11729 = _11724 ^ _11728;
  wire _11730 = _11718 ^ _11729;
  wire _11731 = uncoded_block[1225] ^ uncoded_block[1230];
  wire _11732 = uncoded_block[1234] ^ uncoded_block[1238];
  wire _11733 = _11731 ^ _11732;
  wire _11734 = uncoded_block[1244] ^ uncoded_block[1245];
  wire _11735 = _10627 ^ _11734;
  wire _11736 = _11733 ^ _11735;
  wire _11737 = uncoded_block[1250] ^ uncoded_block[1253];
  wire _11738 = _1449 ^ _11737;
  wire _11739 = uncoded_block[1254] ^ uncoded_block[1256];
  wire _11740 = _11739 ^ _7780;
  wire _11741 = _11738 ^ _11740;
  wire _11742 = _11736 ^ _11741;
  wire _11743 = _4514 ^ _5235;
  wire _11744 = _6550 ^ _2239;
  wire _11745 = _11743 ^ _11744;
  wire _11746 = uncoded_block[1270] ^ uncoded_block[1272];
  wire _11747 = _11746 ^ _4523;
  wire _11748 = _1463 ^ _10638;
  wire _11749 = _11747 ^ _11748;
  wire _11750 = _11745 ^ _11749;
  wire _11751 = _11742 ^ _11750;
  wire _11752 = _11730 ^ _11751;
  wire _11753 = _11710 ^ _11752;
  wire _11754 = _638 ^ _8396;
  wire _11755 = _8399 ^ _3801;
  wire _11756 = _11754 ^ _11755;
  wire _11757 = uncoded_block[1296] ^ uncoded_block[1303];
  wire _11758 = _11757 ^ _2255;
  wire _11759 = uncoded_block[1310] ^ uncoded_block[1313];
  wire _11760 = _8991 ^ _11759;
  wire _11761 = _11758 ^ _11760;
  wire _11762 = _11756 ^ _11761;
  wire _11763 = _6574 ^ _5254;
  wire _11764 = uncoded_block[1326] ^ uncoded_block[1328];
  wire _11765 = _11764 ^ _1494;
  wire _11766 = _11763 ^ _11765;
  wire _11767 = _8413 ^ _3034;
  wire _11768 = _11767 ^ _5267;
  wire _11769 = _11766 ^ _11768;
  wire _11770 = _11762 ^ _11769;
  wire _11771 = uncoded_block[1347] ^ uncoded_block[1349];
  wire _11772 = _11771 ^ _1502;
  wire _11773 = uncoded_block[1359] ^ uncoded_block[1364];
  wire _11774 = _6587 ^ _11773;
  wire _11775 = _11772 ^ _11774;
  wire _11776 = uncoded_block[1368] ^ uncoded_block[1370];
  wire _11777 = _679 ^ _11776;
  wire _11778 = _684 ^ _2290;
  wire _11779 = _11777 ^ _11778;
  wire _11780 = _11775 ^ _11779;
  wire _11781 = uncoded_block[1380] ^ uncoded_block[1383];
  wire _11782 = uncoded_block[1386] ^ uncoded_block[1389];
  wire _11783 = _11781 ^ _11782;
  wire _11784 = _3065 ^ _5293;
  wire _11785 = _11783 ^ _11784;
  wire _11786 = uncoded_block[1410] ^ uncoded_block[1414];
  wire _11787 = _11786 ^ _2306;
  wire _11788 = _7836 ^ _11787;
  wire _11789 = _11785 ^ _11788;
  wire _11790 = _11780 ^ _11789;
  wire _11791 = _11770 ^ _11790;
  wire _11792 = uncoded_block[1418] ^ uncoded_block[1420];
  wire _11793 = _11792 ^ _10683;
  wire _11794 = _11793 ^ _10123;
  wire _11795 = _1534 ^ _3857;
  wire _11796 = uncoded_block[1444] ^ uncoded_block[1448];
  wire _11797 = _10130 ^ _11796;
  wire _11798 = _11795 ^ _11797;
  wire _11799 = _11794 ^ _11798;
  wire _11800 = _6620 ^ _2328;
  wire _11801 = _11800 ^ _7242;
  wire _11802 = _3094 ^ _7247;
  wire _11803 = _4603 ^ _2342;
  wire _11804 = _11802 ^ _11803;
  wire _11805 = _11801 ^ _11804;
  wire _11806 = _11799 ^ _11805;
  wire _11807 = uncoded_block[1479] ^ uncoded_block[1484];
  wire _11808 = _11807 ^ _1562;
  wire _11809 = uncoded_block[1489] ^ uncoded_block[1492];
  wire _11810 = _11809 ^ _6631;
  wire _11811 = _11808 ^ _11810;
  wire _11812 = _6634 ^ _7866;
  wire _11813 = uncoded_block[1504] ^ uncoded_block[1506];
  wire _11814 = _11813 ^ _4617;
  wire _11815 = _11812 ^ _11814;
  wire _11816 = _11811 ^ _11815;
  wire _11817 = _5337 ^ _3900;
  wire _11818 = _3122 ^ _1582;
  wire _11819 = _11817 ^ _11818;
  wire _11820 = uncoded_block[1530] ^ uncoded_block[1533];
  wire _11821 = _11820 ^ _3906;
  wire _11822 = _3908 ^ _3128;
  wire _11823 = _11821 ^ _11822;
  wire _11824 = _11819 ^ _11823;
  wire _11825 = _11816 ^ _11824;
  wire _11826 = _11806 ^ _11825;
  wire _11827 = _11791 ^ _11826;
  wire _11828 = _11753 ^ _11827;
  wire _11829 = uncoded_block[1551] ^ uncoded_block[1555];
  wire _11830 = _11829 ^ _6016;
  wire _11831 = _4635 ^ _11830;
  wire _11832 = _774 ^ _776;
  wire _11833 = uncoded_block[1567] ^ uncoded_block[1569];
  wire _11834 = _11833 ^ _5363;
  wire _11835 = _11832 ^ _11834;
  wire _11836 = _11831 ^ _11835;
  wire _11837 = _9080 ^ _3920;
  wire _11838 = uncoded_block[1582] ^ uncoded_block[1585];
  wire _11839 = _2383 ^ _11838;
  wire _11840 = _11837 ^ _11839;
  wire _11841 = uncoded_block[1588] ^ uncoded_block[1594];
  wire _11842 = _1615 ^ _11841;
  wire _11843 = _792 ^ _11295;
  wire _11844 = _11842 ^ _11843;
  wire _11845 = _11840 ^ _11844;
  wire _11846 = _11836 ^ _11845;
  wire _11847 = uncoded_block[1600] ^ uncoded_block[1601];
  wire _11848 = _11847 ^ _8502;
  wire _11849 = uncoded_block[1605] ^ uncoded_block[1608];
  wire _11850 = _11849 ^ _1632;
  wire _11851 = _11848 ^ _11850;
  wire _11852 = _804 ^ _7911;
  wire _11853 = uncoded_block[1621] ^ uncoded_block[1624];
  wire _11854 = uncoded_block[1626] ^ uncoded_block[1631];
  wire _11855 = _11853 ^ _11854;
  wire _11856 = _11852 ^ _11855;
  wire _11857 = _11851 ^ _11856;
  wire _11858 = uncoded_block[1635] ^ uncoded_block[1638];
  wire _11859 = _812 ^ _11858;
  wire _11860 = _6689 ^ _6691;
  wire _11861 = _11859 ^ _11860;
  wire _11862 = uncoded_block[1654] ^ uncoded_block[1657];
  wire _11863 = _3172 ^ _11862;
  wire _11864 = _4680 ^ _7927;
  wire _11865 = _11863 ^ _11864;
  wire _11866 = _11861 ^ _11865;
  wire _11867 = _11857 ^ _11866;
  wire _11868 = _11846 ^ _11867;
  wire _11869 = _5399 ^ _7322;
  wire _11870 = uncoded_block[1680] ^ uncoded_block[1686];
  wire _11871 = _4690 ^ _11870;
  wire _11872 = _11869 ^ _11871;
  wire _11873 = _3189 ^ _9115;
  wire _11874 = uncoded_block[1693] ^ uncoded_block[1698];
  wire _11875 = uncoded_block[1699] ^ uncoded_block[1703];
  wire _11876 = _11874 ^ _11875;
  wire _11877 = _11873 ^ _11876;
  wire _11878 = _11872 ^ _11877;
  wire _11879 = uncoded_block[1709] ^ uncoded_block[1712];
  wire _11880 = _8536 ^ _11879;
  wire _11881 = _854 ^ uncoded_block[1718];
  wire _11882 = _11880 ^ _11881;
  wire _11883 = _11878 ^ _11882;
  wire _11884 = _11868 ^ _11883;
  wire _11885 = _11828 ^ _11884;
  wire _11886 = _11676 ^ _11885;
  wire _11887 = _3 ^ _9135;
  wire _11888 = _11887 ^ _8546;
  wire _11889 = _10226 ^ _3219;
  wire _11890 = uncoded_block[29] ^ uncoded_block[30];
  wire _11891 = _11890 ^ _6095;
  wire _11892 = _11889 ^ _11891;
  wire _11893 = _11888 ^ _11892;
  wire _11894 = uncoded_block[37] ^ uncoded_block[41];
  wire _11895 = _879 ^ _11894;
  wire _11896 = uncoded_block[51] ^ uncoded_block[57];
  wire _11897 = _885 ^ _11896;
  wire _11898 = _11895 ^ _11897;
  wire _11899 = uncoded_block[58] ^ uncoded_block[62];
  wire _11900 = _11899 ^ _10806;
  wire _11901 = _11900 ^ _4018;
  wire _11902 = _11898 ^ _11901;
  wire _11903 = _11893 ^ _11902;
  wire _11904 = uncoded_block[73] ^ uncoded_block[76];
  wire _11905 = uncoded_block[81] ^ uncoded_block[87];
  wire _11906 = _11904 ^ _11905;
  wire _11907 = _7981 ^ _6115;
  wire _11908 = _11906 ^ _11907;
  wire _11909 = uncoded_block[98] ^ uncoded_block[100];
  wire _11910 = _46 ^ _11909;
  wire _11911 = _49 ^ _6120;
  wire _11912 = _11910 ^ _11911;
  wire _11913 = _11908 ^ _11912;
  wire _11914 = _911 ^ _6123;
  wire _11915 = _10256 ^ _6774;
  wire _11916 = _11914 ^ _11915;
  wire _11917 = _9177 ^ _8581;
  wire _11918 = uncoded_block[140] ^ uncoded_block[141];
  wire _11919 = _9729 ^ _11918;
  wire _11920 = _11917 ^ _11919;
  wire _11921 = _11916 ^ _11920;
  wire _11922 = _11913 ^ _11921;
  wire _11923 = _11903 ^ _11922;
  wire _11924 = uncoded_block[142] ^ uncoded_block[146];
  wire _11925 = _11924 ^ _70;
  wire _11926 = _9186 ^ _5470;
  wire _11927 = _11925 ^ _11926;
  wire _11928 = uncoded_block[164] ^ uncoded_block[167];
  wire _11929 = _4053 ^ _11928;
  wire _11930 = _1752 ^ _6149;
  wire _11931 = _11929 ^ _11930;
  wire _11932 = _11927 ^ _11931;
  wire _11933 = uncoded_block[177] ^ uncoded_block[179];
  wire _11934 = _11933 ^ _8009;
  wire _11935 = uncoded_block[182] ^ uncoded_block[187];
  wire _11936 = _11935 ^ _947;
  wire _11937 = _11934 ^ _11936;
  wire _11938 = _4776 ^ _10277;
  wire _11939 = _6801 ^ _10849;
  wire _11940 = _11938 ^ _11939;
  wire _11941 = _11937 ^ _11940;
  wire _11942 = _11932 ^ _11941;
  wire _11943 = uncoded_block[207] ^ uncoded_block[214];
  wire _11944 = _3289 ^ _11943;
  wire _11945 = uncoded_block[226] ^ uncoded_block[230];
  wire _11946 = _4074 ^ _11945;
  wire _11947 = _11944 ^ _11946;
  wire _11948 = _1775 ^ _968;
  wire _11949 = _7423 ^ _2552;
  wire _11950 = _11948 ^ _11949;
  wire _11951 = _11947 ^ _11950;
  wire _11952 = uncoded_block[244] ^ uncoded_block[246];
  wire _11953 = _6172 ^ _11952;
  wire _11954 = uncoded_block[249] ^ uncoded_block[250];
  wire _11955 = _8617 ^ _11954;
  wire _11956 = _11953 ^ _11955;
  wire _11957 = _3309 ^ _2559;
  wire _11958 = _6185 ^ _4098;
  wire _11959 = _11957 ^ _11958;
  wire _11960 = _11956 ^ _11959;
  wire _11961 = _11951 ^ _11960;
  wire _11962 = _11942 ^ _11961;
  wire _11963 = _11923 ^ _11962;
  wire _11964 = _127 ^ _3320;
  wire _11965 = _5512 ^ _1795;
  wire _11966 = _11964 ^ _11965;
  wire _11967 = uncoded_block[281] ^ uncoded_block[282];
  wire _11968 = _6194 ^ _11967;
  wire _11969 = _3327 ^ _10876;
  wire _11970 = _11968 ^ _11969;
  wire _11971 = _11966 ^ _11970;
  wire _11972 = uncoded_block[294] ^ uncoded_block[300];
  wire _11973 = _4819 ^ _11972;
  wire _11974 = _8052 ^ _1002;
  wire _11975 = _11973 ^ _11974;
  wire _11976 = uncoded_block[312] ^ uncoded_block[315];
  wire _11977 = _8056 ^ _11976;
  wire _11978 = _4118 ^ _11441;
  wire _11979 = _11977 ^ _11978;
  wire _11980 = _11975 ^ _11979;
  wire _11981 = _11971 ^ _11980;
  wire _11982 = _152 ^ _11444;
  wire _11983 = uncoded_block[329] ^ uncoded_block[331];
  wire _11984 = uncoded_block[336] ^ uncoded_block[339];
  wire _11985 = _11983 ^ _11984;
  wire _11986 = _11982 ^ _11985;
  wire _11987 = uncoded_block[340] ^ uncoded_block[344];
  wire _11988 = uncoded_block[345] ^ uncoded_block[349];
  wire _11989 = _11987 ^ _11988;
  wire _11990 = uncoded_block[350] ^ uncoded_block[353];
  wire _11991 = _11990 ^ _2602;
  wire _11992 = _11989 ^ _11991;
  wire _11993 = _11986 ^ _11992;
  wire _11994 = _6864 ^ _11463;
  wire _11995 = uncoded_block[366] ^ uncoded_block[376];
  wire _11996 = _11995 ^ _4854;
  wire _11997 = _11994 ^ _11996;
  wire _11998 = _7476 ^ _2612;
  wire _11999 = uncoded_block[384] ^ uncoded_block[386];
  wire _12000 = _11999 ^ _3381;
  wire _12001 = _11998 ^ _12000;
  wire _12002 = _11997 ^ _12001;
  wire _12003 = _11993 ^ _12002;
  wire _12004 = _11981 ^ _12003;
  wire _12005 = uncoded_block[390] ^ uncoded_block[393];
  wire _12006 = uncoded_block[394] ^ uncoded_block[397];
  wire _12007 = _12005 ^ _12006;
  wire _12008 = _4865 ^ _6244;
  wire _12009 = _12007 ^ _12008;
  wire _12010 = uncoded_block[415] ^ uncoded_block[421];
  wire _12011 = _12010 ^ _4164;
  wire _12012 = _8664 ^ _12011;
  wire _12013 = _12009 ^ _12012;
  wire _12014 = _198 ^ _201;
  wire _12015 = uncoded_block[438] ^ uncoded_block[444];
  wire _12016 = _12015 ^ _7498;
  wire _12017 = _12014 ^ _12016;
  wire _12018 = _4883 ^ _3415;
  wire _12019 = _5586 ^ _1079;
  wire _12020 = _12018 ^ _12019;
  wire _12021 = _12017 ^ _12020;
  wire _12022 = _12013 ^ _12021;
  wire _12023 = uncoded_block[468] ^ uncoded_block[470];
  wire _12024 = _12023 ^ _1082;
  wire _12025 = uncoded_block[475] ^ uncoded_block[477];
  wire _12026 = _12025 ^ _1085;
  wire _12027 = _12024 ^ _12026;
  wire _12028 = uncoded_block[481] ^ uncoded_block[483];
  wire _12029 = _12028 ^ _8694;
  wire _12030 = _1091 ^ _4903;
  wire _12031 = _12029 ^ _12030;
  wire _12032 = _12027 ^ _12031;
  wire _12033 = uncoded_block[498] ^ uncoded_block[501];
  wire _12034 = uncoded_block[505] ^ uncoded_block[506];
  wire _12035 = _12033 ^ _12034;
  wire _12036 = _9294 ^ _8122;
  wire _12037 = _12035 ^ _12036;
  wire _12038 = _4918 ^ _6289;
  wire _12039 = uncoded_block[530] ^ uncoded_block[535];
  wire _12040 = _11513 ^ _12039;
  wire _12041 = _12038 ^ _12040;
  wire _12042 = _12037 ^ _12041;
  wire _12043 = _12032 ^ _12042;
  wire _12044 = _12022 ^ _12043;
  wire _12045 = _12004 ^ _12044;
  wire _12046 = _11963 ^ _12045;
  wire _12047 = _3451 ^ _9311;
  wire _12048 = uncoded_block[543] ^ uncoded_block[548];
  wire _12049 = _12048 ^ _8720;
  wire _12050 = _12047 ^ _12049;
  wire _12051 = uncoded_block[556] ^ uncoded_block[558];
  wire _12052 = _8721 ^ _12051;
  wire _12053 = _8725 ^ _3467;
  wire _12054 = _12052 ^ _12053;
  wire _12055 = _12050 ^ _12054;
  wire _12056 = _3468 ^ _4224;
  wire _12057 = uncoded_block[574] ^ uncoded_block[577];
  wire _12058 = _12057 ^ _1133;
  wire _12059 = _12056 ^ _12058;
  wire _12060 = uncoded_block[584] ^ uncoded_block[592];
  wire _12061 = _3475 ^ _12060;
  wire _12062 = _6316 ^ _1939;
  wire _12063 = _12061 ^ _12062;
  wire _12064 = _12059 ^ _12063;
  wire _12065 = _12055 ^ _12064;
  wire _12066 = uncoded_block[597] ^ uncoded_block[599];
  wire _12067 = _12066 ^ _2710;
  wire _12068 = _2713 ^ _7563;
  wire _12069 = _12067 ^ _12068;
  wire _12070 = _1149 ^ _4243;
  wire _12071 = uncoded_block[629] ^ uncoded_block[630];
  wire _12072 = _7568 ^ _12071;
  wire _12073 = _12070 ^ _12072;
  wire _12074 = _12069 ^ _12073;
  wire _12075 = uncoded_block[633] ^ uncoded_block[636];
  wire _12076 = _12075 ^ _11543;
  wire _12077 = _1163 ^ _6336;
  wire _12078 = _12076 ^ _12077;
  wire _12079 = _3505 ^ _10427;
  wire _12080 = uncoded_block[655] ^ uncoded_block[660];
  wire _12081 = uncoded_block[662] ^ uncoded_block[666];
  wire _12082 = _12080 ^ _12081;
  wire _12083 = _12079 ^ _12082;
  wire _12084 = _12078 ^ _12083;
  wire _12085 = _12074 ^ _12084;
  wire _12086 = _12065 ^ _12085;
  wire _12087 = uncoded_block[672] ^ uncoded_block[678];
  wire _12088 = _1174 ^ _12087;
  wire _12089 = uncoded_block[682] ^ uncoded_block[689];
  wire _12090 = _1181 ^ _12089;
  wire _12091 = _12088 ^ _12090;
  wire _12092 = uncoded_block[693] ^ uncoded_block[697];
  wire _12093 = _326 ^ _12092;
  wire _12094 = _11562 ^ _10447;
  wire _12095 = _12093 ^ _12094;
  wire _12096 = _12091 ^ _12095;
  wire _12097 = _3536 ^ _4999;
  wire _12098 = _4997 ^ _12097;
  wire _12099 = _341 ^ _3544;
  wire _12100 = _4286 ^ _5005;
  wire _12101 = _12099 ^ _12100;
  wire _12102 = _12098 ^ _12101;
  wire _12103 = _12096 ^ _12102;
  wire _12104 = _5006 ^ _1206;
  wire _12105 = _352 ^ _5699;
  wire _12106 = _12104 ^ _12105;
  wire _12107 = uncoded_block[746] ^ uncoded_block[749];
  wire _12108 = _12107 ^ _2002;
  wire _12109 = uncoded_block[755] ^ uncoded_block[760];
  wire _12110 = _12109 ^ _8781;
  wire _12111 = _12108 ^ _12110;
  wire _12112 = _12106 ^ _12111;
  wire _12113 = uncoded_block[768] ^ uncoded_block[770];
  wire _12114 = uncoded_block[771] ^ uncoded_block[773];
  wire _12115 = _12113 ^ _12114;
  wire _12116 = _366 ^ _12115;
  wire _12117 = uncoded_block[774] ^ uncoded_block[777];
  wire _12118 = _12117 ^ _368;
  wire _12119 = _1224 ^ _2019;
  wire _12120 = _12118 ^ _12119;
  wire _12121 = _12116 ^ _12120;
  wire _12122 = _12112 ^ _12121;
  wire _12123 = _12103 ^ _12122;
  wire _12124 = _12086 ^ _12123;
  wire _12125 = _2799 ^ _7628;
  wire _12126 = uncoded_block[800] ^ uncoded_block[803];
  wire _12127 = uncoded_block[805] ^ uncoded_block[806];
  wire _12128 = _12126 ^ _12127;
  wire _12129 = _12125 ^ _12128;
  wire _12130 = _1238 ^ _11596;
  wire _12131 = uncoded_block[818] ^ uncoded_block[821];
  wire _12132 = _11030 ^ _12131;
  wire _12133 = _12130 ^ _12132;
  wire _12134 = _12129 ^ _12133;
  wire _12135 = uncoded_block[827] ^ uncoded_block[829];
  wire _12136 = _11034 ^ _12135;
  wire _12137 = uncoded_block[830] ^ uncoded_block[834];
  wire _12138 = uncoded_block[836] ^ uncoded_block[837];
  wire _12139 = _12137 ^ _12138;
  wire _12140 = _12136 ^ _12139;
  wire _12141 = uncoded_block[848] ^ uncoded_block[850];
  wire _12142 = _7047 ^ _12141;
  wire _12143 = _7044 ^ _12142;
  wire _12144 = _12140 ^ _12143;
  wire _12145 = _12134 ^ _12144;
  wire _12146 = uncoded_block[851] ^ uncoded_block[853];
  wire _12147 = _12146 ^ _7049;
  wire _12148 = _2824 ^ _5069;
  wire _12149 = _12147 ^ _12148;
  wire _12150 = uncoded_block[869] ^ uncoded_block[871];
  wire _12151 = uncoded_block[875] ^ uncoded_block[878];
  wire _12152 = _12150 ^ _12151;
  wire _12153 = _4351 ^ _423;
  wire _12154 = _12152 ^ _12153;
  wire _12155 = _12149 ^ _12154;
  wire _12156 = _11059 ^ _4354;
  wire _12157 = _1277 ^ _8250;
  wire _12158 = _12156 ^ _12157;
  wire _12159 = uncoded_block[903] ^ uncoded_block[906];
  wire _12160 = _12159 ^ _2070;
  wire _12161 = _2845 ^ _12160;
  wire _12162 = _12158 ^ _12161;
  wire _12163 = _12155 ^ _12162;
  wire _12164 = _12145 ^ _12163;
  wire _12165 = uncoded_block[910] ^ uncoded_block[916];
  wire _12166 = _12165 ^ _439;
  wire _12167 = _5766 ^ _5772;
  wire _12168 = _12166 ^ _12167;
  wire _12169 = uncoded_block[931] ^ uncoded_block[936];
  wire _12170 = _12169 ^ _452;
  wire _12171 = uncoded_block[942] ^ uncoded_block[943];
  wire _12172 = _9971 ^ _12171;
  wire _12173 = _12170 ^ _12172;
  wire _12174 = _12168 ^ _12173;
  wire _12175 = uncoded_block[949] ^ uncoded_block[952];
  wire _12176 = _456 ^ _12175;
  wire _12177 = _461 ^ _2871;
  wire _12178 = _12176 ^ _12177;
  wire _12179 = uncoded_block[963] ^ uncoded_block[964];
  wire _12180 = uncoded_block[965] ^ uncoded_block[967];
  wire _12181 = _12179 ^ _12180;
  wire _12182 = _468 ^ _8853;
  wire _12183 = _12181 ^ _12182;
  wire _12184 = _12178 ^ _12183;
  wire _12185 = _12174 ^ _12184;
  wire _12186 = uncoded_block[985] ^ uncoded_block[986];
  wire _12187 = _5792 ^ _12186;
  wire _12188 = uncoded_block[989] ^ uncoded_block[999];
  wire _12189 = _8856 ^ _12188;
  wire _12190 = _12187 ^ _12189;
  wire _12191 = _4405 ^ _4410;
  wire _12192 = _485 ^ _12191;
  wire _12193 = _12190 ^ _12192;
  wire _12194 = _8868 ^ _5135;
  wire _12195 = _9454 ^ _495;
  wire _12196 = _12194 ^ _12195;
  wire _12197 = _6472 ^ _11668;
  wire _12198 = uncoded_block[1036] ^ uncoded_block[1037];
  wire _12199 = uncoded_block[1038] ^ uncoded_block[1041];
  wire _12200 = _12198 ^ _12199;
  wire _12201 = _12197 ^ _12200;
  wire _12202 = _12196 ^ _12201;
  wire _12203 = _12193 ^ _12202;
  wire _12204 = _12185 ^ _12203;
  wire _12205 = _12164 ^ _12204;
  wire _12206 = _12124 ^ _12205;
  wire _12207 = _12046 ^ _12206;
  wire _12208 = uncoded_block[1042] ^ uncoded_block[1046];
  wire _12209 = _12208 ^ _2134;
  wire _12210 = _2136 ^ _1359;
  wire _12211 = _12209 ^ _12210;
  wire _12212 = _1360 ^ _10566;
  wire _12213 = uncoded_block[1067] ^ uncoded_block[1069];
  wire _12214 = _2917 ^ _12213;
  wire _12215 = _12212 ^ _12214;
  wire _12216 = _12211 ^ _12215;
  wire _12217 = uncoded_block[1071] ^ uncoded_block[1073];
  wire _12218 = _12217 ^ _2924;
  wire _12219 = uncoded_block[1080] ^ uncoded_block[1082];
  wire _12220 = _12219 ^ _533;
  wire _12221 = _12218 ^ _12220;
  wire _12222 = uncoded_block[1089] ^ uncoded_block[1095];
  wire _12223 = _534 ^ _12222;
  wire _12224 = uncoded_block[1099] ^ uncoded_block[1102];
  wire _12225 = _5843 ^ _12224;
  wire _12226 = _12223 ^ _12225;
  wire _12227 = _12221 ^ _12226;
  wire _12228 = _12216 ^ _12227;
  wire _12229 = _3708 ^ _2164;
  wire _12230 = _4451 ^ _2938;
  wire _12231 = _12229 ^ _12230;
  wire _12232 = uncoded_block[1120] ^ uncoded_block[1125];
  wire _12233 = _11147 ^ _12232;
  wire _12234 = uncoded_block[1127] ^ uncoded_block[1133];
  wire _12235 = _12234 ^ _564;
  wire _12236 = _12233 ^ _12235;
  wire _12237 = _12231 ^ _12236;
  wire _12238 = _3721 ^ _2952;
  wire _12239 = _2953 ^ _5862;
  wire _12240 = _12238 ^ _12239;
  wire _12241 = uncoded_block[1149] ^ uncoded_block[1153];
  wire _12242 = _12241 ^ _3727;
  wire _12243 = uncoded_block[1156] ^ uncoded_block[1159];
  wire _12244 = _12243 ^ _2958;
  wire _12245 = _12242 ^ _12244;
  wire _12246 = _12240 ^ _12245;
  wire _12247 = _12237 ^ _12246;
  wire _12248 = _12228 ^ _12247;
  wire _12249 = _6511 ^ _11160;
  wire _12250 = _11161 ^ _3739;
  wire _12251 = _12249 ^ _12250;
  wire _12252 = _585 ^ _10608;
  wire _12253 = _592 ^ _2200;
  wire _12254 = _12252 ^ _12253;
  wire _12255 = _12251 ^ _12254;
  wire _12256 = uncoded_block[1191] ^ uncoded_block[1198];
  wire _12257 = _12256 ^ _2206;
  wire _12258 = uncoded_block[1203] ^ uncoded_block[1210];
  wire _12259 = uncoded_block[1211] ^ uncoded_block[1214];
  wire _12260 = _12258 ^ _12259;
  wire _12261 = _12257 ^ _12260;
  wire _12262 = _5215 ^ _11731;
  wire _12263 = _2221 ^ _12262;
  wire _12264 = _12261 ^ _12263;
  wire _12265 = _12255 ^ _12264;
  wire _12266 = _2225 ^ _5219;
  wire _12267 = _8382 ^ _5229;
  wire _12268 = _12266 ^ _12267;
  wire _12269 = uncoded_block[1256] ^ uncoded_block[1268];
  wire _12270 = _5231 ^ _12269;
  wire _12271 = _9533 ^ _9538;
  wire _12272 = _12270 ^ _12271;
  wire _12273 = _12268 ^ _12272;
  wire _12274 = _5908 ^ _631;
  wire _12275 = _4525 ^ _638;
  wire _12276 = _12274 ^ _12275;
  wire _12277 = _5243 ^ _641;
  wire _12278 = _7193 ^ _7799;
  wire _12279 = _12277 ^ _12278;
  wire _12280 = _12276 ^ _12279;
  wire _12281 = _12273 ^ _12280;
  wire _12282 = _12265 ^ _12281;
  wire _12283 = _12248 ^ _12282;
  wire _12284 = _2254 ^ _6571;
  wire _12285 = _649 ^ _4539;
  wire _12286 = _12284 ^ _12285;
  wire _12287 = uncoded_block[1318] ^ uncoded_block[1320];
  wire _12288 = _2262 ^ _12287;
  wire _12289 = _3814 ^ _656;
  wire _12290 = _12288 ^ _12289;
  wire _12291 = _12286 ^ _12290;
  wire _12292 = uncoded_block[1337] ^ uncoded_block[1340];
  wire _12293 = _1494 ^ _12292;
  wire _12294 = _5262 ^ _5266;
  wire _12295 = _12293 ^ _12294;
  wire _12296 = _4556 ^ _8418;
  wire _12297 = _12296 ^ _7210;
  wire _12298 = _12295 ^ _12297;
  wire _12299 = _12291 ^ _12298;
  wire _12300 = uncoded_block[1360] ^ uncoded_block[1362];
  wire _12301 = _12300 ^ _677;
  wire _12302 = uncoded_block[1367] ^ uncoded_block[1368];
  wire _12303 = _10665 ^ _12302;
  wire _12304 = _12301 ^ _12303;
  wire _12305 = uncoded_block[1375] ^ uncoded_block[1376];
  wire _12306 = _9572 ^ _12305;
  wire _12307 = uncoded_block[1382] ^ uncoded_block[1384];
  wire _12308 = _4564 ^ _12307;
  wire _12309 = _12306 ^ _12308;
  wire _12310 = _12304 ^ _12309;
  wire _12311 = uncoded_block[1385] ^ uncoded_block[1386];
  wire _12312 = _12311 ^ _5950;
  wire _12313 = _6597 ^ _4569;
  wire _12314 = _12312 ^ _12313;
  wire _12315 = uncoded_block[1400] ^ uncoded_block[1403];
  wire _12316 = _5955 ^ _12315;
  wire _12317 = _4578 ^ _5294;
  wire _12318 = _12316 ^ _12317;
  wire _12319 = _12314 ^ _12318;
  wire _12320 = _12310 ^ _12319;
  wire _12321 = _12299 ^ _12320;
  wire _12322 = uncoded_block[1415] ^ uncoded_block[1418];
  wire _12323 = _12322 ^ _7842;
  wire _12324 = _2308 ^ _2311;
  wire _12325 = _12323 ^ _12324;
  wire _12326 = _5968 ^ _1533;
  wire _12327 = _1534 ^ _2318;
  wire _12328 = _12326 ^ _12327;
  wire _12329 = _12325 ^ _12328;
  wire _12330 = uncoded_block[1442] ^ uncoded_block[1447];
  wire _12331 = _4590 ^ _12330;
  wire _12332 = uncoded_block[1451] ^ uncoded_block[1454];
  wire _12333 = _12332 ^ _5309;
  wire _12334 = _12331 ^ _12333;
  wire _12335 = uncoded_block[1457] ^ uncoded_block[1460];
  wire _12336 = _12335 ^ _3871;
  wire _12337 = uncoded_block[1474] ^ uncoded_block[1480];
  wire _12338 = _3097 ^ _12337;
  wire _12339 = _12336 ^ _12338;
  wire _12340 = _12334 ^ _12339;
  wire _12341 = _12329 ^ _12340;
  wire _12342 = uncoded_block[1481] ^ uncoded_block[1483];
  wire _12343 = _12342 ^ _8462;
  wire _12344 = uncoded_block[1497] ^ uncoded_block[1500];
  wire _12345 = _12344 ^ _7866;
  wire _12346 = _12343 ^ _12345;
  wire _12347 = _7259 ^ _3112;
  wire _12348 = uncoded_block[1512] ^ uncoded_block[1518];
  wire _12349 = _5333 ^ _12348;
  wire _12350 = _12347 ^ _12349;
  wire _12351 = _12346 ^ _12350;
  wire _12352 = uncoded_block[1519] ^ uncoded_block[1521];
  wire _12353 = _12352 ^ _4621;
  wire _12354 = uncoded_block[1529] ^ uncoded_block[1534];
  wire _12355 = _5343 ^ _12354;
  wire _12356 = _12353 ^ _12355;
  wire _12357 = uncoded_block[1540] ^ uncoded_block[1546];
  wire _12358 = _5348 ^ _12357;
  wire _12359 = _7275 ^ _7277;
  wire _12360 = _12358 ^ _12359;
  wire _12361 = _12356 ^ _12360;
  wire _12362 = _12351 ^ _12361;
  wire _12363 = _12341 ^ _12362;
  wire _12364 = _12321 ^ _12363;
  wire _12365 = _12283 ^ _12364;
  wire _12366 = _8484 ^ _776;
  wire _12367 = _11284 ^ _4645;
  wire _12368 = _12366 ^ _12367;
  wire _12369 = uncoded_block[1581] ^ uncoded_block[1583];
  wire _12370 = _12369 ^ _1616;
  wire _12371 = _6664 ^ _12370;
  wire _12372 = _12368 ^ _12371;
  wire _12373 = uncoded_block[1603] ^ uncoded_block[1606];
  wire _12374 = _11847 ^ _12373;
  wire _12375 = _11843 ^ _12374;
  wire _12376 = uncoded_block[1618] ^ uncoded_block[1620];
  wire _12377 = _7906 ^ _12376;
  wire _12378 = _11853 ^ _4665;
  wire _12379 = _12377 ^ _12378;
  wire _12380 = _12375 ^ _12379;
  wire _12381 = _12372 ^ _12380;
  wire _12382 = _3166 ^ _9099;
  wire _12383 = uncoded_block[1639] ^ uncoded_block[1641];
  wire _12384 = _12383 ^ _815;
  wire _12385 = _12382 ^ _12384;
  wire _12386 = uncoded_block[1646] ^ uncoded_block[1647];
  wire _12387 = uncoded_block[1649] ^ uncoded_block[1652];
  wire _12388 = _12386 ^ _12387;
  wire _12389 = uncoded_block[1653] ^ uncoded_block[1655];
  wire _12390 = uncoded_block[1656] ^ uncoded_block[1657];
  wire _12391 = _12389 ^ _12390;
  wire _12392 = _12388 ^ _12391;
  wire _12393 = _12385 ^ _12392;
  wire _12394 = uncoded_block[1658] ^ uncoded_block[1662];
  wire _12395 = uncoded_block[1665] ^ uncoded_block[1668];
  wire _12396 = _12394 ^ _12395;
  wire _12397 = _12396 ^ _8523;
  wire _12398 = uncoded_block[1676] ^ uncoded_block[1677];
  wire _12399 = _12398 ^ _3186;
  wire _12400 = uncoded_block[1691] ^ uncoded_block[1698];
  wire _12401 = _12400 ^ _8533;
  wire _12402 = _12399 ^ _12401;
  wire _12403 = _12397 ^ _12402;
  wire _12404 = _12393 ^ _12403;
  wire _12405 = _12381 ^ _12404;
  wire _12406 = _3976 ^ _8536;
  wire _12407 = uncoded_block[1710] ^ uncoded_block[1713];
  wire _12408 = _12407 ^ _854;
  wire _12409 = _12406 ^ _12408;
  wire _12410 = _7946 ^ uncoded_block[1721];
  wire _12411 = _12409 ^ _12410;
  wire _12412 = _12405 ^ _12411;
  wire _12413 = _12365 ^ _12412;
  wire _12414 = _12207 ^ _12413;
  wire _12415 = uncoded_block[1] ^ uncoded_block[4];
  wire _12416 = _12415 ^ _1684;
  wire _12417 = _7 ^ _3998;
  wire _12418 = _12416 ^ _12417;
  wire _12419 = _6087 ^ _3217;
  wire _12420 = uncoded_block[22] ^ uncoded_block[27];
  wire _12421 = _12420 ^ _11890;
  wire _12422 = _12419 ^ _12421;
  wire _12423 = _12418 ^ _12422;
  wire _12424 = _875 ^ _2462;
  wire _12425 = uncoded_block[44] ^ uncoded_block[45];
  wire _12426 = _7965 ^ _12425;
  wire _12427 = _12424 ^ _12426;
  wire _12428 = uncoded_block[47] ^ uncoded_block[52];
  wire _12429 = uncoded_block[53] ^ uncoded_block[55];
  wire _12430 = _12428 ^ _12429;
  wire _12431 = _26 ^ _7365;
  wire _12432 = _12430 ^ _12431;
  wire _12433 = _12427 ^ _12432;
  wire _12434 = _12423 ^ _12433;
  wire _12435 = uncoded_block[64] ^ uncoded_block[65];
  wire _12436 = uncoded_block[67] ^ uncoded_block[72];
  wire _12437 = _12435 ^ _12436;
  wire _12438 = uncoded_block[73] ^ uncoded_block[77];
  wire _12439 = _12438 ^ _11363;
  wire _12440 = _12437 ^ _12439;
  wire _12441 = _41 ^ _4025;
  wire _12442 = uncoded_block[90] ^ uncoded_block[94];
  wire _12443 = uncoded_block[96] ^ uncoded_block[98];
  wire _12444 = _12442 ^ _12443;
  wire _12445 = _12441 ^ _12444;
  wire _12446 = _12440 ^ _12445;
  wire _12447 = uncoded_block[99] ^ uncoded_block[102];
  wire _12448 = _12447 ^ _1721;
  wire _12449 = _4032 ^ _914;
  wire _12450 = _12448 ^ _12449;
  wire _12451 = uncoded_block[120] ^ uncoded_block[121];
  wire _12452 = _2495 ^ _12451;
  wire _12453 = _3255 ^ _1730;
  wire _12454 = _12452 ^ _12453;
  wire _12455 = _12450 ^ _12454;
  wire _12456 = _12446 ^ _12455;
  wire _12457 = _12434 ^ _12456;
  wire _12458 = _1733 ^ _4042;
  wire _12459 = uncoded_block[137] ^ uncoded_block[142];
  wire _12460 = uncoded_block[144] ^ uncoded_block[149];
  wire _12461 = _12459 ^ _12460;
  wire _12462 = _12458 ^ _12461;
  wire _12463 = uncoded_block[162] ^ uncoded_block[164];
  wire _12464 = _2514 ^ _12463;
  wire _12465 = _6782 ^ _12464;
  wire _12466 = _12462 ^ _12465;
  wire _12467 = uncoded_block[168] ^ uncoded_block[172];
  wire _12468 = _8589 ^ _12467;
  wire _12469 = _4057 ^ _85;
  wire _12470 = _12468 ^ _12469;
  wire _12471 = _941 ^ _86;
  wire _12472 = _1759 ^ _945;
  wire _12473 = _12471 ^ _12472;
  wire _12474 = _12470 ^ _12473;
  wire _12475 = _12466 ^ _12474;
  wire _12476 = _5483 ^ _4776;
  wire _12477 = _3284 ^ _94;
  wire _12478 = _12476 ^ _12477;
  wire _12479 = uncoded_block[203] ^ uncoded_block[204];
  wire _12480 = _12479 ^ _10852;
  wire _12481 = _11939 ^ _12480;
  wire _12482 = _12478 ^ _12481;
  wire _12483 = uncoded_block[210] ^ uncoded_block[214];
  wire _12484 = uncoded_block[216] ^ uncoded_block[220];
  wire _12485 = _12483 ^ _12484;
  wire _12486 = _7419 ^ _3299;
  wire _12487 = _12485 ^ _12486;
  wire _12488 = _109 ^ _4081;
  wire _12489 = _7422 ^ _10289;
  wire _12490 = _12488 ^ _12489;
  wire _12491 = _12487 ^ _12490;
  wire _12492 = _12482 ^ _12491;
  wire _12493 = _12475 ^ _12492;
  wire _12494 = _12457 ^ _12493;
  wire _12495 = uncoded_block[237] ^ uncoded_block[239];
  wire _12496 = _12495 ^ _10860;
  wire _12497 = _8616 ^ _7432;
  wire _12498 = _12496 ^ _12497;
  wire _12499 = uncoded_block[255] ^ uncoded_block[261];
  wire _12500 = _4800 ^ _12499;
  wire _12501 = uncoded_block[262] ^ uncoded_block[266];
  wire _12502 = _12501 ^ _127;
  wire _12503 = _12500 ^ _12502;
  wire _12504 = _12498 ^ _12503;
  wire _12505 = _3320 ^ _3324;
  wire _12506 = uncoded_block[279] ^ uncoded_block[281];
  wire _12507 = _12506 ^ _11424;
  wire _12508 = _12505 ^ _12507;
  wire _12509 = uncoded_block[288] ^ uncoded_block[294];
  wire _12510 = _134 ^ _12509;
  wire _12511 = _1807 ^ _4111;
  wire _12512 = _12510 ^ _12511;
  wire _12513 = _12508 ^ _12512;
  wire _12514 = _12504 ^ _12513;
  wire _12515 = uncoded_block[304] ^ uncoded_block[306];
  wire _12516 = uncoded_block[308] ^ uncoded_block[314];
  wire _12517 = _12515 ^ _12516;
  wire _12518 = _146 ^ _149;
  wire _12519 = _12517 ^ _12518;
  wire _12520 = _3346 ^ _4123;
  wire _12521 = uncoded_block[327] ^ uncoded_block[329];
  wire _12522 = _12521 ^ _3352;
  wire _12523 = _12520 ^ _12522;
  wire _12524 = _12519 ^ _12523;
  wire _12525 = _6857 ^ _7463;
  wire _12526 = uncoded_block[342] ^ uncoded_block[348];
  wire _12527 = _9242 ^ _12526;
  wire _12528 = _12525 ^ _12527;
  wire _12529 = _11454 ^ _9249;
  wire _12530 = uncoded_block[360] ^ uncoded_block[362];
  wire _12531 = _12530 ^ _4851;
  wire _12532 = _12529 ^ _12531;
  wire _12533 = _12528 ^ _12532;
  wire _12534 = _12524 ^ _12533;
  wire _12535 = _12514 ^ _12534;
  wire _12536 = uncoded_block[366] ^ uncoded_block[370];
  wire _12537 = _12536 ^ _4140;
  wire _12538 = uncoded_block[379] ^ uncoded_block[381];
  wire _12539 = _12538 ^ _6876;
  wire _12540 = _12537 ^ _12539;
  wire _12541 = uncoded_block[390] ^ uncoded_block[392];
  wire _12542 = _12541 ^ _1048;
  wire _12543 = _3382 ^ _12542;
  wire _12544 = _12540 ^ _12543;
  wire _12545 = uncoded_block[405] ^ uncoded_block[406];
  wire _12546 = _10341 ^ _12545;
  wire _12547 = uncoded_block[409] ^ uncoded_block[413];
  wire _12548 = uncoded_block[414] ^ uncoded_block[418];
  wire _12549 = _12547 ^ _12548;
  wire _12550 = _12546 ^ _12549;
  wire _12551 = uncoded_block[423] ^ uncoded_block[426];
  wire _12552 = _4163 ^ _12551;
  wire _12553 = uncoded_block[427] ^ uncoded_block[433];
  wire _12554 = _12553 ^ _2640;
  wire _12555 = _12552 ^ _12554;
  wire _12556 = _12550 ^ _12555;
  wire _12557 = _12544 ^ _12556;
  wire _12558 = _4169 ^ _3405;
  wire _12559 = uncoded_block[444] ^ uncoded_block[445];
  wire _12560 = _205 ^ _12559;
  wire _12561 = _12558 ^ _12560;
  wire _12562 = uncoded_block[451] ^ uncoded_block[453];
  wire _12563 = _12562 ^ _2650;
  wire _12564 = _213 ^ _4185;
  wire _12565 = _12563 ^ _12564;
  wire _12566 = _12561 ^ _12565;
  wire _12567 = _8683 ^ _9283;
  wire _12568 = _12567 ^ _4892;
  wire _12569 = _11494 ^ _5592;
  wire _12570 = _5593 ^ _1086;
  wire _12571 = _12569 ^ _12570;
  wire _12572 = _12568 ^ _12571;
  wire _12573 = _12566 ^ _12572;
  wire _12574 = _12557 ^ _12573;
  wire _12575 = _12535 ^ _12574;
  wire _12576 = _12494 ^ _12575;
  wire _12577 = uncoded_block[486] ^ uncoded_block[489];
  wire _12578 = uncoded_block[492] ^ uncoded_block[493];
  wire _12579 = _12577 ^ _12578;
  wire _12580 = _12579 ^ _1095;
  wire _12581 = uncoded_block[499] ^ uncoded_block[506];
  wire _12582 = _12581 ^ _10376;
  wire _12583 = _4908 ^ _4910;
  wire _12584 = _12582 ^ _12583;
  wire _12585 = _12580 ^ _12584;
  wire _12586 = uncoded_block[528] ^ uncoded_block[531];
  wire _12587 = _6289 ^ _12586;
  wire _12588 = _8130 ^ _12587;
  wire _12589 = uncoded_block[535] ^ uncoded_block[538];
  wire _12590 = _9309 ^ _12589;
  wire _12591 = uncoded_block[540] ^ uncoded_block[545];
  wire _12592 = uncoded_block[547] ^ uncoded_block[549];
  wire _12593 = _12591 ^ _12592;
  wire _12594 = _12590 ^ _12593;
  wire _12595 = _12588 ^ _12594;
  wire _12596 = _12585 ^ _12595;
  wire _12597 = uncoded_block[552] ^ uncoded_block[562];
  wire _12598 = _247 ^ _12597;
  wire _12599 = uncoded_block[563] ^ uncoded_block[572];
  wire _12600 = _12599 ^ _262;
  wire _12601 = _12598 ^ _12600;
  wire _12602 = uncoded_block[579] ^ uncoded_block[582];
  wire _12603 = _10399 ^ _12602;
  wire _12604 = _266 ^ _4236;
  wire _12605 = _12603 ^ _12604;
  wire _12606 = _12601 ^ _12605;
  wire _12607 = _2706 ^ _9332;
  wire _12608 = uncoded_block[603] ^ uncoded_block[608];
  wire _12609 = uncoded_block[609] ^ uncoded_block[612];
  wire _12610 = _12608 ^ _12609;
  wire _12611 = _12607 ^ _12610;
  wire _12612 = _5652 ^ _1149;
  wire _12613 = _281 ^ _7568;
  wire _12614 = _12612 ^ _12613;
  wire _12615 = _12611 ^ _12614;
  wire _12616 = _12606 ^ _12615;
  wire _12617 = _12596 ^ _12616;
  wire _12618 = uncoded_block[623] ^ uncoded_block[624];
  wire _12619 = _12618 ^ _2720;
  wire _12620 = uncoded_block[628] ^ uncoded_block[632];
  wire _12621 = uncoded_block[633] ^ uncoded_block[638];
  wire _12622 = _12620 ^ _12621;
  wire _12623 = _12619 ^ _12622;
  wire _12624 = uncoded_block[641] ^ uncoded_block[644];
  wire _12625 = _12624 ^ _296;
  wire _12626 = _297 ^ _301;
  wire _12627 = _12625 ^ _12626;
  wire _12628 = _12623 ^ _12627;
  wire _12629 = uncoded_block[654] ^ uncoded_block[657];
  wire _12630 = uncoded_block[662] ^ uncoded_block[663];
  wire _12631 = _12629 ^ _12630;
  wire _12632 = _3516 ^ _1177;
  wire _12633 = _12631 ^ _12632;
  wire _12634 = uncoded_block[675] ^ uncoded_block[679];
  wire _12635 = _1178 ^ _12634;
  wire _12636 = uncoded_block[682] ^ uncoded_block[684];
  wire _12637 = _12636 ^ _4271;
  wire _12638 = _12635 ^ _12637;
  wire _12639 = _12633 ^ _12638;
  wire _12640 = _12628 ^ _12639;
  wire _12641 = uncoded_block[697] ^ uncoded_block[699];
  wire _12642 = _328 ^ _12641;
  wire _12643 = _5681 ^ _12642;
  wire _12644 = uncoded_block[700] ^ uncoded_block[706];
  wire _12645 = uncoded_block[707] ^ uncoded_block[712];
  wire _12646 = _12644 ^ _12645;
  wire _12647 = uncoded_block[714] ^ uncoded_block[716];
  wire _12648 = uncoded_block[720] ^ uncoded_block[723];
  wire _12649 = _12647 ^ _12648;
  wire _12650 = _12646 ^ _12649;
  wire _12651 = _12643 ^ _12650;
  wire _12652 = _10457 ^ _2768;
  wire _12653 = uncoded_block[732] ^ uncoded_block[735];
  wire _12654 = _12653 ^ _3549;
  wire _12655 = _12652 ^ _12654;
  wire _12656 = _5010 ^ _11576;
  wire _12657 = _2775 ^ _4295;
  wire _12658 = _12656 ^ _12657;
  wire _12659 = _12655 ^ _12658;
  wire _12660 = _12651 ^ _12659;
  wire _12661 = _12640 ^ _12660;
  wire _12662 = _12617 ^ _12661;
  wire _12663 = uncoded_block[753] ^ uncoded_block[755];
  wire _12664 = uncoded_block[756] ^ uncoded_block[762];
  wire _12665 = _12663 ^ _12664;
  wire _12666 = _4301 ^ _1218;
  wire _12667 = _12665 ^ _12666;
  wire _12668 = _12114 ^ _2792;
  wire _12669 = uncoded_block[780] ^ uncoded_block[781];
  wire _12670 = _9382 ^ _12669;
  wire _12671 = _12668 ^ _12670;
  wire _12672 = _12667 ^ _12671;
  wire _12673 = uncoded_block[782] ^ uncoded_block[784];
  wire _12674 = _12673 ^ _2018;
  wire _12675 = uncoded_block[788] ^ uncoded_block[790];
  wire _12676 = uncoded_block[792] ^ uncoded_block[795];
  wire _12677 = _12675 ^ _12676;
  wire _12678 = _12674 ^ _12677;
  wire _12679 = uncoded_block[799] ^ uncoded_block[804];
  wire _12680 = _382 ^ _12679;
  wire _12681 = _5042 ^ _2806;
  wire _12682 = _12680 ^ _12681;
  wire _12683 = _12678 ^ _12682;
  wire _12684 = _12672 ^ _12683;
  wire _12685 = _1241 ^ _2029;
  wire _12686 = uncoded_block[830] ^ uncoded_block[833];
  wire _12687 = _6401 ^ _12686;
  wire _12688 = _12685 ^ _12687;
  wire _12689 = _4336 ^ _2035;
  wire _12690 = uncoded_block[848] ^ uncoded_block[852];
  wire _12691 = _11046 ^ _12690;
  wire _12692 = _12689 ^ _12691;
  wire _12693 = _12688 ^ _12692;
  wire _12694 = _8812 ^ _5747;
  wire _12695 = _12694 ^ _1267;
  wire _12696 = uncoded_block[871] ^ uncoded_block[873];
  wire _12697 = _12696 ^ _9954;
  wire _12698 = uncoded_block[880] ^ uncoded_block[887];
  wire _12699 = _12698 ^ _9416;
  wire _12700 = _12697 ^ _12699;
  wire _12701 = _12695 ^ _12700;
  wire _12702 = _12693 ^ _12701;
  wire _12703 = _12684 ^ _12702;
  wire _12704 = uncoded_block[892] ^ uncoded_block[893];
  wire _12705 = _2061 ^ _12704;
  wire _12706 = _4355 ^ _5758;
  wire _12707 = _12705 ^ _12706;
  wire _12708 = uncoded_block[911] ^ uncoded_block[912];
  wire _12709 = _12159 ^ _12708;
  wire _12710 = _2845 ^ _12709;
  wire _12711 = _12707 ^ _12710;
  wire _12712 = uncoded_block[915] ^ uncoded_block[917];
  wire _12713 = _1287 ^ _12712;
  wire _12714 = uncoded_block[919] ^ uncoded_block[923];
  wire _12715 = _12714 ^ _4370;
  wire _12716 = _12713 ^ _12715;
  wire _12717 = uncoded_block[932] ^ uncoded_block[934];
  wire _12718 = _4371 ^ _12717;
  wire _12719 = _8268 ^ _7080;
  wire _12720 = _12718 ^ _12719;
  wire _12721 = _12716 ^ _12720;
  wire _12722 = _12711 ^ _12721;
  wire _12723 = uncoded_block[943] ^ uncoded_block[946];
  wire _12724 = _6439 ^ _12723;
  wire _12725 = uncoded_block[947] ^ uncoded_block[949];
  wire _12726 = uncoded_block[955] ^ uncoded_block[958];
  wire _12727 = _12725 ^ _12726;
  wire _12728 = _12724 ^ _12727;
  wire _12729 = _4385 ^ _1310;
  wire _12730 = _7682 ^ _11649;
  wire _12731 = _12729 ^ _12730;
  wire _12732 = _12728 ^ _12731;
  wire _12733 = uncoded_block[979] ^ uncoded_block[982];
  wire _12734 = uncoded_block[985] ^ uncoded_block[989];
  wire _12735 = _12733 ^ _12734;
  wire _12736 = _11654 ^ _12735;
  wire _12737 = uncoded_block[990] ^ uncoded_block[993];
  wire _12738 = _12737 ^ _8293;
  wire _12739 = _5798 ^ _2111;
  wire _12740 = _12738 ^ _12739;
  wire _12741 = _12736 ^ _12740;
  wire _12742 = _12732 ^ _12741;
  wire _12743 = _12722 ^ _12742;
  wire _12744 = _12703 ^ _12743;
  wire _12745 = _12662 ^ _12744;
  wire _12746 = _12576 ^ _12745;
  wire _12747 = uncoded_block[1003] ^ uncoded_block[1008];
  wire _12748 = _12747 ^ _4409;
  wire _12749 = _12748 ^ _5132;
  wire _12750 = uncoded_block[1017] ^ uncoded_block[1021];
  wire _12751 = _12750 ^ _5137;
  wire _12752 = uncoded_block[1024] ^ uncoded_block[1026];
  wire _12753 = _12752 ^ _1339;
  wire _12754 = _12751 ^ _12753;
  wire _12755 = _12749 ^ _12754;
  wire _12756 = uncoded_block[1030] ^ uncoded_block[1033];
  wire _12757 = _12756 ^ _7707;
  wire _12758 = uncoded_block[1037] ^ uncoded_block[1040];
  wire _12759 = _12758 ^ _512;
  wire _12760 = _12757 ^ _12759;
  wire _12761 = uncoded_block[1044] ^ uncoded_block[1050];
  wire _12762 = uncoded_block[1052] ^ uncoded_block[1053];
  wire _12763 = _12761 ^ _12762;
  wire _12764 = uncoded_block[1056] ^ uncoded_block[1058];
  wire _12765 = _12764 ^ _5825;
  wire _12766 = _12763 ^ _12765;
  wire _12767 = _12760 ^ _12766;
  wire _12768 = _12755 ^ _12767;
  wire _12769 = _2142 ^ _11122;
  wire _12770 = uncoded_block[1072] ^ uncoded_block[1075];
  wire _12771 = _12770 ^ _2147;
  wire _12772 = _12769 ^ _12771;
  wire _12773 = _5834 ^ _7724;
  wire _12774 = uncoded_block[1088] ^ uncoded_block[1090];
  wire _12775 = _533 ^ _12774;
  wire _12776 = _12773 ^ _12775;
  wire _12777 = _12772 ^ _12776;
  wire _12778 = _5840 ^ _3698;
  wire _12779 = _5169 ^ _11142;
  wire _12780 = _12778 ^ _12779;
  wire _12781 = _9484 ^ _4450;
  wire _12782 = uncoded_block[1114] ^ uncoded_block[1115];
  wire _12783 = _4451 ^ _12782;
  wire _12784 = _12781 ^ _12783;
  wire _12785 = _12780 ^ _12784;
  wire _12786 = _12777 ^ _12785;
  wire _12787 = _12768 ^ _12786;
  wire _12788 = uncoded_block[1117] ^ uncoded_block[1122];
  wire _12789 = uncoded_block[1123] ^ uncoded_block[1124];
  wire _12790 = _12788 ^ _12789;
  wire _12791 = uncoded_block[1125] ^ uncoded_block[1128];
  wire _12792 = _12791 ^ _560;
  wire _12793 = _12790 ^ _12792;
  wire _12794 = _5856 ^ _8929;
  wire _12795 = uncoded_block[1138] ^ uncoded_block[1143];
  wire _12796 = _12795 ^ _2180;
  wire _12797 = _12794 ^ _12796;
  wire _12798 = _12793 ^ _12797;
  wire _12799 = _7143 ^ _11157;
  wire _12800 = _7748 ^ _3734;
  wire _12801 = _12799 ^ _12800;
  wire _12802 = uncoded_block[1169] ^ uncoded_block[1175];
  wire _12803 = _7151 ^ _12802;
  wire _12804 = _3740 ^ _2195;
  wire _12805 = _12803 ^ _12804;
  wire _12806 = _12801 ^ _12805;
  wire _12807 = _12798 ^ _12806;
  wire _12808 = uncoded_block[1188] ^ uncoded_block[1189];
  wire _12809 = _12808 ^ _4488;
  wire _12810 = uncoded_block[1195] ^ uncoded_block[1199];
  wire _12811 = _12810 ^ _3753;
  wire _12812 = _12809 ^ _12811;
  wire _12813 = uncoded_block[1213] ^ uncoded_block[1215];
  wire _12814 = _5885 ^ _12813;
  wire _12815 = uncoded_block[1219] ^ uncoded_block[1222];
  wire _12816 = _3763 ^ _12815;
  wire _12817 = _12814 ^ _12816;
  wire _12818 = _12812 ^ _12817;
  wire _12819 = uncoded_block[1226] ^ uncoded_block[1228];
  wire _12820 = uncoded_block[1229] ^ uncoded_block[1234];
  wire _12821 = _12819 ^ _12820;
  wire _12822 = _3771 ^ _1448;
  wire _12823 = _12821 ^ _12822;
  wire _12824 = _5901 ^ _11739;
  wire _12825 = uncoded_block[1258] ^ uncoded_block[1260];
  wire _12826 = _12825 ^ _7178;
  wire _12827 = _12824 ^ _12826;
  wire _12828 = _12823 ^ _12827;
  wire _12829 = _12818 ^ _12828;
  wire _12830 = _12807 ^ _12829;
  wire _12831 = _12787 ^ _12830;
  wire _12832 = uncoded_block[1269] ^ uncoded_block[1272];
  wire _12833 = _12832 ^ _7791;
  wire _12834 = uncoded_block[1279] ^ uncoded_block[1281];
  wire _12835 = _7792 ^ _12834;
  wire _12836 = _12833 ^ _12835;
  wire _12837 = uncoded_block[1282] ^ uncoded_block[1284];
  wire _12838 = uncoded_block[1285] ^ uncoded_block[1291];
  wire _12839 = _12837 ^ _12838;
  wire _12840 = _7193 ^ _4531;
  wire _12841 = _12839 ^ _12840;
  wire _12842 = _12836 ^ _12841;
  wire _12843 = uncoded_block[1298] ^ uncoded_block[1301];
  wire _12844 = _12843 ^ _1472;
  wire _12845 = _1479 ^ _8407;
  wire _12846 = _12844 ^ _12845;
  wire _12847 = uncoded_block[1316] ^ uncoded_block[1319];
  wire _12848 = _12847 ^ _3032;
  wire _12849 = _10655 ^ _6578;
  wire _12850 = _12848 ^ _12849;
  wire _12851 = _12846 ^ _12850;
  wire _12852 = _12842 ^ _12851;
  wire _12853 = _11767 ^ _11214;
  wire _12854 = uncoded_block[1341] ^ uncoded_block[1345];
  wire _12855 = uncoded_block[1347] ^ uncoded_block[1350];
  wire _12856 = _12854 ^ _12855;
  wire _12857 = uncoded_block[1355] ^ uncoded_block[1356];
  wire _12858 = _5938 ^ _12857;
  wire _12859 = _12856 ^ _12858;
  wire _12860 = _12853 ^ _12859;
  wire _12861 = uncoded_block[1362] ^ uncoded_block[1364];
  wire _12862 = _7821 ^ _12861;
  wire _12863 = _10665 ^ _10668;
  wire _12864 = _12862 ^ _12863;
  wire _12865 = _3832 ^ _9572;
  wire _12866 = uncoded_block[1376] ^ uncoded_block[1381];
  wire _12867 = uncoded_block[1388] ^ uncoded_block[1390];
  wire _12868 = _12866 ^ _12867;
  wire _12869 = _12865 ^ _12868;
  wire _12870 = _12864 ^ _12869;
  wire _12871 = _12860 ^ _12870;
  wire _12872 = _12852 ^ _12871;
  wire _12873 = _7828 ^ _3065;
  wire _12874 = uncoded_block[1400] ^ uncoded_block[1409];
  wire _12875 = _4572 ^ _12874;
  wire _12876 = _12873 ^ _12875;
  wire _12877 = uncoded_block[1410] ^ uncoded_block[1413];
  wire _12878 = _12877 ^ _10120;
  wire _12879 = _7844 ^ _10684;
  wire _12880 = _12878 ^ _12879;
  wire _12881 = _12876 ^ _12880;
  wire _12882 = uncoded_block[1434] ^ uncoded_block[1438];
  wire _12883 = _3081 ^ _12882;
  wire _12884 = uncoded_block[1441] ^ uncoded_block[1454];
  wire _12885 = _3861 ^ _12884;
  wire _12886 = _12883 ^ _12885;
  wire _12887 = uncoded_block[1458] ^ uncoded_block[1463];
  wire _12888 = _12887 ^ _9602;
  wire _12889 = _7247 ^ _5983;
  wire _12890 = _12888 ^ _12889;
  wire _12891 = _12886 ^ _12890;
  wire _12892 = _12881 ^ _12891;
  wire _12893 = _3097 ^ _2342;
  wire _12894 = _3884 ^ _739;
  wire _12895 = _12893 ^ _12894;
  wire _12896 = uncoded_block[1493] ^ uncoded_block[1494];
  wire _12897 = _740 ^ _12896;
  wire _12898 = uncoded_block[1495] ^ uncoded_block[1497];
  wire _12899 = uncoded_block[1498] ^ uncoded_block[1501];
  wire _12900 = _12898 ^ _12899;
  wire _12901 = _12897 ^ _12900;
  wire _12902 = _12895 ^ _12901;
  wire _12903 = _3112 ^ _6637;
  wire _12904 = _1575 ^ _9055;
  wire _12905 = _12903 ^ _12904;
  wire _12906 = _9058 ^ _3118;
  wire _12907 = _9626 ^ _6647;
  wire _12908 = _12906 ^ _12907;
  wire _12909 = _12905 ^ _12908;
  wire _12910 = _12902 ^ _12909;
  wire _12911 = _12892 ^ _12910;
  wire _12912 = _12872 ^ _12911;
  wire _12913 = _12831 ^ _12912;
  wire _12914 = uncoded_block[1533] ^ uncoded_block[1534];
  wire _12915 = uncoded_block[1535] ^ uncoded_block[1537];
  wire _12916 = _12914 ^ _12915;
  wire _12917 = uncoded_block[1538] ^ uncoded_block[1540];
  wire _12918 = _12917 ^ _1590;
  wire _12919 = _12916 ^ _12918;
  wire _12920 = uncoded_block[1547] ^ uncoded_block[1552];
  wire _12921 = _5355 ^ _12920;
  wire _12922 = _3131 ^ _11281;
  wire _12923 = _12921 ^ _12922;
  wire _12924 = _12919 ^ _12923;
  wire _12925 = uncoded_block[1569] ^ uncoded_block[1573];
  wire _12926 = _1606 ^ _12925;
  wire _12927 = _11832 ^ _12926;
  wire _12928 = _4648 ^ _3921;
  wire _12929 = uncoded_block[1583] ^ uncoded_block[1588];
  wire _12930 = _6031 ^ _12929;
  wire _12931 = _12928 ^ _12930;
  wire _12932 = _12927 ^ _12931;
  wire _12933 = _12924 ^ _12932;
  wire _12934 = uncoded_block[1589] ^ uncoded_block[1590];
  wire _12935 = uncoded_block[1591] ^ uncoded_block[1594];
  wire _12936 = _12934 ^ _12935;
  wire _12937 = uncoded_block[1600] ^ uncoded_block[1602];
  wire _12938 = _792 ^ _12937;
  wire _12939 = _12936 ^ _12938;
  wire _12940 = uncoded_block[1612] ^ uncoded_block[1614];
  wire _12941 = _9089 ^ _12940;
  wire _12942 = _8503 ^ _12941;
  wire _12943 = _12939 ^ _12942;
  wire _12944 = _10181 ^ _804;
  wire _12945 = _3160 ^ _3941;
  wire _12946 = _12944 ^ _12945;
  wire _12947 = uncoded_block[1626] ^ uncoded_block[1627];
  wire _12948 = _12947 ^ _1636;
  wire _12949 = uncoded_block[1636] ^ uncoded_block[1639];
  wire _12950 = _1639 ^ _12949;
  wire _12951 = _12948 ^ _12950;
  wire _12952 = _12946 ^ _12951;
  wire _12953 = _12943 ^ _12952;
  wire _12954 = _12933 ^ _12953;
  wire _12955 = uncoded_block[1640] ^ uncoded_block[1644];
  wire _12956 = _12955 ^ _6691;
  wire _12957 = uncoded_block[1654] ^ uncoded_block[1658];
  wire _12958 = _4677 ^ _12957;
  wire _12959 = _12956 ^ _12958;
  wire _12960 = uncoded_block[1660] ^ uncoded_block[1663];
  wire _12961 = _12960 ^ _9666;
  wire _12962 = _7928 ^ _6700;
  wire _12963 = _12961 ^ _12962;
  wire _12964 = _12959 ^ _12963;
  wire _12965 = _3965 ^ _2429;
  wire _12966 = _12399 ^ _12965;
  wire _12967 = _11325 ^ _6710;
  wire _12968 = _3973 ^ _3976;
  wire _12969 = _12967 ^ _12968;
  wire _12970 = _12966 ^ _12969;
  wire _12971 = _12964 ^ _12970;
  wire _12972 = uncoded_block[1709] ^ uncoded_block[1714];
  wire _12973 = _2435 ^ _12972;
  wire _12974 = _2441 ^ _3988;
  wire _12975 = _12973 ^ _12974;
  wire _12976 = uncoded_block[1720] ^ uncoded_block[1721];
  wire _12977 = _12976 ^ uncoded_block[1722];
  wire _12978 = _12975 ^ _12977;
  wire _12979 = _12971 ^ _12978;
  wire _12980 = _12954 ^ _12979;
  wire _12981 = _12913 ^ _12980;
  wire _12982 = _12746 ^ _12981;
  wire _12983 = _3213 ^ _7956;
  wire _12984 = _4711 ^ _12983;
  wire _12985 = uncoded_block[18] ^ uncoded_block[23];
  wire _12986 = _8545 ^ _12985;
  wire _12987 = uncoded_block[24] ^ uncoded_block[30];
  wire _12988 = _12987 ^ _6095;
  wire _12989 = _12986 ^ _12988;
  wire _12990 = _12984 ^ _12989;
  wire _12991 = _8549 ^ _2466;
  wire _12992 = _4723 ^ _8554;
  wire _12993 = _12991 ^ _12992;
  wire _12994 = uncoded_block[48] ^ uncoded_block[52];
  wire _12995 = _12994 ^ _5436;
  wire _12996 = uncoded_block[56] ^ uncoded_block[60];
  wire _12997 = _12996 ^ _7365;
  wire _12998 = _12995 ^ _12997;
  wire _12999 = _12993 ^ _12998;
  wire _13000 = _12990 ^ _12999;
  wire _13001 = _35 ^ _7976;
  wire _13002 = _897 ^ _900;
  wire _13003 = _13001 ^ _13002;
  wire _13004 = uncoded_block[81] ^ uncoded_block[86];
  wire _13005 = _7979 ^ _13004;
  wire _13006 = _6113 ^ _1718;
  wire _13007 = _13005 ^ _13006;
  wire _13008 = _13003 ^ _13007;
  wire _13009 = _46 ^ _4745;
  wire _13010 = uncoded_block[102] ^ uncoded_block[105];
  wire _13011 = uncoded_block[106] ^ uncoded_block[109];
  wire _13012 = _13010 ^ _13011;
  wire _13013 = _13009 ^ _13012;
  wire _13014 = uncoded_block[114] ^ uncoded_block[117];
  wire _13015 = _13014 ^ _2498;
  wire _13016 = uncoded_block[121] ^ uncoded_block[125];
  wire _13017 = uncoded_block[126] ^ uncoded_block[129];
  wire _13018 = _13016 ^ _13017;
  wire _13019 = _13015 ^ _13018;
  wire _13020 = _13013 ^ _13019;
  wire _13021 = _13008 ^ _13020;
  wire _13022 = _13000 ^ _13021;
  wire _13023 = _9177 ^ _12459;
  wire _13024 = uncoded_block[148] ^ uncoded_block[154];
  wire _13025 = _2511 ^ _13024;
  wire _13026 = _13023 ^ _13025;
  wire _13027 = uncoded_block[160] ^ uncoded_block[165];
  wire _13028 = _73 ^ _13027;
  wire _13029 = _1751 ^ _7399;
  wire _13030 = _13028 ^ _13029;
  wire _13031 = _13026 ^ _13030;
  wire _13032 = uncoded_block[176] ^ uncoded_block[178];
  wire _13033 = _11392 ^ _13032;
  wire _13034 = uncoded_block[179] ^ uncoded_block[183];
  wire _13035 = _13034 ^ _1759;
  wire _13036 = _13033 ^ _13035;
  wire _13037 = _2529 ^ _2531;
  wire _13038 = uncoded_block[195] ^ uncoded_block[202];
  wire _13039 = _13038 ^ _12479;
  wire _13040 = _13037 ^ _13039;
  wire _13041 = _13036 ^ _13040;
  wire _13042 = _13031 ^ _13041;
  wire _13043 = _4780 ^ _955;
  wire _13044 = _3296 ^ _2543;
  wire _13045 = _13043 ^ _13044;
  wire _13046 = _6168 ^ _7422;
  wire _13047 = _6166 ^ _13046;
  wire _13048 = _13045 ^ _13047;
  wire _13049 = _2552 ^ _9756;
  wire _13050 = uncoded_block[242] ^ uncoded_block[246];
  wire _13051 = _13050 ^ _116;
  wire _13052 = _13049 ^ _13051;
  wire _13053 = uncoded_block[251] ^ uncoded_block[252];
  wire _13054 = _13053 ^ _9761;
  wire _13055 = uncoded_block[258] ^ uncoded_block[259];
  wire _13056 = _13055 ^ _6185;
  wire _13057 = _13054 ^ _13056;
  wire _13058 = _13052 ^ _13057;
  wire _13059 = _13048 ^ _13058;
  wire _13060 = _13042 ^ _13059;
  wire _13061 = _13022 ^ _13060;
  wire _13062 = _6187 ^ _11421;
  wire _13063 = _4102 ^ _1795;
  wire _13064 = _13062 ^ _13063;
  wire _13065 = _10304 ^ _4105;
  wire _13066 = _8632 ^ _5522;
  wire _13067 = _13065 ^ _13066;
  wire _13068 = _13064 ^ _13067;
  wire _13069 = uncoded_block[289] ^ uncoded_block[291];
  wire _13070 = _13069 ^ _7449;
  wire _13071 = uncoded_block[299] ^ uncoded_block[303];
  wire _13072 = _10312 ^ _13071;
  wire _13073 = _13070 ^ _13072;
  wire _13074 = uncoded_block[307] ^ uncoded_block[310];
  wire _13075 = _12515 ^ _13074;
  wire _13076 = _3338 ^ _11439;
  wire _13077 = _13075 ^ _13076;
  wire _13078 = _13073 ^ _13077;
  wire _13079 = _13068 ^ _13078;
  wire _13080 = _1814 ^ _6850;
  wire _13081 = uncoded_block[326] ^ uncoded_block[329];
  wire _13082 = _4123 ^ _13081;
  wire _13083 = _13080 ^ _13082;
  wire _13084 = _2586 ^ _3352;
  wire _13085 = _8646 ^ _9242;
  wire _13086 = _13084 ^ _13085;
  wire _13087 = _13083 ^ _13086;
  wire _13088 = _2595 ^ _159;
  wire _13089 = uncoded_block[353] ^ uncoded_block[356];
  wire _13090 = _2599 ^ _13089;
  wire _13091 = _13088 ^ _13090;
  wire _13092 = _3362 ^ _12530;
  wire _13093 = uncoded_block[367] ^ uncoded_block[370];
  wire _13094 = uncoded_block[372] ^ uncoded_block[373];
  wire _13095 = _13093 ^ _13094;
  wire _13096 = _13092 ^ _13095;
  wire _13097 = _13091 ^ _13096;
  wire _13098 = _13087 ^ _13097;
  wire _13099 = _13079 ^ _13098;
  wire _13100 = _1036 ^ _7474;
  wire _13101 = uncoded_block[380] ^ uncoded_block[383];
  wire _13102 = uncoded_block[386] ^ uncoded_block[389];
  wire _13103 = _13101 ^ _13102;
  wire _13104 = _13100 ^ _13103;
  wire _13105 = _2615 ^ _1849;
  wire _13106 = uncoded_block[406] ^ uncoded_block[408];
  wire _13107 = _2625 ^ _13106;
  wire _13108 = _13105 ^ _13107;
  wire _13109 = _13104 ^ _13108;
  wire _13110 = uncoded_block[412] ^ uncoded_block[416];
  wire _13111 = _2629 ^ _13110;
  wire _13112 = uncoded_block[417] ^ uncoded_block[418];
  wire _13113 = _13112 ^ _2633;
  wire _13114 = _13111 ^ _13113;
  wire _13115 = uncoded_block[429] ^ uncoded_block[431];
  wire _13116 = _2637 ^ _13115;
  wire _13117 = uncoded_block[433] ^ uncoded_block[437];
  wire _13118 = _13117 ^ _2641;
  wire _13119 = _13116 ^ _13118;
  wire _13120 = _13114 ^ _13119;
  wire _13121 = _13109 ^ _13120;
  wire _13122 = uncoded_block[443] ^ uncoded_block[446];
  wire _13123 = _205 ^ _13122;
  wire _13124 = uncoded_block[452] ^ uncoded_block[456];
  wire _13125 = _1866 ^ _13124;
  wire _13126 = _13123 ^ _13125;
  wire _13127 = uncoded_block[458] ^ uncoded_block[461];
  wire _13128 = _13127 ^ _4890;
  wire _13129 = _3416 ^ _8686;
  wire _13130 = _13128 ^ _13129;
  wire _13131 = _13126 ^ _13130;
  wire _13132 = uncoded_block[475] ^ uncoded_block[478];
  wire _13133 = _1083 ^ _13132;
  wire _13134 = uncoded_block[479] ^ uncoded_block[484];
  wire _13135 = uncoded_block[485] ^ uncoded_block[488];
  wire _13136 = _13134 ^ _13135;
  wire _13137 = _13133 ^ _13136;
  wire _13138 = _10370 ^ _1093;
  wire _13139 = uncoded_block[496] ^ uncoded_block[497];
  wire _13140 = _13139 ^ _4905;
  wire _13141 = _13138 ^ _13140;
  wire _13142 = _13137 ^ _13141;
  wire _13143 = _13131 ^ _13142;
  wire _13144 = _13121 ^ _13143;
  wire _13145 = _13099 ^ _13144;
  wire _13146 = _13061 ^ _13145;
  wire _13147 = _5606 ^ _1892;
  wire _13148 = uncoded_block[511] ^ uncoded_block[514];
  wire _13149 = _3437 ^ _13148;
  wire _13150 = _13147 ^ _13149;
  wire _13151 = _8706 ^ _1895;
  wire _13152 = uncoded_block[520] ^ uncoded_block[524];
  wire _13153 = _13152 ^ _9301;
  wire _13154 = _13151 ^ _13153;
  wire _13155 = _13150 ^ _13154;
  wire _13156 = _1115 ^ _1908;
  wire _13157 = _9310 ^ _13156;
  wire _13158 = _1909 ^ _12592;
  wire _13159 = uncoded_block[551] ^ uncoded_block[554];
  wire _13160 = _13159 ^ _8724;
  wire _13161 = _13158 ^ _13160;
  wire _13162 = _13157 ^ _13161;
  wire _13163 = _13155 ^ _13162;
  wire _13164 = _1924 ^ _3465;
  wire _13165 = uncoded_block[568] ^ uncoded_block[570];
  wire _13166 = _3467 ^ _13165;
  wire _13167 = _13164 ^ _13166;
  wire _13168 = uncoded_block[571] ^ uncoded_block[575];
  wire _13169 = _13168 ^ _10400;
  wire _13170 = _9325 ^ _1139;
  wire _13171 = _13169 ^ _13170;
  wire _13172 = _13167 ^ _13171;
  wire _13173 = _4233 ^ _9330;
  wire _13174 = _8149 ^ _9332;
  wire _13175 = _13173 ^ _13174;
  wire _13176 = uncoded_block[609] ^ uncoded_block[613];
  wire _13177 = _11535 ^ _13176;
  wire _13178 = uncoded_block[615] ^ uncoded_block[618];
  wire _13179 = _13178 ^ _3495;
  wire _13180 = _13177 ^ _13179;
  wire _13181 = _13175 ^ _13180;
  wire _13182 = _13172 ^ _13181;
  wire _13183 = _13163 ^ _13182;
  wire _13184 = uncoded_block[630] ^ uncoded_block[642];
  wire _13185 = _12618 ^ _13184;
  wire _13186 = _13185 ^ _9345;
  wire _13187 = uncoded_block[650] ^ uncoded_block[655];
  wire _13188 = uncoded_block[656] ^ uncoded_block[660];
  wire _13189 = _13187 ^ _13188;
  wire _13190 = uncoded_block[667] ^ uncoded_block[670];
  wire _13191 = _13190 ^ _6353;
  wire _13192 = _13189 ^ _13191;
  wire _13193 = _13186 ^ _13192;
  wire _13194 = uncoded_block[684] ^ uncoded_block[686];
  wire _13195 = _13194 ^ _4271;
  wire _13196 = _326 ^ _8186;
  wire _13197 = _13195 ^ _13196;
  wire _13198 = uncoded_block[697] ^ uncoded_block[704];
  wire _13199 = _13198 ^ _4998;
  wire _13200 = uncoded_block[718] ^ uncoded_block[723];
  wire _13201 = _13200 ^ _3544;
  wire _13202 = _13199 ^ _13201;
  wire _13203 = _13197 ^ _13202;
  wire _13204 = _13193 ^ _13203;
  wire _13205 = _344 ^ _1991;
  wire _13206 = _3547 ^ _8204;
  wire _13207 = _13205 ^ _13206;
  wire _13208 = uncoded_block[740] ^ uncoded_block[743];
  wire _13209 = _13208 ^ _2775;
  wire _13210 = _4293 ^ _5016;
  wire _13211 = _13209 ^ _13210;
  wire _13212 = _13207 ^ _13211;
  wire _13213 = uncoded_block[757] ^ uncoded_block[762];
  wire _13214 = _13213 ^ _1217;
  wire _13215 = uncoded_block[767] ^ uncoded_block[770];
  wire _13216 = uncoded_block[773] ^ uncoded_block[774];
  wire _13217 = _13215 ^ _13216;
  wire _13218 = _13214 ^ _13217;
  wire _13219 = uncoded_block[779] ^ uncoded_block[780];
  wire _13220 = _2014 ^ _13219;
  wire _13221 = _2794 ^ _4309;
  wire _13222 = _13220 ^ _13221;
  wire _13223 = _13218 ^ _13222;
  wire _13224 = _13212 ^ _13223;
  wire _13225 = _13204 ^ _13224;
  wire _13226 = _13183 ^ _13225;
  wire _13227 = _1232 ^ _9928;
  wire _13228 = _373 ^ _13227;
  wire _13229 = _1238 ^ _8228;
  wire _13230 = _2806 ^ _7634;
  wire _13231 = _13229 ^ _13230;
  wire _13232 = _13228 ^ _13231;
  wire _13233 = _1246 ^ _12135;
  wire _13234 = uncoded_block[832] ^ uncoded_block[837];
  wire _13235 = _3590 ^ _13234;
  wire _13236 = _13233 ^ _13235;
  wire _13237 = _4337 ^ _5737;
  wire _13238 = uncoded_block[846] ^ uncoded_block[849];
  wire _13239 = _1256 ^ _13238;
  wire _13240 = _13237 ^ _13239;
  wire _13241 = _13236 ^ _13240;
  wire _13242 = _13232 ^ _13241;
  wire _13243 = _2821 ^ _2046;
  wire _13244 = uncoded_block[861] ^ uncoded_block[864];
  wire _13245 = _408 ^ _13244;
  wire _13246 = _13243 ^ _13245;
  wire _13247 = _414 ^ _5072;
  wire _13248 = _1269 ^ _3608;
  wire _13249 = _13247 ^ _13248;
  wire _13250 = _13246 ^ _13249;
  wire _13251 = uncoded_block[894] ^ uncoded_block[897];
  wire _13252 = _2061 ^ _13251;
  wire _13253 = _6424 ^ _2065;
  wire _13254 = _13252 ^ _13253;
  wire _13255 = _1281 ^ _11067;
  wire _13256 = _5092 ^ _3631;
  wire _13257 = _13255 ^ _13256;
  wire _13258 = _13254 ^ _13257;
  wire _13259 = _13250 ^ _13258;
  wire _13260 = _13242 ^ _13259;
  wire _13261 = uncoded_block[923] ^ uncoded_block[928];
  wire _13262 = _13261 ^ _8835;
  wire _13263 = uncoded_block[942] ^ uncoded_block[944];
  wire _13264 = _9971 ^ _13263;
  wire _13265 = _13262 ^ _13264;
  wire _13266 = uncoded_block[949] ^ uncoded_block[950];
  wire _13267 = _9975 ^ _13266;
  wire _13268 = _7086 ^ _7682;
  wire _13269 = _13267 ^ _13268;
  wire _13270 = _13265 ^ _13269;
  wire _13271 = _1314 ^ _2877;
  wire _13272 = uncoded_block[974] ^ uncoded_block[979];
  wire _13273 = _13272 ^ _5790;
  wire _13274 = _13271 ^ _13273;
  wire _13275 = uncoded_block[982] ^ uncoded_block[991];
  wire _13276 = _13275 ^ _4401;
  wire _13277 = uncoded_block[996] ^ uncoded_block[997];
  wire _13278 = _479 ^ _13277;
  wire _13279 = _13276 ^ _13278;
  wire _13280 = _13274 ^ _13279;
  wire _13281 = _13270 ^ _13280;
  wire _13282 = uncoded_block[1006] ^ uncoded_block[1009];
  wire _13283 = uncoded_block[1010] ^ uncoded_block[1011];
  wire _13284 = _13282 ^ _13283;
  wire _13285 = _2113 ^ _13284;
  wire _13286 = uncoded_block[1019] ^ uncoded_block[1026];
  wire _13287 = _10547 ^ _13286;
  wire _13288 = uncoded_block[1028] ^ uncoded_block[1030];
  wire _13289 = _13288 ^ _4418;
  wire _13290 = _13287 ^ _13289;
  wire _13291 = _13285 ^ _13290;
  wire _13292 = _6474 ^ _6478;
  wire _13293 = _514 ^ _3681;
  wire _13294 = _13292 ^ _13293;
  wire _13295 = uncoded_block[1053] ^ uncoded_block[1055];
  wire _13296 = _9464 ^ _13295;
  wire _13297 = uncoded_block[1058] ^ uncoded_block[1063];
  wire _13298 = _519 ^ _13297;
  wire _13299 = _13296 ^ _13298;
  wire _13300 = _13294 ^ _13299;
  wire _13301 = _13291 ^ _13300;
  wire _13302 = _13281 ^ _13301;
  wire _13303 = _13260 ^ _13302;
  wire _13304 = _13226 ^ _13303;
  wire _13305 = _13146 ^ _13304;
  wire _13306 = _9475 ^ _5156;
  wire _13307 = uncoded_block[1074] ^ uncoded_block[1077];
  wire _13308 = _5158 ^ _13307;
  wire _13309 = _13306 ^ _13308;
  wire _13310 = uncoded_block[1078] ^ uncoded_block[1085];
  wire _13311 = uncoded_block[1087] ^ uncoded_block[1089];
  wire _13312 = _13310 ^ _13311;
  wire _13313 = _5840 ^ _10026;
  wire _13314 = _13312 ^ _13313;
  wire _13315 = _13309 ^ _13314;
  wire _13316 = uncoded_block[1098] ^ uncoded_block[1101];
  wire _13317 = _13316 ^ _2160;
  wire _13318 = uncoded_block[1105] ^ uncoded_block[1107];
  wire _13319 = uncoded_block[1109] ^ uncoded_block[1112];
  wire _13320 = _13318 ^ _13319;
  wire _13321 = _13317 ^ _13320;
  wire _13322 = uncoded_block[1116] ^ uncoded_block[1117];
  wire _13323 = _12782 ^ _13322;
  wire _13324 = _13323 ^ _11698;
  wire _13325 = _13321 ^ _13324;
  wire _13326 = _13315 ^ _13325;
  wire _13327 = uncoded_block[1124] ^ uncoded_block[1127];
  wire _13328 = _13327 ^ _6499;
  wire _13329 = _13328 ^ _562;
  wire _13330 = _564 ^ _8930;
  wire _13331 = _2179 ^ _5862;
  wire _13332 = _13330 ^ _13331;
  wire _13333 = _13329 ^ _13332;
  wire _13334 = _7143 ^ _5188;
  wire _13335 = uncoded_block[1164] ^ uncoded_block[1166];
  wire _13336 = _10043 ^ _13335;
  wire _13337 = _13334 ^ _13336;
  wire _13338 = uncoded_block[1167] ^ uncoded_block[1172];
  wire _13339 = uncoded_block[1174] ^ uncoded_block[1176];
  wire _13340 = _13338 ^ _13339;
  wire _13341 = _8944 ^ _3746;
  wire _13342 = _13340 ^ _13341;
  wire _13343 = _13337 ^ _13342;
  wire _13344 = _13333 ^ _13343;
  wire _13345 = _13326 ^ _13344;
  wire _13346 = uncoded_block[1188] ^ uncoded_block[1191];
  wire _13347 = uncoded_block[1192] ^ uncoded_block[1196];
  wire _13348 = _13346 ^ _13347;
  wire _13349 = uncoded_block[1201] ^ uncoded_block[1205];
  wire _13350 = _7758 ^ _13349;
  wire _13351 = _13348 ^ _13350;
  wire _13352 = _3762 ^ _605;
  wire _13353 = _2218 ^ _13352;
  wire _13354 = _13351 ^ _13353;
  wire _13355 = uncoded_block[1221] ^ uncoded_block[1224];
  wire _13356 = _4499 ^ _13355;
  wire _13357 = uncoded_block[1228] ^ uncoded_block[1229];
  wire _13358 = _612 ^ _13357;
  wire _13359 = _13356 ^ _13358;
  wire _13360 = uncoded_block[1234] ^ uncoded_block[1237];
  wire _13361 = _2225 ^ _13360;
  wire _13362 = _13361 ^ _9527;
  wire _13363 = _13359 ^ _13362;
  wire _13364 = _13354 ^ _13363;
  wire _13365 = uncoded_block[1244] ^ uncoded_block[1246];
  wire _13366 = _13365 ^ _1451;
  wire _13367 = _8385 ^ _5231;
  wire _13368 = _13366 ^ _13367;
  wire _13369 = uncoded_block[1258] ^ uncoded_block[1262];
  wire _13370 = _3001 ^ _13369;
  wire _13371 = _4516 ^ _2239;
  wire _13372 = _13370 ^ _13371;
  wire _13373 = _13368 ^ _13372;
  wire _13374 = uncoded_block[1270] ^ uncoded_block[1273];
  wire _13375 = _13374 ^ _1463;
  wire _13376 = _5908 ^ _12834;
  wire _13377 = _13375 ^ _13376;
  wire _13378 = uncoded_block[1284] ^ uncoded_block[1287];
  wire _13379 = _6557 ^ _13378;
  wire _13380 = uncoded_block[1288] ^ uncoded_block[1289];
  wire _13381 = _13380 ^ _1468;
  wire _13382 = _13379 ^ _13381;
  wire _13383 = _13377 ^ _13382;
  wire _13384 = _13373 ^ _13383;
  wire _13385 = _13364 ^ _13384;
  wire _13386 = _13345 ^ _13385;
  wire _13387 = _10646 ^ _3015;
  wire _13388 = uncoded_block[1299] ^ uncoded_block[1303];
  wire _13389 = _3017 ^ _13388;
  wire _13390 = _13387 ^ _13389;
  wire _13391 = _3025 ^ _1480;
  wire _13392 = _3026 ^ _654;
  wire _13393 = _13391 ^ _13392;
  wire _13394 = _13390 ^ _13393;
  wire _13395 = uncoded_block[1323] ^ uncoded_block[1326];
  wire _13396 = _13395 ^ _10655;
  wire _13397 = _1494 ^ _661;
  wire _13398 = _13396 ^ _13397;
  wire _13399 = uncoded_block[1338] ^ uncoded_block[1339];
  wire _13400 = _13399 ^ _11215;
  wire _13401 = uncoded_block[1349] ^ uncoded_block[1352];
  wire _13402 = _664 ^ _13401;
  wire _13403 = _13400 ^ _13402;
  wire _13404 = _13398 ^ _13403;
  wire _13405 = _13394 ^ _13404;
  wire _13406 = _5272 ^ _3045;
  wire _13407 = uncoded_block[1363] ^ uncoded_block[1367];
  wire _13408 = _13407 ^ _3052;
  wire _13409 = _13406 ^ _13408;
  wire _13410 = uncoded_block[1379] ^ uncoded_block[1382];
  wire _13411 = _10103 ^ _13410;
  wire _13412 = uncoded_block[1390] ^ uncoded_block[1391];
  wire _13413 = _10108 ^ _13412;
  wire _13414 = _13411 ^ _13413;
  wire _13415 = _13409 ^ _13414;
  wire _13416 = uncoded_block[1394] ^ uncoded_block[1397];
  wire _13417 = _13416 ^ _4572;
  wire _13418 = _2297 ^ _3846;
  wire _13419 = _13417 ^ _13418;
  wire _13420 = uncoded_block[1406] ^ uncoded_block[1409];
  wire _13421 = _13420 ^ _12877;
  wire _13422 = uncoded_block[1414] ^ uncoded_block[1415];
  wire _13423 = _13422 ^ _10118;
  wire _13424 = _13421 ^ _13423;
  wire _13425 = _13419 ^ _13424;
  wire _13426 = _13415 ^ _13425;
  wire _13427 = _13405 ^ _13426;
  wire _13428 = uncoded_block[1419] ^ uncoded_block[1422];
  wire _13429 = uncoded_block[1424] ^ uncoded_block[1426];
  wire _13430 = _13428 ^ _13429;
  wire _13431 = _13430 ^ _9592;
  wire _13432 = uncoded_block[1438] ^ uncoded_block[1440];
  wire _13433 = _10690 ^ _13432;
  wire _13434 = _13433 ^ _4592;
  wire _13435 = _13431 ^ _13434;
  wire _13436 = _3865 ^ _2326;
  wire _13437 = uncoded_block[1457] ^ uncoded_block[1459];
  wire _13438 = _5309 ^ _13437;
  wire _13439 = _13436 ^ _13438;
  wire _13440 = uncoded_block[1460] ^ uncoded_block[1464];
  wire _13441 = _13440 ^ _10136;
  wire _13442 = _7247 ^ _1551;
  wire _13443 = _13441 ^ _13442;
  wire _13444 = _13439 ^ _13443;
  wire _13445 = _13435 ^ _13444;
  wire _13446 = uncoded_block[1477] ^ uncoded_block[1479];
  wire _13447 = _4603 ^ _13446;
  wire _13448 = uncoded_block[1481] ^ uncoded_block[1482];
  wire _13449 = _13448 ^ _5320;
  wire _13450 = _13447 ^ _13449;
  wire _13451 = _2349 ^ _1563;
  wire _13452 = uncoded_block[1497] ^ uncoded_block[1501];
  wire _13453 = _2350 ^ _13452;
  wire _13454 = _13451 ^ _13453;
  wire _13455 = _13450 ^ _13454;
  wire _13456 = _5333 ^ _9620;
  wire _13457 = _5331 ^ _13456;
  wire _13458 = uncoded_block[1516] ^ uncoded_block[1521];
  wire _13459 = uncoded_block[1526] ^ uncoded_block[1528];
  wire _13460 = _13458 ^ _13459;
  wire _13461 = _5344 ^ _12914;
  wire _13462 = _13460 ^ _13461;
  wire _13463 = _13457 ^ _13462;
  wire _13464 = _13455 ^ _13463;
  wire _13465 = _13445 ^ _13464;
  wire _13466 = _13427 ^ _13465;
  wire _13467 = _13386 ^ _13466;
  wire _13468 = _6006 ^ _6651;
  wire _13469 = _6008 ^ _5355;
  wire _13470 = _13468 ^ _13469;
  wire _13471 = uncoded_block[1547] ^ uncoded_block[1548];
  wire _13472 = uncoded_block[1549] ^ uncoded_block[1550];
  wire _13473 = _13471 ^ _13472;
  wire _13474 = _13473 ^ _6658;
  wire _13475 = _13470 ^ _13474;
  wire _13476 = _10160 ^ _2372;
  wire _13477 = _13476 ^ _12367;
  wire _13478 = uncoded_block[1573] ^ uncoded_block[1575];
  wire _13479 = uncoded_block[1578] ^ uncoded_block[1580];
  wire _13480 = _13478 ^ _13479;
  wire _13481 = _6031 ^ _2386;
  wire _13482 = _13480 ^ _13481;
  wire _13483 = _13477 ^ _13482;
  wire _13484 = _13475 ^ _13483;
  wire _13485 = _789 ^ _2394;
  wire _13486 = uncoded_block[1596] ^ uncoded_block[1597];
  wire _13487 = _13486 ^ _6039;
  wire _13488 = _13485 ^ _13487;
  wire _13489 = _4660 ^ _5380;
  wire _13490 = uncoded_block[1611] ^ uncoded_block[1615];
  wire _13491 = _13490 ^ _804;
  wire _13492 = _13489 ^ _13491;
  wire _13493 = _13488 ^ _13492;
  wire _13494 = uncoded_block[1623] ^ uncoded_block[1625];
  wire _13495 = _3160 ^ _13494;
  wire _13496 = uncoded_block[1629] ^ uncoded_block[1633];
  wire _13497 = _3942 ^ _13496;
  wire _13498 = _13495 ^ _13497;
  wire _13499 = _11858 ^ _6689;
  wire _13500 = uncoded_block[1642] ^ uncoded_block[1643];
  wire _13501 = _13500 ^ _7312;
  wire _13502 = _13499 ^ _13501;
  wire _13503 = _13498 ^ _13502;
  wire _13504 = _13493 ^ _13503;
  wire _13505 = _13484 ^ _13504;
  wire _13506 = uncoded_block[1651] ^ uncoded_block[1655];
  wire _13507 = _9661 ^ _13506;
  wire _13508 = uncoded_block[1656] ^ uncoded_block[1658];
  wire _13509 = _13508 ^ _3958;
  wire _13510 = _13507 ^ _13509;
  wire _13511 = uncoded_block[1664] ^ uncoded_block[1667];
  wire _13512 = _13511 ^ _7928;
  wire _13513 = uncoded_block[1674] ^ uncoded_block[1677];
  wire _13514 = _6700 ^ _13513;
  wire _13515 = _13512 ^ _13514;
  wire _13516 = _13510 ^ _13515;
  wire _13517 = uncoded_block[1681] ^ uncoded_block[1683];
  wire _13518 = _11321 ^ _13517;
  wire _13519 = uncoded_block[1687] ^ uncoded_block[1689];
  wire _13520 = _13519 ^ _7331;
  wire _13521 = _13518 ^ _13520;
  wire _13522 = uncoded_block[1692] ^ uncoded_block[1697];
  wire _13523 = _13522 ^ _2434;
  wire _13524 = _848 ^ _12407;
  wire _13525 = _13523 ^ _13524;
  wire _13526 = _13521 ^ _13525;
  wire _13527 = _13516 ^ _13526;
  wire _13528 = uncoded_block[1716] ^ uncoded_block[1719];
  wire _13529 = _13528 ^ uncoded_block[1720];
  wire _13530 = _13527 ^ _13529;
  wire _13531 = _13505 ^ _13530;
  wire _13532 = _13467 ^ _13531;
  wire _13533 = _13305 ^ _13532;
  wire _13534 = _10223 ^ _3993;
  wire _13535 = _3213 ^ _6086;
  wire _13536 = _13534 ^ _13535;
  wire _13537 = uncoded_block[18] ^ uncoded_block[20];
  wire _13538 = _871 ^ _13537;
  wire _13539 = uncoded_block[25] ^ uncoded_block[27];
  wire _13540 = _10 ^ _13539;
  wire _13541 = _13538 ^ _13540;
  wire _13542 = _13536 ^ _13541;
  wire _13543 = uncoded_block[31] ^ uncoded_block[34];
  wire _13544 = _13543 ^ _8549;
  wire _13545 = _13544 ^ _2467;
  wire _13546 = _22 ^ _8554;
  wire _13547 = uncoded_block[50] ^ uncoded_block[52];
  wire _13548 = _13547 ^ _25;
  wire _13549 = _13546 ^ _13548;
  wire _13550 = _13545 ^ _13549;
  wire _13551 = _13542 ^ _13550;
  wire _13552 = uncoded_block[57] ^ uncoded_block[60];
  wire _13553 = uncoded_block[61] ^ uncoded_block[62];
  wire _13554 = _13552 ^ _13553;
  wire _13555 = _6744 ^ _3241;
  wire _13556 = _13554 ^ _13555;
  wire _13557 = _1712 ^ _901;
  wire _13558 = uncoded_block[82] ^ uncoded_block[84];
  wire _13559 = _13558 ^ _2484;
  wire _13560 = _13557 ^ _13559;
  wire _13561 = _13556 ^ _13560;
  wire _13562 = _9713 ^ _1718;
  wire _13563 = _4026 ^ _47;
  wire _13564 = _13562 ^ _13563;
  wire _13565 = _910 ^ _13010;
  wire _13566 = _6123 ^ _7990;
  wire _13567 = _13565 ^ _13566;
  wire _13568 = _13564 ^ _13567;
  wire _13569 = _13561 ^ _13568;
  wire _13570 = _13551 ^ _13569;
  wire _13571 = uncoded_block[118] ^ uncoded_block[122];
  wire _13572 = _13571 ^ _9727;
  wire _13573 = uncoded_block[144] ^ uncoded_block[148];
  wire _13574 = _926 ^ _13573;
  wire _13575 = _13572 ^ _13574;
  wire _13576 = _1744 ^ _3271;
  wire _13577 = _4049 ^ _6144;
  wire _13578 = _13576 ^ _13577;
  wire _13579 = _13575 ^ _13578;
  wire _13580 = _1749 ^ _4056;
  wire _13581 = _13580 ^ _8008;
  wire _13582 = _940 ^ _4770;
  wire _13583 = uncoded_block[182] ^ uncoded_block[183];
  wire _13584 = _13583 ^ _4062;
  wire _13585 = _13582 ^ _13584;
  wire _13586 = _13581 ^ _13585;
  wire _13587 = _13579 ^ _13586;
  wire _13588 = uncoded_block[188] ^ uncoded_block[189];
  wire _13589 = _13588 ^ _5483;
  wire _13590 = uncoded_block[195] ^ uncoded_block[199];
  wire _13591 = _4776 ^ _13590;
  wire _13592 = _13589 ^ _13591;
  wire _13593 = _10849 ^ _4780;
  wire _13594 = _955 ^ _1767;
  wire _13595 = _13593 ^ _13594;
  wire _13596 = _13592 ^ _13595;
  wire _13597 = uncoded_block[221] ^ uncoded_block[224];
  wire _13598 = _102 ^ _13597;
  wire _13599 = _10287 ^ _7422;
  wire _13600 = _13598 ^ _13599;
  wire _13601 = _1780 ^ _8616;
  wire _13602 = _11949 ^ _13601;
  wire _13603 = _13600 ^ _13602;
  wire _13604 = _13596 ^ _13603;
  wire _13605 = _13587 ^ _13604;
  wire _13606 = _13570 ^ _13605;
  wire _13607 = _3309 ^ _3311;
  wire _13608 = _11955 ^ _13607;
  wire _13609 = uncoded_block[258] ^ uncoded_block[261];
  wire _13610 = _13609 ^ _2568;
  wire _13611 = _5515 ^ _6197;
  wire _13612 = _13610 ^ _13611;
  wire _13613 = _13608 ^ _13612;
  wire _13614 = _1804 ^ _4819;
  wire _13615 = uncoded_block[295] ^ uncoded_block[298];
  wire _13616 = _13615 ^ _142;
  wire _13617 = _13614 ^ _13616;
  wire _13618 = _4826 ^ _6845;
  wire _13619 = uncoded_block[310] ^ uncoded_block[313];
  wire _13620 = _3334 ^ _13619;
  wire _13621 = _13618 ^ _13620;
  wire _13622 = _13617 ^ _13621;
  wire _13623 = _13613 ^ _13622;
  wire _13624 = uncoded_block[316] ^ uncoded_block[319];
  wire _13625 = uncoded_block[321] ^ uncoded_block[323];
  wire _13626 = _13624 ^ _13625;
  wire _13627 = _8058 ^ _2586;
  wire _13628 = _13626 ^ _13627;
  wire _13629 = uncoded_block[335] ^ uncoded_block[338];
  wire _13630 = _1821 ^ _13629;
  wire _13631 = _9242 ^ _3355;
  wire _13632 = _13630 ^ _13631;
  wire _13633 = _13628 ^ _13632;
  wire _13634 = _10892 ^ _2603;
  wire _13635 = _6227 ^ _11463;
  wire _13636 = _1835 ^ _8076;
  wire _13637 = _13635 ^ _13636;
  wire _13638 = _13634 ^ _13637;
  wire _13639 = _13633 ^ _13638;
  wire _13640 = _13623 ^ _13639;
  wire _13641 = _10334 ^ _4143;
  wire _13642 = _1038 ^ _11999;
  wire _13643 = _13641 ^ _13642;
  wire _13644 = uncoded_block[387] ^ uncoded_block[392];
  wire _13645 = _13644 ^ _6881;
  wire _13646 = uncoded_block[401] ^ uncoded_block[403];
  wire _13647 = _2622 ^ _13646;
  wire _13648 = _13645 ^ _13647;
  wire _13649 = _13643 ^ _13648;
  wire _13650 = uncoded_block[412] ^ uncoded_block[415];
  wire _13651 = _2626 ^ _13650;
  wire _13652 = uncoded_block[424] ^ uncoded_block[429];
  wire _13653 = _11477 ^ _13652;
  wire _13654 = _13651 ^ _13653;
  wire _13655 = uncoded_block[431] ^ uncoded_block[435];
  wire _13656 = _13655 ^ _4169;
  wire _13657 = _1863 ^ _7498;
  wire _13658 = _13656 ^ _13657;
  wire _13659 = _13654 ^ _13658;
  wire _13660 = _13649 ^ _13659;
  wire _13661 = _1866 ^ _2645;
  wire _13662 = uncoded_block[462] ^ uncoded_block[463];
  wire _13663 = _10926 ^ _13662;
  wire _13664 = _13661 ^ _13663;
  wire _13665 = uncoded_block[467] ^ uncoded_block[471];
  wire _13666 = _8683 ^ _13665;
  wire _13667 = _13666 ^ _5591;
  wire _13668 = _13664 ^ _13667;
  wire _13669 = uncoded_block[485] ^ uncoded_block[491];
  wire _13670 = _7513 ^ _13669;
  wire _13671 = uncoded_block[495] ^ uncoded_block[502];
  wire _13672 = _3432 ^ _13671;
  wire _13673 = _13670 ^ _13672;
  wire _13674 = uncoded_block[505] ^ uncoded_block[509];
  wire _13675 = _6921 ^ _13674;
  wire _13676 = uncoded_block[513] ^ uncoded_block[514];
  wire _13677 = _4908 ^ _13676;
  wire _13678 = _13675 ^ _13677;
  wire _13679 = _13673 ^ _13678;
  wire _13680 = _13668 ^ _13679;
  wire _13681 = _13660 ^ _13680;
  wire _13682 = _13640 ^ _13681;
  wire _13683 = _13606 ^ _13682;
  wire _13684 = uncoded_block[524] ^ uncoded_block[525];
  wire _13685 = _9299 ^ _13684;
  wire _13686 = _6929 ^ _10384;
  wire _13687 = _13685 ^ _13686;
  wire _13688 = uncoded_block[537] ^ uncoded_block[543];
  wire _13689 = uncoded_block[545] ^ uncoded_block[547];
  wire _13690 = _13688 ^ _13689;
  wire _13691 = _1912 ^ _3459;
  wire _13692 = _13690 ^ _13691;
  wire _13693 = _13687 ^ _13692;
  wire _13694 = _8724 ^ _1916;
  wire _13695 = _8139 ^ _3464;
  wire _13696 = _13694 ^ _13695;
  wire _13697 = uncoded_block[567] ^ uncoded_block[569];
  wire _13698 = uncoded_block[571] ^ uncoded_block[573];
  wire _13699 = _13697 ^ _13698;
  wire _13700 = uncoded_block[574] ^ uncoded_block[578];
  wire _13701 = _13700 ^ _6947;
  wire _13702 = _13699 ^ _13701;
  wire _13703 = _13696 ^ _13702;
  wire _13704 = _13693 ^ _13703;
  wire _13705 = uncoded_block[589] ^ uncoded_block[591];
  wire _13706 = _8143 ^ _13705;
  wire _13707 = _3480 ^ _6952;
  wire _13708 = _13706 ^ _13707;
  wire _13709 = _8152 ^ _1942;
  wire _13710 = _3488 ^ _13709;
  wire _13711 = _13708 ^ _13710;
  wire _13712 = _8154 ^ _7564;
  wire _13713 = uncoded_block[616] ^ uncoded_block[617];
  wire _13714 = _13713 ^ _4243;
  wire _13715 = _13712 ^ _13714;
  wire _13716 = _2719 ^ _1154;
  wire _13717 = uncoded_block[634] ^ uncoded_block[638];
  wire _13718 = _12620 ^ _13717;
  wire _13719 = _13716 ^ _13718;
  wire _13720 = _13715 ^ _13719;
  wire _13721 = _13711 ^ _13720;
  wire _13722 = _13704 ^ _13721;
  wire _13723 = _1163 ^ _2729;
  wire _13724 = _6338 ^ _6973;
  wire _13725 = _13723 ^ _13724;
  wire _13726 = uncoded_block[665] ^ uncoded_block[667];
  wire _13727 = _4262 ^ _13726;
  wire _13728 = _306 ^ _13727;
  wire _13729 = _13725 ^ _13728;
  wire _13730 = _311 ^ _1178;
  wire _13731 = uncoded_block[677] ^ uncoded_block[678];
  wire _13732 = _10434 ^ _13731;
  wire _13733 = _13730 ^ _13732;
  wire _13734 = _3522 ^ _2750;
  wire _13735 = uncoded_block[690] ^ uncoded_block[692];
  wire _13736 = _13735 ^ _328;
  wire _13737 = _13734 ^ _13736;
  wire _13738 = _13733 ^ _13737;
  wire _13739 = _13729 ^ _13738;
  wire _13740 = uncoded_block[699] ^ uncoded_block[702];
  wire _13741 = _13740 ^ _5685;
  wire _13742 = uncoded_block[711] ^ uncoded_block[716];
  wire _13743 = _4995 ^ _13742;
  wire _13744 = _13741 ^ _13743;
  wire _13745 = _5002 ^ _6367;
  wire _13746 = _9369 ^ _4283;
  wire _13747 = _13745 ^ _13746;
  wire _13748 = _13744 ^ _13747;
  wire _13749 = uncoded_block[728] ^ uncoded_block[730];
  wire _13750 = _13749 ^ _1991;
  wire _13751 = _13750 ^ _12104;
  wire _13752 = uncoded_block[744] ^ uncoded_block[748];
  wire _13753 = _13752 ^ _1210;
  wire _13754 = uncoded_block[751] ^ uncoded_block[755];
  wire _13755 = _13754 ^ _3559;
  wire _13756 = _13753 ^ _13755;
  wire _13757 = _13751 ^ _13756;
  wire _13758 = _13748 ^ _13757;
  wire _13759 = _13739 ^ _13758;
  wire _13760 = _13722 ^ _13759;
  wire _13761 = uncoded_block[761] ^ uncoded_block[763];
  wire _13762 = uncoded_block[764] ^ uncoded_block[766];
  wire _13763 = _13761 ^ _13762;
  wire _13764 = _5027 ^ _11019;
  wire _13765 = _13763 ^ _13764;
  wire _13766 = uncoded_block[775] ^ uncoded_block[778];
  wire _13767 = _1221 ^ _13766;
  wire _13768 = uncoded_block[779] ^ uncoded_block[783];
  wire _13769 = _13768 ^ _3570;
  wire _13770 = _13767 ^ _13769;
  wire _13771 = _13765 ^ _13770;
  wire _13772 = _3571 ^ _375;
  wire _13773 = _13772 ^ _384;
  wire _13774 = _389 ^ _2026;
  wire _13775 = _387 ^ _13774;
  wire _13776 = _13773 ^ _13775;
  wire _13777 = _13771 ^ _13776;
  wire _13778 = _2808 ^ _2028;
  wire _13779 = _6399 ^ _2812;
  wire _13780 = _13778 ^ _13779;
  wire _13781 = uncoded_block[833] ^ uncoded_block[836];
  wire _13782 = _13781 ^ _11043;
  wire _13783 = uncoded_block[841] ^ uncoded_block[845];
  wire _13784 = _13783 ^ _2820;
  wire _13785 = _13782 ^ _13784;
  wire _13786 = _13780 ^ _13785;
  wire _13787 = _8809 ^ _3600;
  wire _13788 = _5747 ^ _413;
  wire _13789 = _13787 ^ _13788;
  wire _13790 = _414 ^ _7054;
  wire _13791 = uncoded_block[872] ^ uncoded_block[874];
  wire _13792 = _6415 ^ _13791;
  wire _13793 = _13790 ^ _13792;
  wire _13794 = _13789 ^ _13793;
  wire _13795 = _13786 ^ _13794;
  wire _13796 = _13777 ^ _13795;
  wire _13797 = uncoded_block[885] ^ uncoded_block[887];
  wire _13798 = _3608 ^ _13797;
  wire _13799 = uncoded_block[888] ^ uncoded_block[891];
  wire _13800 = _13799 ^ _12704;
  wire _13801 = _13798 ^ _13800;
  wire _13802 = _5758 ^ _429;
  wire _13803 = _9960 ^ _8254;
  wire _13804 = _13802 ^ _13803;
  wire _13805 = _13801 ^ _13804;
  wire _13806 = _1285 ^ _6430;
  wire _13807 = _10513 ^ _2073;
  wire _13808 = _13806 ^ _13807;
  wire _13809 = uncoded_block[931] ^ uncoded_block[937];
  wire _13810 = _13809 ^ _7080;
  wire _13811 = _9426 ^ _13810;
  wire _13812 = _13808 ^ _13811;
  wire _13813 = _13805 ^ _13812;
  wire _13814 = _8271 ^ _9975;
  wire _13815 = _13266 ^ _461;
  wire _13816 = _13814 ^ _13815;
  wire _13817 = _11642 ^ _1308;
  wire _13818 = _13817 ^ _9982;
  wire _13819 = _13816 ^ _13818;
  wire _13820 = _11648 ^ _468;
  wire _13821 = uncoded_block[973] ^ uncoded_block[976];
  wire _13822 = uncoded_block[981] ^ uncoded_block[984];
  wire _13823 = _13821 ^ _13822;
  wire _13824 = _13820 ^ _13823;
  wire _13825 = uncoded_block[985] ^ uncoded_block[990];
  wire _13826 = _13825 ^ _10543;
  wire _13827 = _4402 ^ _1326;
  wire _13828 = _13826 ^ _13827;
  wire _13829 = _13824 ^ _13828;
  wire _13830 = _13819 ^ _13829;
  wire _13831 = _13813 ^ _13830;
  wire _13832 = _13796 ^ _13831;
  wire _13833 = _13760 ^ _13832;
  wire _13834 = _13683 ^ _13833;
  wire _13835 = uncoded_block[1007] ^ uncoded_block[1012];
  wire _13836 = _13835 ^ _2891;
  wire _13837 = uncoded_block[1021] ^ uncoded_block[1025];
  wire _13838 = _13837 ^ _8874;
  wire _13839 = _13836 ^ _13838;
  wire _13840 = _13288 ^ _2127;
  wire _13841 = _13840 ^ _8881;
  wire _13842 = _13839 ^ _13841;
  wire _13843 = uncoded_block[1040] ^ uncoded_block[1045];
  wire _13844 = uncoded_block[1049] ^ uncoded_block[1051];
  wire _13845 = _13843 ^ _13844;
  wire _13846 = uncoded_block[1052] ^ uncoded_block[1056];
  wire _13847 = _13846 ^ _7117;
  wire _13848 = _13845 ^ _13847;
  wire _13849 = uncoded_block[1059] ^ uncoded_block[1062];
  wire _13850 = _13849 ^ _8888;
  wire _13851 = uncoded_block[1068] ^ uncoded_block[1071];
  wire _13852 = _13851 ^ _8895;
  wire _13853 = _13850 ^ _13852;
  wire _13854 = _13848 ^ _13853;
  wire _13855 = _13842 ^ _13854;
  wire _13856 = _5834 ^ _533;
  wire _13857 = uncoded_block[1089] ^ uncoded_block[1092];
  wire _13858 = _3696 ^ _13857;
  wire _13859 = _13856 ^ _13858;
  wire _13860 = _5842 ^ _1380;
  wire _13861 = uncoded_block[1111] ^ uncoded_block[1116];
  wire _13862 = _545 ^ _13861;
  wire _13863 = _13860 ^ _13862;
  wire _13864 = _13859 ^ _13863;
  wire _13865 = _1388 ^ _4455;
  wire _13866 = uncoded_block[1131] ^ uncoded_block[1133];
  wire _13867 = _13327 ^ _13866;
  wire _13868 = _13865 ^ _13867;
  wire _13869 = uncoded_block[1134] ^ uncoded_block[1137];
  wire _13870 = _13869 ^ _565;
  wire _13871 = _13870 ^ _569;
  wire _13872 = _13868 ^ _13871;
  wire _13873 = _13864 ^ _13872;
  wire _13874 = _13855 ^ _13873;
  wire _13875 = _8932 ^ _1401;
  wire _13876 = _4468 ^ _3727;
  wire _13877 = _13875 ^ _13876;
  wire _13878 = _3728 ^ _2958;
  wire _13879 = _13878 ^ _3737;
  wire _13880 = _13877 ^ _13879;
  wire _13881 = _3740 ^ _10608;
  wire _13882 = uncoded_block[1182] ^ uncoded_block[1185];
  wire _13883 = uncoded_block[1186] ^ uncoded_block[1189];
  wire _13884 = _13882 ^ _13883;
  wire _13885 = _13881 ^ _13884;
  wire _13886 = uncoded_block[1196] ^ uncoded_block[1200];
  wire _13887 = _13886 ^ _6529;
  wire _13888 = _8950 ^ _13887;
  wire _13889 = _13885 ^ _13888;
  wire _13890 = _13880 ^ _13889;
  wire _13891 = _6530 ^ _10617;
  wire _13892 = _13891 ^ _13352;
  wire _13893 = uncoded_block[1218] ^ uncoded_block[1223];
  wire _13894 = _13893 ^ _1435;
  wire _13895 = _1436 ^ _5218;
  wire _13896 = _13894 ^ _13895;
  wire _13897 = _13892 ^ _13896;
  wire _13898 = uncoded_block[1233] ^ uncoded_block[1238];
  wire _13899 = _13898 ^ _4509;
  wire _13900 = _11734 ^ _5229;
  wire _13901 = _13899 ^ _13900;
  wire _13902 = _1455 ^ _5234;
  wire _13903 = _13367 ^ _13902;
  wire _13904 = _13901 ^ _13903;
  wire _13905 = _13897 ^ _13904;
  wire _13906 = _13890 ^ _13905;
  wire _13907 = _13874 ^ _13906;
  wire _13908 = _8391 ^ _7179;
  wire _13909 = _10075 ^ _1463;
  wire _13910 = _13908 ^ _13909;
  wire _13911 = _631 ^ _6557;
  wire _13912 = _13378 ^ _13380;
  wire _13913 = _13911 ^ _13912;
  wire _13914 = _13910 ^ _13913;
  wire _13915 = uncoded_block[1298] ^ uncoded_block[1304];
  wire _13916 = _9545 ^ _13915;
  wire _13917 = uncoded_block[1309] ^ uncoded_block[1312];
  wire _13918 = _3025 ^ _13917;
  wire _13919 = _13916 ^ _13918;
  wire _13920 = uncoded_block[1315] ^ uncoded_block[1320];
  wire _13921 = _13920 ^ _3029;
  wire _13922 = uncoded_block[1329] ^ uncoded_block[1332];
  wire _13923 = _8411 ^ _13922;
  wire _13924 = _13921 ^ _13923;
  wire _13925 = _13919 ^ _13924;
  wire _13926 = _13914 ^ _13925;
  wire _13927 = uncoded_block[1341] ^ uncoded_block[1343];
  wire _13928 = _13927 ^ _1498;
  wire _13929 = _13928 ^ _13402;
  wire _13930 = _4558 ^ _5275;
  wire _13931 = _677 ^ _679;
  wire _13932 = _13930 ^ _13931;
  wire _13933 = _13929 ^ _13932;
  wire _13934 = _10668 ^ _8423;
  wire _13935 = _5284 ^ _4564;
  wire _13936 = _13934 ^ _13935;
  wire _13937 = _12311 ^ _6597;
  wire _13938 = uncoded_block[1396] ^ uncoded_block[1397];
  wire _13939 = uncoded_block[1398] ^ uncoded_block[1401];
  wire _13940 = _13938 ^ _13939;
  wire _13941 = _13937 ^ _13940;
  wire _13942 = _13936 ^ _13941;
  wire _13943 = _13933 ^ _13942;
  wire _13944 = _13926 ^ _13943;
  wire _13945 = uncoded_block[1402] ^ uncoded_block[1405];
  wire _13946 = _13945 ^ _701;
  wire _13947 = uncoded_block[1409] ^ uncoded_block[1411];
  wire _13948 = _13947 ^ _5962;
  wire _13949 = _13946 ^ _13948;
  wire _13950 = _7842 ^ _7844;
  wire _13951 = uncoded_block[1431] ^ uncoded_block[1438];
  wire _13952 = _10684 ^ _13951;
  wire _13953 = _13950 ^ _13952;
  wire _13954 = _13949 ^ _13953;
  wire _13955 = _3861 ^ _1541;
  wire _13956 = _13955 ^ _10695;
  wire _13957 = _720 ^ _3870;
  wire _13958 = _10699 ^ _3879;
  wire _13959 = _13957 ^ _13958;
  wire _13960 = _13956 ^ _13959;
  wire _13961 = _13954 ^ _13960;
  wire _13962 = _3097 ^ _1555;
  wire _13963 = uncoded_block[1478] ^ uncoded_block[1481];
  wire _13964 = _13963 ^ _7861;
  wire _13965 = _13962 ^ _13964;
  wire _13966 = uncoded_block[1488] ^ uncoded_block[1491];
  wire _13967 = uncoded_block[1493] ^ uncoded_block[1495];
  wire _13968 = _13966 ^ _13967;
  wire _13969 = uncoded_block[1496] ^ uncoded_block[1502];
  wire _13970 = _13969 ^ _7259;
  wire _13971 = _13968 ^ _13970;
  wire _13972 = _13965 ^ _13971;
  wire _13973 = uncoded_block[1508] ^ uncoded_block[1512];
  wire _13974 = _3112 ^ _13973;
  wire _13975 = uncoded_block[1513] ^ uncoded_block[1519];
  wire _13976 = _13975 ^ _1579;
  wire _13977 = _13974 ^ _13976;
  wire _13978 = uncoded_block[1523] ^ uncoded_block[1528];
  wire _13979 = uncoded_block[1532] ^ uncoded_block[1536];
  wire _13980 = _13978 ^ _13979;
  wire _13981 = _6650 ^ _5350;
  wire _13982 = _13980 ^ _13981;
  wire _13983 = _13977 ^ _13982;
  wire _13984 = _13972 ^ _13983;
  wire _13985 = _13961 ^ _13984;
  wire _13986 = _13944 ^ _13985;
  wire _13987 = _13907 ^ _13986;
  wire _13988 = _6008 ^ _7274;
  wire _13989 = _10157 ^ _10732;
  wire _13990 = _13988 ^ _13989;
  wire _13991 = uncoded_block[1561] ^ uncoded_block[1563];
  wire _13992 = _13991 ^ _9072;
  wire _13993 = _4647 ^ _784;
  wire _13994 = _13992 ^ _13993;
  wire _13995 = _13990 ^ _13994;
  wire _13996 = uncoded_block[1595] ^ uncoded_block[1598];
  wire _13997 = _788 ^ _13996;
  wire _13998 = _1621 ^ _3151;
  wire _13999 = _13997 ^ _13998;
  wire _14000 = uncoded_block[1604] ^ uncoded_block[1608];
  wire _14001 = _14000 ^ _801;
  wire _14002 = _10181 ^ _7911;
  wire _14003 = _14001 ^ _14002;
  wire _14004 = _13999 ^ _14003;
  wire _14005 = _13995 ^ _14004;
  wire _14006 = uncoded_block[1625] ^ uncoded_block[1628];
  wire _14007 = _7300 ^ _14006;
  wire _14008 = _14007 ^ _5389;
  wire _14009 = uncoded_block[1636] ^ uncoded_block[1642];
  wire _14010 = _14009 ^ _4673;
  wire _14011 = uncoded_block[1654] ^ uncoded_block[1655];
  wire _14012 = _3953 ^ _14011;
  wire _14013 = _14010 ^ _14012;
  wire _14014 = _14008 ^ _14013;
  wire _14015 = _12390 ^ _1653;
  wire _14016 = _7927 ^ _4687;
  wire _14017 = _14015 ^ _14016;
  wire _14018 = _7323 ^ _12398;
  wire _14019 = _10766 ^ _4693;
  wire _14020 = _14018 ^ _14019;
  wire _14021 = _14017 ^ _14020;
  wire _14022 = _14014 ^ _14021;
  wire _14023 = _14005 ^ _14022;
  wire _14024 = uncoded_block[1692] ^ uncoded_block[1695];
  wire _14025 = uncoded_block[1697] ^ uncoded_block[1701];
  wire _14026 = _14024 ^ _14025;
  wire _14027 = _9671 ^ _14026;
  wire _14028 = uncoded_block[1703] ^ uncoded_block[1706];
  wire _14029 = _14028 ^ _10778;
  wire _14030 = _854 ^ _1677;
  wire _14031 = _14029 ^ _14030;
  wire _14032 = _14027 ^ _14031;
  wire _14033 = _3988 ^ uncoded_block[1720];
  wire _14034 = _14032 ^ _14033;
  wire _14035 = _14023 ^ _14034;
  wire _14036 = _13987 ^ _14035;
  wire _14037 = _13834 ^ _14036;
  wire _14038 = uncoded_block[4] ^ uncoded_block[8];
  wire _14039 = _4710 ^ _14038;
  wire _14040 = _14039 ^ _10789;
  wire _14041 = _3998 ^ _10226;
  wire _14042 = _4000 ^ _13539;
  wire _14043 = _14041 ^ _14042;
  wire _14044 = _14040 ^ _14043;
  wire _14045 = _6095 ^ _8549;
  wire _14046 = _876 ^ _14045;
  wire _14047 = uncoded_block[38] ^ uncoded_block[41];
  wire _14048 = uncoded_block[42] ^ uncoded_block[47];
  wire _14049 = _14047 ^ _14048;
  wire _14050 = _9150 ^ _4014;
  wire _14051 = _14049 ^ _14050;
  wire _14052 = _14046 ^ _14051;
  wire _14053 = _14044 ^ _14052;
  wire _14054 = _5436 ^ _7364;
  wire _14055 = uncoded_block[63] ^ uncoded_block[66];
  wire _14056 = _14055 ^ _11357;
  wire _14057 = _14054 ^ _14056;
  wire _14058 = uncoded_block[72] ^ uncoded_block[74];
  wire _14059 = _7976 ^ _14058;
  wire _14060 = uncoded_block[76] ^ uncoded_block[78];
  wire _14061 = _14060 ^ _6749;
  wire _14062 = _14059 ^ _14061;
  wire _14063 = _14057 ^ _14062;
  wire _14064 = _6750 ^ _6754;
  wire _14065 = uncoded_block[87] ^ uncoded_block[89];
  wire _14066 = _14065 ^ _9715;
  wire _14067 = _14064 ^ _14066;
  wire _14068 = uncoded_block[96] ^ uncoded_block[97];
  wire _14069 = _14068 ^ _9718;
  wire _14070 = _14069 ^ _6121;
  wire _14071 = _14067 ^ _14070;
  wire _14072 = _14063 ^ _14071;
  wire _14073 = _14053 ^ _14072;
  wire _14074 = uncoded_block[115] ^ uncoded_block[119];
  wire _14075 = _6123 ^ _14074;
  wire _14076 = _10256 ^ _1730;
  wire _14077 = _14075 ^ _14076;
  wire _14078 = _3263 ^ _64;
  wire _14079 = _12458 ^ _14078;
  wire _14080 = _14077 ^ _14079;
  wire _14081 = _7392 ^ _4046;
  wire _14082 = uncoded_block[148] ^ uncoded_block[149];
  wire _14083 = _14082 ^ _1745;
  wire _14084 = _14081 ^ _14083;
  wire _14085 = uncoded_block[156] ^ uncoded_block[160];
  wire _14086 = _7397 ^ _14085;
  wire _14087 = _74 ^ _8589;
  wire _14088 = _14086 ^ _14087;
  wire _14089 = _14084 ^ _14088;
  wire _14090 = _14080 ^ _14089;
  wire _14091 = _6788 ^ _2521;
  wire _14092 = uncoded_block[177] ^ uncoded_block[180];
  wire _14093 = _1756 ^ _14092;
  wire _14094 = _14091 ^ _14093;
  wire _14095 = _2525 ^ _10275;
  wire _14096 = _4773 ^ _7411;
  wire _14097 = _14095 ^ _14096;
  wire _14098 = _14094 ^ _14097;
  wire _14099 = uncoded_block[201] ^ uncoded_block[204];
  wire _14100 = _6801 ^ _14099;
  wire _14101 = uncoded_block[206] ^ uncoded_block[207];
  wire _14102 = _14101 ^ _97;
  wire _14103 = _14100 ^ _14102;
  wire _14104 = _98 ^ _959;
  wire _14105 = uncoded_block[219] ^ uncoded_block[221];
  wire _14106 = _14105 ^ _4076;
  wire _14107 = _14104 ^ _14106;
  wire _14108 = _14103 ^ _14107;
  wire _14109 = _14098 ^ _14108;
  wire _14110 = _14090 ^ _14109;
  wire _14111 = _14073 ^ _14110;
  wire _14112 = _4080 ^ _2549;
  wire _14113 = uncoded_block[238] ^ uncoded_block[245];
  wire _14114 = _14113 ^ _6180;
  wire _14115 = _14112 ^ _14114;
  wire _14116 = uncoded_block[249] ^ uncoded_block[251];
  wire _14117 = uncoded_block[253] ^ uncoded_block[255];
  wire _14118 = _14116 ^ _14117;
  wire _14119 = _1786 ^ _119;
  wire _14120 = _14118 ^ _14119;
  wire _14121 = _14115 ^ _14120;
  wire _14122 = uncoded_block[265] ^ uncoded_block[269];
  wire _14123 = _14122 ^ _2566;
  wire _14124 = uncoded_block[272] ^ uncoded_block[274];
  wire _14125 = _14124 ^ _4814;
  wire _14126 = _14123 ^ _14125;
  wire _14127 = _11967 ^ _1803;
  wire _14128 = uncoded_block[289] ^ uncoded_block[294];
  wire _14129 = _14128 ^ _137;
  wire _14130 = _14127 ^ _14129;
  wire _14131 = _14126 ^ _14130;
  wire _14132 = _14121 ^ _14131;
  wire _14133 = uncoded_block[299] ^ uncoded_block[301];
  wire _14134 = _14133 ^ _4826;
  wire _14135 = uncoded_block[311] ^ uncoded_block[319];
  wire _14136 = _14135 ^ _8642;
  wire _14137 = _14134 ^ _14136;
  wire _14138 = _11984 ^ _6217;
  wire _14139 = _13084 ^ _14138;
  wire _14140 = _14137 ^ _14139;
  wire _14141 = _4841 ^ _8652;
  wire _14142 = _4132 ^ _11455;
  wire _14143 = _14141 ^ _14142;
  wire _14144 = uncoded_block[365] ^ uncoded_block[372];
  wire _14145 = _14144 ^ _4853;
  wire _14146 = _8074 ^ _14145;
  wire _14147 = _14143 ^ _14146;
  wire _14148 = _14140 ^ _14147;
  wire _14149 = _14132 ^ _14148;
  wire _14150 = uncoded_block[377] ^ uncoded_block[381];
  wire _14151 = _14150 ^ _1039;
  wire _14152 = uncoded_block[387] ^ uncoded_block[396];
  wire _14153 = _14152 ^ _2622;
  wire _14154 = _14151 ^ _14153;
  wire _14155 = _4155 ^ _3389;
  wire _14156 = _190 ^ _11473;
  wire _14157 = _14155 ^ _14156;
  wire _14158 = _14154 ^ _14157;
  wire _14159 = _5565 ^ _13112;
  wire _14160 = uncoded_block[421] ^ uncoded_block[422];
  wire _14161 = _4872 ^ _14160;
  wire _14162 = _14159 ^ _14161;
  wire _14163 = uncoded_block[427] ^ uncoded_block[429];
  wire _14164 = _8672 ^ _14163;
  wire _14165 = _7495 ^ _1066;
  wire _14166 = _14164 ^ _14165;
  wire _14167 = _14162 ^ _14166;
  wire _14168 = _14158 ^ _14167;
  wire _14169 = uncoded_block[440] ^ uncoded_block[445];
  wire _14170 = _14169 ^ _11486;
  wire _14171 = _3411 ^ _4177;
  wire _14172 = _14170 ^ _14171;
  wire _14173 = uncoded_block[453] ^ uncoded_block[457];
  wire _14174 = _14173 ^ _10926;
  wire _14175 = uncoded_block[467] ^ uncoded_block[469];
  wire _14176 = uncoded_block[474] ^ uncoded_block[477];
  wire _14177 = _14175 ^ _14176;
  wire _14178 = _14174 ^ _14177;
  wire _14179 = _14172 ^ _14178;
  wire _14180 = _7513 ^ _4895;
  wire _14181 = _8694 ^ _4898;
  wire _14182 = _14180 ^ _14181;
  wire _14183 = uncoded_block[492] ^ uncoded_block[495];
  wire _14184 = _14183 ^ _1094;
  wire _14185 = _3434 ^ _12034;
  wire _14186 = _14184 ^ _14185;
  wire _14187 = _14182 ^ _14186;
  wire _14188 = _14179 ^ _14187;
  wire _14189 = _14168 ^ _14188;
  wire _14190 = _14149 ^ _14189;
  wire _14191 = _14111 ^ _14190;
  wire _14192 = _3437 ^ _13676;
  wire _14193 = uncoded_block[515] ^ uncoded_block[519];
  wire _14194 = _14193 ^ _4210;
  wire _14195 = _14192 ^ _14194;
  wire _14196 = _7534 ^ _1114;
  wire _14197 = uncoded_block[536] ^ uncoded_block[539];
  wire _14198 = uncoded_block[540] ^ uncoded_block[541];
  wire _14199 = _14197 ^ _14198;
  wire _14200 = _14196 ^ _14199;
  wire _14201 = _14195 ^ _14200;
  wire _14202 = uncoded_block[544] ^ uncoded_block[549];
  wire _14203 = _9854 ^ _14202;
  wire _14204 = uncoded_block[555] ^ uncoded_block[558];
  wire _14205 = _14204 ^ _3461;
  wire _14206 = _14203 ^ _14205;
  wire _14207 = _7545 ^ _3467;
  wire _14208 = uncoded_block[568] ^ uncoded_block[572];
  wire _14209 = uncoded_block[573] ^ uncoded_block[577];
  wire _14210 = _14208 ^ _14209;
  wire _14211 = _14207 ^ _14210;
  wire _14212 = _14206 ^ _14211;
  wire _14213 = _14201 ^ _14212;
  wire _14214 = uncoded_block[582] ^ uncoded_block[586];
  wire _14215 = _10400 ^ _14214;
  wire _14216 = _14215 ^ _9331;
  wire _14217 = _10408 ^ _2709;
  wire _14218 = uncoded_block[605] ^ uncoded_block[606];
  wire _14219 = _14218 ^ _1942;
  wire _14220 = _14217 ^ _14219;
  wire _14221 = _14216 ^ _14220;
  wire _14222 = _2713 ^ _4242;
  wire _14223 = uncoded_block[614] ^ uncoded_block[618];
  wire _14224 = uncoded_block[622] ^ uncoded_block[624];
  wire _14225 = _14223 ^ _14224;
  wire _14226 = _14222 ^ _14225;
  wire _14227 = _8159 ^ _12071;
  wire _14228 = uncoded_block[631] ^ uncoded_block[632];
  wire _14229 = _14228 ^ _12621;
  wire _14230 = _14227 ^ _14229;
  wire _14231 = _14226 ^ _14230;
  wire _14232 = _14221 ^ _14231;
  wire _14233 = _14213 ^ _14232;
  wire _14234 = uncoded_block[649] ^ uncoded_block[650];
  wire _14235 = _2730 ^ _14234;
  wire _14236 = _6974 ^ _2738;
  wire _14237 = _14235 ^ _14236;
  wire _14238 = uncoded_block[660] ^ uncoded_block[664];
  wire _14239 = _14238 ^ _1173;
  wire _14240 = uncoded_block[667] ^ uncoded_block[673];
  wire _14241 = uncoded_block[674] ^ uncoded_block[678];
  wire _14242 = _14240 ^ _14241;
  wire _14243 = _14239 ^ _14242;
  wire _14244 = _14237 ^ _14243;
  wire _14245 = _1971 ^ _12636;
  wire _14246 = _4271 ^ _2754;
  wire _14247 = _14245 ^ _14246;
  wire _14248 = _2755 ^ _8186;
  wire _14249 = uncoded_block[698] ^ uncoded_block[701];
  wire _14250 = uncoded_block[702] ^ uncoded_block[703];
  wire _14251 = _14249 ^ _14250;
  wire _14252 = _14248 ^ _14251;
  wire _14253 = _14247 ^ _14252;
  wire _14254 = _14244 ^ _14253;
  wire _14255 = uncoded_block[704] ^ uncoded_block[706];
  wire _14256 = _14255 ^ _10448;
  wire _14257 = uncoded_block[709] ^ uncoded_block[719];
  wire _14258 = _14257 ^ _8198;
  wire _14259 = _14256 ^ _14258;
  wire _14260 = _1988 ^ _1990;
  wire _14261 = _349 ^ _7605;
  wire _14262 = _14260 ^ _14261;
  wire _14263 = _14259 ^ _14262;
  wire _14264 = uncoded_block[742] ^ uncoded_block[745];
  wire _14265 = _1996 ^ _14264;
  wire _14266 = uncoded_block[750] ^ uncoded_block[752];
  wire _14267 = _12107 ^ _14266;
  wire _14268 = _14265 ^ _14267;
  wire _14269 = _359 ^ _9914;
  wire _14270 = uncoded_block[762] ^ uncoded_block[769];
  wire _14271 = uncoded_block[770] ^ uncoded_block[772];
  wire _14272 = _14270 ^ _14271;
  wire _14273 = _14269 ^ _14272;
  wire _14274 = _14268 ^ _14273;
  wire _14275 = _14263 ^ _14274;
  wire _14276 = _14254 ^ _14275;
  wire _14277 = _14233 ^ _14276;
  wire _14278 = uncoded_block[776] ^ uncoded_block[778];
  wire _14279 = _14278 ^ _9384;
  wire _14280 = _4309 ^ _5033;
  wire _14281 = _14279 ^ _14280;
  wire _14282 = uncoded_block[794] ^ uncoded_block[796];
  wire _14283 = _14282 ^ _8223;
  wire _14284 = _385 ^ _8793;
  wire _14285 = _14283 ^ _14284;
  wire _14286 = _14281 ^ _14285;
  wire _14287 = uncoded_block[807] ^ uncoded_block[810];
  wire _14288 = _14287 ^ _2808;
  wire _14289 = _14288 ^ _2030;
  wire _14290 = uncoded_block[822] ^ uncoded_block[823];
  wire _14291 = uncoded_block[824] ^ uncoded_block[828];
  wire _14292 = _14290 ^ _14291;
  wire _14293 = _7039 ^ _4331;
  wire _14294 = _14292 ^ _14293;
  wire _14295 = _14289 ^ _14294;
  wire _14296 = _14286 ^ _14295;
  wire _14297 = _3596 ^ _5737;
  wire _14298 = _1257 ^ _4340;
  wire _14299 = _14297 ^ _14298;
  wire _14300 = uncoded_block[857] ^ uncoded_block[858];
  wire _14301 = _7049 ^ _14300;
  wire _14302 = uncoded_block[863] ^ uncoded_block[865];
  wire _14303 = _14302 ^ _5071;
  wire _14304 = _14301 ^ _14303;
  wire _14305 = _14299 ^ _14304;
  wire _14306 = _5749 ^ _416;
  wire _14307 = _6416 ^ _3608;
  wire _14308 = _14306 ^ _14307;
  wire _14309 = _4351 ^ _1272;
  wire _14310 = _2061 ^ _5085;
  wire _14311 = _14309 ^ _14310;
  wire _14312 = _14308 ^ _14311;
  wire _14313 = _14305 ^ _14312;
  wire _14314 = _14296 ^ _14313;
  wire _14315 = _428 ^ _2843;
  wire _14316 = uncoded_block[901] ^ uncoded_block[908];
  wire _14317 = uncoded_block[910] ^ uncoded_block[915];
  wire _14318 = _14316 ^ _14317;
  wire _14319 = _14315 ^ _14318;
  wire _14320 = _2852 ^ _4368;
  wire _14321 = uncoded_block[931] ^ uncoded_block[934];
  wire _14322 = _14321 ^ _2862;
  wire _14323 = _14320 ^ _14322;
  wire _14324 = _14319 ^ _14323;
  wire _14325 = _7080 ^ _453;
  wire _14326 = uncoded_block[948] ^ uncoded_block[951];
  wire _14327 = _13263 ^ _14326;
  wire _14328 = _14325 ^ _14327;
  wire _14329 = uncoded_block[952] ^ uncoded_block[955];
  wire _14330 = _14329 ^ _2090;
  wire _14331 = _14330 ^ _12729;
  wire _14332 = _14328 ^ _14331;
  wire _14333 = _14324 ^ _14332;
  wire _14334 = _8847 ^ _5112;
  wire _14335 = _11647 ^ _14334;
  wire _14336 = uncoded_block[979] ^ uncoded_block[984];
  wire _14337 = _11091 ^ _14336;
  wire _14338 = _5118 ^ _8859;
  wire _14339 = _14337 ^ _14338;
  wire _14340 = _14335 ^ _14339;
  wire _14341 = _9991 ^ _1330;
  wire _14342 = _4403 ^ _14341;
  wire _14343 = _5131 ^ _2893;
  wire _14344 = _5135 ^ _12752;
  wire _14345 = _14343 ^ _14344;
  wire _14346 = _14342 ^ _14345;
  wire _14347 = _14340 ^ _14346;
  wire _14348 = _14333 ^ _14347;
  wire _14349 = _14314 ^ _14348;
  wire _14350 = _14277 ^ _14349;
  wire _14351 = _14191 ^ _14350;
  wire _14352 = uncoded_block[1035] ^ uncoded_block[1040];
  wire _14353 = _11668 ^ _14352;
  wire _14354 = _14353 ^ _5148;
  wire _14355 = uncoded_block[1055] ^ uncoded_block[1059];
  wire _14356 = _14355 ^ _3684;
  wire _14357 = uncoded_block[1063] ^ uncoded_block[1065];
  wire _14358 = _14357 ^ _8889;
  wire _14359 = _14356 ^ _14358;
  wire _14360 = _14354 ^ _14359;
  wire _14361 = uncoded_block[1073] ^ uncoded_block[1077];
  wire _14362 = _13851 ^ _14361;
  wire _14363 = _11126 ^ _1371;
  wire _14364 = _14362 ^ _14363;
  wire _14365 = uncoded_block[1089] ^ uncoded_block[1093];
  wire _14366 = uncoded_block[1094] ^ uncoded_block[1099];
  wire _14367 = _14365 ^ _14366;
  wire _14368 = _11688 ^ _14367;
  wire _14369 = _14364 ^ _14368;
  wire _14370 = _14360 ^ _14369;
  wire _14371 = _545 ^ _2160;
  wire _14372 = uncoded_block[1105] ^ uncoded_block[1108];
  wire _14373 = _14372 ^ _2165;
  wire _14374 = _14371 ^ _14373;
  wire _14375 = _2167 ^ _3714;
  wire _14376 = uncoded_block[1122] ^ uncoded_block[1125];
  wire _14377 = _14376 ^ _6499;
  wire _14378 = _14375 ^ _14377;
  wire _14379 = _14374 ^ _14378;
  wire _14380 = uncoded_block[1135] ^ uncoded_block[1136];
  wire _14381 = _10590 ^ _14380;
  wire _14382 = _14381 ^ _10594;
  wire _14383 = _2179 ^ _10597;
  wire _14384 = _3725 ^ _8937;
  wire _14385 = _14383 ^ _14384;
  wire _14386 = _14382 ^ _14385;
  wire _14387 = _14379 ^ _14386;
  wire _14388 = _14370 ^ _14387;
  wire _14389 = uncoded_block[1157] ^ uncoded_block[1162];
  wire _14390 = _14389 ^ _13335;
  wire _14391 = _2189 ^ _11161;
  wire _14392 = _14390 ^ _14391;
  wire _14393 = uncoded_block[1176] ^ uncoded_block[1180];
  wire _14394 = _14393 ^ _2195;
  wire _14395 = _5201 ^ _3747;
  wire _14396 = _14394 ^ _14395;
  wire _14397 = _14392 ^ _14396;
  wire _14398 = uncoded_block[1194] ^ uncoded_block[1196];
  wire _14399 = _3749 ^ _14398;
  wire _14400 = _2206 ^ _2209;
  wire _14401 = _14399 ^ _14400;
  wire _14402 = _5885 ^ _5209;
  wire _14403 = _12259 ^ _2219;
  wire _14404 = _14402 ^ _14403;
  wire _14405 = _14401 ^ _14404;
  wire _14406 = _14397 ^ _14405;
  wire _14407 = uncoded_block[1218] ^ uncoded_block[1221];
  wire _14408 = _14407 ^ _7168;
  wire _14409 = _1435 ^ _12819;
  wire _14410 = _14408 ^ _14409;
  wire _14411 = _1439 ^ _2225;
  wire _14412 = uncoded_block[1234] ^ uncoded_block[1241];
  wire _14413 = _14412 ^ _1448;
  wire _14414 = _14411 ^ _14413;
  wire _14415 = _14410 ^ _14414;
  wire _14416 = uncoded_block[1248] ^ uncoded_block[1252];
  wire _14417 = _14416 ^ _8389;
  wire _14418 = uncoded_block[1262] ^ uncoded_block[1264];
  wire _14419 = _3784 ^ _14418;
  wire _14420 = _14417 ^ _14419;
  wire _14421 = _9538 ^ _7183;
  wire _14422 = _10635 ^ _14421;
  wire _14423 = _14420 ^ _14422;
  wire _14424 = _14415 ^ _14423;
  wire _14425 = _14406 ^ _14424;
  wire _14426 = _14388 ^ _14425;
  wire _14427 = _9541 ^ _3798;
  wire _14428 = _3801 ^ _645;
  wire _14429 = _14427 ^ _14428;
  wire _14430 = uncoded_block[1312] ^ uncoded_block[1313];
  wire _14431 = _8984 ^ _14430;
  wire _14432 = uncoded_block[1314] ^ uncoded_block[1315];
  wire _14433 = _14432 ^ _5926;
  wire _14434 = _14431 ^ _14433;
  wire _14435 = _14429 ^ _14434;
  wire _14436 = uncoded_block[1325] ^ uncoded_block[1331];
  wire _14437 = uncoded_block[1332] ^ uncoded_block[1335];
  wire _14438 = _14436 ^ _14437;
  wire _14439 = _4544 ^ _14438;
  wire _14440 = uncoded_block[1337] ^ uncoded_block[1342];
  wire _14441 = _14440 ^ _5268;
  wire _14442 = uncoded_block[1349] ^ uncoded_block[1351];
  wire _14443 = _14442 ^ _5272;
  wire _14444 = _14441 ^ _14443;
  wire _14445 = _14439 ^ _14444;
  wire _14446 = _14435 ^ _14445;
  wire _14447 = uncoded_block[1357] ^ uncoded_block[1360];
  wire _14448 = _14447 ^ _5275;
  wire _14449 = uncoded_block[1363] ^ uncoded_block[1369];
  wire _14450 = _14449 ^ _9573;
  wire _14451 = _14448 ^ _14450;
  wire _14452 = _7219 ^ _5288;
  wire _14453 = _12867 ^ _4568;
  wire _14454 = _14452 ^ _14453;
  wire _14455 = _14451 ^ _14454;
  wire _14456 = _3065 ^ _1517;
  wire _14457 = uncoded_block[1403] ^ uncoded_block[1405];
  wire _14458 = _14457 ^ _2300;
  wire _14459 = _14456 ^ _14458;
  wire _14460 = _8436 ^ _5962;
  wire _14461 = _705 ^ _708;
  wire _14462 = _14460 ^ _14461;
  wire _14463 = _14459 ^ _14462;
  wire _14464 = _14455 ^ _14463;
  wire _14465 = _14446 ^ _14464;
  wire _14466 = uncoded_block[1426] ^ uncoded_block[1428];
  wire _14467 = uncoded_block[1430] ^ uncoded_block[1435];
  wire _14468 = _14466 ^ _14467;
  wire _14469 = uncoded_block[1439] ^ uncoded_block[1442];
  wire _14470 = _14469 ^ _3862;
  wire _14471 = _14468 ^ _14470;
  wire _14472 = _1544 ^ _5309;
  wire _14473 = _723 ^ _2336;
  wire _14474 = _14472 ^ _14473;
  wire _14475 = _14471 ^ _14474;
  wire _14476 = _7247 ^ _9608;
  wire _14477 = _4603 ^ _3881;
  wire _14478 = _14476 ^ _14477;
  wire _14479 = uncoded_block[1480] ^ uncoded_block[1485];
  wire _14480 = _13446 ^ _14479;
  wire _14481 = _14480 ^ _13451;
  wire _14482 = _14478 ^ _14481;
  wire _14483 = _14475 ^ _14482;
  wire _14484 = uncoded_block[1496] ^ uncoded_block[1500];
  wire _14485 = _12896 ^ _14484;
  wire _14486 = _7866 ^ _7259;
  wire _14487 = _14485 ^ _14486;
  wire _14488 = uncoded_block[1515] ^ uncoded_block[1517];
  wire _14489 = _9053 ^ _14488;
  wire _14490 = _5335 ^ _14489;
  wire _14491 = _14487 ^ _14490;
  wire _14492 = uncoded_block[1531] ^ uncoded_block[1540];
  wire _14493 = _13978 ^ _14492;
  wire _14494 = _3129 ^ _13471;
  wire _14495 = _14493 ^ _14494;
  wire _14496 = uncoded_block[1550] ^ uncoded_block[1551];
  wire _14497 = _14496 ^ _7885;
  wire _14498 = uncoded_block[1562] ^ uncoded_block[1566];
  wire _14499 = _10732 ^ _14498;
  wire _14500 = _14497 ^ _14499;
  wire _14501 = _14495 ^ _14500;
  wire _14502 = _14491 ^ _14501;
  wire _14503 = _14483 ^ _14502;
  wire _14504 = _14465 ^ _14503;
  wire _14505 = _14426 ^ _14504;
  wire _14506 = uncoded_block[1573] ^ uncoded_block[1577];
  wire _14507 = uncoded_block[1578] ^ uncoded_block[1581];
  wire _14508 = _14506 ^ _14507;
  wire _14509 = _6021 ^ _14508;
  wire _14510 = _1612 ^ _3925;
  wire _14511 = uncoded_block[1588] ^ uncoded_block[1589];
  wire _14512 = uncoded_block[1591] ^ uncoded_block[1593];
  wire _14513 = _14511 ^ _14512;
  wire _14514 = _14510 ^ _14513;
  wire _14515 = _14509 ^ _14514;
  wire _14516 = _792 ^ _1620;
  wire _14517 = uncoded_block[1602] ^ uncoded_block[1605];
  wire _14518 = _11847 ^ _14517;
  wire _14519 = _14516 ^ _14518;
  wire _14520 = uncoded_block[1610] ^ uncoded_block[1614];
  wire _14521 = _6677 ^ _14520;
  wire _14522 = _14521 ^ _8508;
  wire _14523 = _14519 ^ _14522;
  wire _14524 = _14515 ^ _14523;
  wire _14525 = uncoded_block[1627] ^ uncoded_block[1628];
  wire _14526 = _14525 ^ _7305;
  wire _14527 = _7306 ^ _1642;
  wire _14528 = _14526 ^ _14527;
  wire _14529 = _2408 ^ _4673;
  wire _14530 = uncoded_block[1649] ^ uncoded_block[1651];
  wire _14531 = _12386 ^ _14530;
  wire _14532 = _14529 ^ _14531;
  wire _14533 = _14528 ^ _14532;
  wire _14534 = _9106 ^ _7925;
  wire _14535 = _823 ^ _3179;
  wire _14536 = _14534 ^ _14535;
  wire _14537 = _2422 ^ _3182;
  wire _14538 = _11319 ^ _3962;
  wire _14539 = _14537 ^ _14538;
  wire _14540 = _14536 ^ _14539;
  wire _14541 = _14533 ^ _14540;
  wire _14542 = _14524 ^ _14541;
  wire _14543 = uncoded_block[1685] ^ uncoded_block[1686];
  wire _14544 = _14543 ^ _3189;
  wire _14545 = uncoded_block[1689] ^ uncoded_block[1695];
  wire _14546 = _14545 ^ _844;
  wire _14547 = _14544 ^ _14546;
  wire _14548 = _6068 ^ _3196;
  wire _14549 = _848 ^ _3980;
  wire _14550 = _14548 ^ _14549;
  wire _14551 = _14547 ^ _14550;
  wire _14552 = uncoded_block[1715] ^ uncoded_block[1717];
  wire _14553 = _3200 ^ _14552;
  wire _14554 = _14553 ^ _14033;
  wire _14555 = _14551 ^ _14554;
  wire _14556 = _14542 ^ _14555;
  wire _14557 = _14505 ^ _14556;
  wire _14558 = _14351 ^ _14557;
  wire _14559 = _12415 ^ _3212;
  wire _14560 = uncoded_block[11] ^ uncoded_block[14];
  wire _14561 = _4 ^ _14560;
  wire _14562 = _14559 ^ _14561;
  wire _14563 = uncoded_block[17] ^ uncoded_block[22];
  wire _14564 = _5423 ^ _14563;
  wire _14565 = uncoded_block[24] ^ uncoded_block[27];
  wire _14566 = _14565 ^ _11;
  wire _14567 = _14564 ^ _14566;
  wire _14568 = _14562 ^ _14567;
  wire _14569 = uncoded_block[33] ^ uncoded_block[36];
  wire _14570 = _14569 ^ _18;
  wire _14571 = uncoded_block[39] ^ uncoded_block[41];
  wire _14572 = _14571 ^ _7965;
  wire _14573 = _14570 ^ _14572;
  wire _14574 = _23 ^ _3232;
  wire _14575 = uncoded_block[52] ^ uncoded_block[54];
  wire _14576 = _3233 ^ _14575;
  wire _14577 = _14574 ^ _14576;
  wire _14578 = _14573 ^ _14577;
  wire _14579 = _14568 ^ _14578;
  wire _14580 = _1703 ^ _7364;
  wire _14581 = _10806 ^ _9705;
  wire _14582 = _14580 ^ _14581;
  wire _14583 = uncoded_block[72] ^ uncoded_block[76];
  wire _14584 = _14583 ^ _901;
  wire _14585 = uncoded_block[79] ^ uncoded_block[82];
  wire _14586 = uncoded_block[84] ^ uncoded_block[85];
  wire _14587 = _14585 ^ _14586;
  wire _14588 = _14584 ^ _14587;
  wire _14589 = _14582 ^ _14588;
  wire _14590 = uncoded_block[86] ^ uncoded_block[90];
  wire _14591 = uncoded_block[91] ^ uncoded_block[94];
  wire _14592 = _14590 ^ _14591;
  wire _14593 = _14068 ^ _7377;
  wire _14594 = _14592 ^ _14593;
  wire _14595 = uncoded_block[105] ^ uncoded_block[107];
  wire _14596 = _14595 ^ _6123;
  wire _14597 = _6126 ^ _6769;
  wire _14598 = _14596 ^ _14597;
  wire _14599 = _14594 ^ _14598;
  wire _14600 = _14589 ^ _14599;
  wire _14601 = _14579 ^ _14600;
  wire _14602 = uncoded_block[118] ^ uncoded_block[121];
  wire _14603 = _14602 ^ _3255;
  wire _14604 = _3256 ^ _3262;
  wire _14605 = _14603 ^ _14604;
  wire _14606 = _8581 ^ _9729;
  wire _14607 = _11924 ^ _7397;
  wire _14608 = _14606 ^ _14607;
  wire _14609 = _14605 ^ _14608;
  wire _14610 = uncoded_block[156] ^ uncoded_block[163];
  wire _14611 = _14610 ^ _2516;
  wire _14612 = _11390 ^ _8591;
  wire _14613 = _14611 ^ _14612;
  wire _14614 = uncoded_block[172] ^ uncoded_block[174];
  wire _14615 = _14614 ^ _2524;
  wire _14616 = uncoded_block[187] ^ uncoded_block[190];
  wire _14617 = _5479 ^ _14616;
  wire _14618 = _14615 ^ _14617;
  wire _14619 = _14613 ^ _14618;
  wire _14620 = _14609 ^ _14619;
  wire _14621 = _6798 ^ _10277;
  wire _14622 = uncoded_block[201] ^ uncoded_block[203];
  wire _14623 = _14622 ^ _8600;
  wire _14624 = _14621 ^ _14623;
  wire _14625 = _12483 ^ _3296;
  wire _14626 = _4787 ^ _5492;
  wire _14627 = _14625 ^ _14626;
  wire _14628 = _14624 ^ _14627;
  wire _14629 = _11410 ^ _4791;
  wire _14630 = _6171 ^ _2552;
  wire _14631 = _14629 ^ _14630;
  wire _14632 = _9211 ^ _8616;
  wire _14633 = _2556 ^ _11419;
  wire _14634 = _14632 ^ _14633;
  wire _14635 = _14631 ^ _14634;
  wire _14636 = _14628 ^ _14635;
  wire _14637 = _14620 ^ _14636;
  wire _14638 = _14601 ^ _14637;
  wire _14639 = uncoded_block[257] ^ uncoded_block[258];
  wire _14640 = _14639 ^ _7438;
  wire _14641 = uncoded_block[263] ^ uncoded_block[265];
  wire _14642 = uncoded_block[269] ^ uncoded_block[270];
  wire _14643 = _14641 ^ _14642;
  wire _14644 = _14640 ^ _14643;
  wire _14645 = _6194 ^ _988;
  wire _14646 = _8625 ^ _14645;
  wire _14647 = _14644 ^ _14646;
  wire _14648 = _11428 ^ _10876;
  wire _14649 = uncoded_block[293] ^ uncoded_block[298];
  wire _14650 = _14649 ^ _1810;
  wire _14651 = _14648 ^ _14650;
  wire _14652 = uncoded_block[302] ^ uncoded_block[304];
  wire _14653 = _14652 ^ _4114;
  wire _14654 = uncoded_block[311] ^ uncoded_block[315];
  wire _14655 = _14654 ^ _13625;
  wire _14656 = _14653 ^ _14655;
  wire _14657 = _14651 ^ _14656;
  wire _14658 = _14647 ^ _14657;
  wire _14659 = _2586 ^ _1017;
  wire _14660 = _13082 ^ _14659;
  wire _14661 = _4129 ^ _4131;
  wire _14662 = uncoded_block[350] ^ uncoded_block[352];
  wire _14663 = _1023 ^ _14662;
  wire _14664 = _14661 ^ _14663;
  wire _14665 = _14660 ^ _14664;
  wire _14666 = _1028 ^ _3361;
  wire _14667 = _3362 ^ _6866;
  wire _14668 = _14666 ^ _14667;
  wire _14669 = uncoded_block[365] ^ uncoded_block[371];
  wire _14670 = _14669 ^ _1036;
  wire _14671 = uncoded_block[376] ^ uncoded_block[379];
  wire _14672 = _14671 ^ _3377;
  wire _14673 = _14670 ^ _14672;
  wire _14674 = _14668 ^ _14673;
  wire _14675 = _14665 ^ _14674;
  wire _14676 = _14658 ^ _14675;
  wire _14677 = uncoded_block[385] ^ uncoded_block[389];
  wire _14678 = uncoded_block[391] ^ uncoded_block[396];
  wire _14679 = _14677 ^ _14678;
  wire _14680 = _1051 ^ _190;
  wire _14681 = _14679 ^ _14680;
  wire _14682 = uncoded_block[413] ^ uncoded_block[416];
  wire _14683 = _8091 ^ _14682;
  wire _14684 = _4161 ^ _11477;
  wire _14685 = _14683 ^ _14684;
  wire _14686 = _14681 ^ _14685;
  wire _14687 = uncoded_block[427] ^ uncoded_block[431];
  wire _14688 = _11479 ^ _14687;
  wire _14689 = uncoded_block[432] ^ uncoded_block[435];
  wire _14690 = uncoded_block[436] ^ uncoded_block[439];
  wire _14691 = _14689 ^ _14690;
  wire _14692 = _14688 ^ _14691;
  wire _14693 = _4177 ^ _5584;
  wire _14694 = _5579 ^ _14693;
  wire _14695 = _14692 ^ _14694;
  wire _14696 = _14686 ^ _14695;
  wire _14697 = _2653 ^ _13662;
  wire _14698 = _8683 ^ _3418;
  wire _14699 = _14697 ^ _14698;
  wire _14700 = _3421 ^ _8110;
  wire _14701 = _7515 ^ _5600;
  wire _14702 = _14700 ^ _14701;
  wire _14703 = _14699 ^ _14702;
  wire _14704 = uncoded_block[500] ^ uncoded_block[504];
  wire _14705 = _2667 ^ _14704;
  wire _14706 = _9836 ^ _14705;
  wire _14707 = uncoded_block[505] ^ uncoded_block[510];
  wire _14708 = _14707 ^ _9295;
  wire _14709 = _13676 ^ _9840;
  wire _14710 = _14708 ^ _14709;
  wire _14711 = _14706 ^ _14710;
  wire _14712 = _14703 ^ _14711;
  wire _14713 = _14696 ^ _14712;
  wire _14714 = _14676 ^ _14713;
  wire _14715 = _14638 ^ _14714;
  wire _14716 = uncoded_block[527] ^ uncoded_block[529];
  wire _14717 = _13684 ^ _14716;
  wire _14718 = _8130 ^ _14717;
  wire _14719 = uncoded_block[535] ^ uncoded_block[539];
  wire _14720 = _240 ^ _14719;
  wire _14721 = uncoded_block[540] ^ uncoded_block[543];
  wire _14722 = _14721 ^ _1117;
  wire _14723 = _14720 ^ _14722;
  wire _14724 = _14718 ^ _14723;
  wire _14725 = uncoded_block[548] ^ uncoded_block[552];
  wire _14726 = _5628 ^ _14725;
  wire _14727 = _1122 ^ _6940;
  wire _14728 = _14726 ^ _14727;
  wire _14729 = _9320 ^ _7550;
  wire _14730 = _13168 ^ _11526;
  wire _14731 = _14729 ^ _14730;
  wire _14732 = _14728 ^ _14731;
  wire _14733 = _14724 ^ _14732;
  wire _14734 = _1139 ^ _3478;
  wire _14735 = _13705 ^ _4236;
  wire _14736 = _14734 ^ _14735;
  wire _14737 = uncoded_block[599] ^ uncoded_block[602];
  wire _14738 = _14737 ^ _8152;
  wire _14739 = uncoded_block[607] ^ uncoded_block[610];
  wire _14740 = _14739 ^ _7564;
  wire _14741 = _14738 ^ _14740;
  wire _14742 = _14736 ^ _14741;
  wire _14743 = uncoded_block[618] ^ uncoded_block[621];
  wire _14744 = _13713 ^ _14743;
  wire _14745 = uncoded_block[630] ^ uncoded_block[631];
  wire _14746 = _6966 ^ _14745;
  wire _14747 = _14744 ^ _14746;
  wire _14748 = _2723 ^ _4255;
  wire _14749 = _4972 ^ _296;
  wire _14750 = _14748 ^ _14749;
  wire _14751 = _14747 ^ _14750;
  wire _14752 = _14742 ^ _14751;
  wire _14753 = _14733 ^ _14752;
  wire _14754 = _8165 ^ _6974;
  wire _14755 = uncoded_block[655] ^ uncoded_block[657];
  wire _14756 = _14755 ^ _2739;
  wire _14757 = _14754 ^ _14756;
  wire _14758 = _12630 ^ _5671;
  wire _14759 = uncoded_block[671] ^ uncoded_block[676];
  wire _14760 = _311 ^ _14759;
  wire _14761 = _14758 ^ _14760;
  wire _14762 = _14757 ^ _14761;
  wire _14763 = _10440 ^ _3522;
  wire _14764 = _10442 ^ _6985;
  wire _14765 = _14763 ^ _14764;
  wire _14766 = uncoded_block[698] ^ uncoded_block[702];
  wire _14767 = _3529 ^ _14766;
  wire _14768 = _6361 ^ _6364;
  wire _14769 = _14767 ^ _14768;
  wire _14770 = _14765 ^ _14769;
  wire _14771 = _14762 ^ _14770;
  wire _14772 = _8190 ^ _10452;
  wire _14773 = _14772 ^ _10454;
  wire _14774 = uncoded_block[726] ^ uncoded_block[729];
  wire _14775 = _9904 ^ _14774;
  wire _14776 = uncoded_block[733] ^ uncoded_block[738];
  wire _14777 = _8200 ^ _14776;
  wire _14778 = _14775 ^ _14777;
  wire _14779 = _14773 ^ _14778;
  wire _14780 = _5703 ^ _9376;
  wire _14781 = _2778 ^ _9914;
  wire _14782 = _2781 ^ _2783;
  wire _14783 = _14781 ^ _14782;
  wire _14784 = _14780 ^ _14783;
  wire _14785 = _14779 ^ _14784;
  wire _14786 = _14771 ^ _14785;
  wire _14787 = _14753 ^ _14786;
  wire _14788 = uncoded_block[768] ^ uncoded_block[772];
  wire _14789 = _365 ^ _14788;
  wire _14790 = _13216 ^ _3562;
  wire _14791 = _14789 ^ _14790;
  wire _14792 = _368 ^ _12669;
  wire _14793 = uncoded_block[784] ^ uncoded_block[786];
  wire _14794 = _14793 ^ _1225;
  wire _14795 = _14792 ^ _14794;
  wire _14796 = _14791 ^ _14795;
  wire _14797 = uncoded_block[792] ^ uncoded_block[796];
  wire _14798 = _14797 ^ _8223;
  wire _14799 = _12679 ^ _5727;
  wire _14800 = _14798 ^ _14799;
  wire _14801 = _11596 ^ _5045;
  wire _14802 = uncoded_block[821] ^ uncoded_block[825];
  wire _14803 = _4325 ^ _14802;
  wire _14804 = _14801 ^ _14803;
  wire _14805 = _14800 ^ _14804;
  wire _14806 = _14796 ^ _14805;
  wire _14807 = uncoded_block[831] ^ uncoded_block[834];
  wire _14808 = _6401 ^ _14807;
  wire _14809 = uncoded_block[837] ^ uncoded_block[840];
  wire _14810 = _14809 ^ _2036;
  wire _14811 = _14808 ^ _14810;
  wire _14812 = uncoded_block[843] ^ uncoded_block[846];
  wire _14813 = _14812 ^ _3599;
  wire _14814 = uncoded_block[850] ^ uncoded_block[851];
  wire _14815 = _14814 ^ _11048;
  wire _14816 = _14813 ^ _14815;
  wire _14817 = _14811 ^ _14816;
  wire _14818 = _8812 ^ _5066;
  wire _14819 = _4344 ^ _5749;
  wire _14820 = _14818 ^ _14819;
  wire _14821 = uncoded_block[884] ^ uncoded_block[886];
  wire _14822 = _2836 ^ _14821;
  wire _14823 = _7061 ^ _14822;
  wire _14824 = _14820 ^ _14823;
  wire _14825 = _14817 ^ _14824;
  wire _14826 = _14806 ^ _14825;
  wire _14827 = uncoded_block[891] ^ uncoded_block[892];
  wire _14828 = _9416 ^ _14827;
  wire _14829 = uncoded_block[895] ^ uncoded_block[898];
  wire _14830 = _14829 ^ _2844;
  wire _14831 = _14828 ^ _14830;
  wire _14832 = _2065 ^ _9421;
  wire _14833 = _12165 ^ _3629;
  wire _14834 = _14832 ^ _14833;
  wire _14835 = _14831 ^ _14834;
  wire _14836 = _2073 ^ _2855;
  wire _14837 = _4371 ^ _2858;
  wire _14838 = _14836 ^ _14837;
  wire _14839 = _1299 ^ _8269;
  wire _14840 = _5104 ^ _10529;
  wire _14841 = _14839 ^ _14840;
  wire _14842 = _14838 ^ _14841;
  wire _14843 = _14835 ^ _14842;
  wire _14844 = uncoded_block[963] ^ uncoded_block[965];
  wire _14845 = _14844 ^ _467;
  wire _14846 = _14845 ^ _11089;
  wire _14847 = _11091 ^ _5790;
  wire _14848 = _14847 ^ _3660;
  wire _14849 = _14846 ^ _14848;
  wire _14850 = uncoded_block[988] ^ uncoded_block[991];
  wire _14851 = uncoded_block[995] ^ uncoded_block[1005];
  wire _14852 = _14850 ^ _14851;
  wire _14853 = _4410 ^ _4412;
  wire _14854 = _14852 ^ _14853;
  wire _14855 = uncoded_block[1020] ^ uncoded_block[1023];
  wire _14856 = _8871 ^ _14855;
  wire _14857 = uncoded_block[1032] ^ uncoded_block[1038];
  wire _14858 = _2121 ^ _14857;
  wire _14859 = _14856 ^ _14858;
  wire _14860 = _14854 ^ _14859;
  wire _14861 = _14849 ^ _14860;
  wire _14862 = _14843 ^ _14861;
  wire _14863 = _14826 ^ _14862;
  wire _14864 = _14787 ^ _14863;
  wire _14865 = _14715 ^ _14864;
  wire _14866 = _2130 ^ _8309;
  wire _14867 = uncoded_block[1049] ^ uncoded_block[1053];
  wire _14868 = _14867 ^ _4430;
  wire _14869 = _14866 ^ _14868;
  wire _14870 = _1363 ^ _3685;
  wire _14871 = _12213 ^ _5158;
  wire _14872 = _14870 ^ _14871;
  wire _14873 = _14869 ^ _14872;
  wire _14874 = _2924 ^ _11126;
  wire _14875 = _10575 ^ _2928;
  wire _14876 = _14874 ^ _14875;
  wire _14877 = _1374 ^ _5840;
  wire _14878 = _5166 ^ _4444;
  wire _14879 = _14877 ^ _14878;
  wire _14880 = _14876 ^ _14879;
  wire _14881 = _14873 ^ _14880;
  wire _14882 = uncoded_block[1111] ^ uncoded_block[1113];
  wire _14883 = uncoded_block[1114] ^ uncoded_block[1124];
  wire _14884 = _14882 ^ _14883;
  wire _14885 = _10028 ^ _14884;
  wire _14886 = _5854 ^ _6499;
  wire _14887 = uncoded_block[1131] ^ uncoded_block[1134];
  wire _14888 = _14887 ^ _2950;
  wire _14889 = _14886 ^ _14888;
  wire _14890 = _14885 ^ _14889;
  wire _14891 = _5859 ^ _2179;
  wire _14892 = _5862 ^ _2956;
  wire _14893 = _14891 ^ _14892;
  wire _14894 = uncoded_block[1154] ^ uncoded_block[1159];
  wire _14895 = _8351 ^ _14894;
  wire _14896 = _6511 ^ _5193;
  wire _14897 = _14895 ^ _14896;
  wire _14898 = _14893 ^ _14897;
  wire _14899 = _14890 ^ _14898;
  wire _14900 = _14881 ^ _14899;
  wire _14901 = uncoded_block[1173] ^ uncoded_block[1175];
  wire _14902 = _5870 ^ _14901;
  wire _14903 = _3740 ^ _3742;
  wire _14904 = _14902 ^ _14903;
  wire _14905 = _1417 ^ _4486;
  wire _14906 = _9508 ^ _596;
  wire _14907 = _14905 ^ _14906;
  wire _14908 = _14904 ^ _14907;
  wire _14909 = _8951 ^ _2206;
  wire _14910 = _2978 ^ _2216;
  wire _14911 = _14909 ^ _14910;
  wire _14912 = uncoded_block[1209] ^ uncoded_block[1212];
  wire _14913 = _14912 ^ _2982;
  wire _14914 = uncoded_block[1216] ^ uncoded_block[1219];
  wire _14915 = _14914 ^ _1433;
  wire _14916 = _14913 ^ _14915;
  wire _14917 = _14911 ^ _14916;
  wire _14918 = _14908 ^ _14917;
  wire _14919 = uncoded_block[1230] ^ uncoded_block[1232];
  wire _14920 = _1435 ^ _14919;
  wire _14921 = uncoded_block[1233] ^ uncoded_block[1235];
  wire _14922 = _14921 ^ _1443;
  wire _14923 = _14920 ^ _14922;
  wire _14924 = _9527 ^ _6544;
  wire _14925 = _14923 ^ _14924;
  wire _14926 = uncoded_block[1256] ^ uncoded_block[1265];
  wire _14927 = _6545 ^ _14926;
  wire _14928 = uncoded_block[1269] ^ uncoded_block[1275];
  wire _14929 = _3008 ^ _14928;
  wire _14930 = _14927 ^ _14929;
  wire _14931 = uncoded_block[1282] ^ uncoded_block[1290];
  wire _14932 = _5908 ^ _14931;
  wire _14933 = _10646 ^ _4531;
  wire _14934 = _14932 ^ _14933;
  wire _14935 = _14930 ^ _14934;
  wire _14936 = _14925 ^ _14935;
  wire _14937 = _14918 ^ _14936;
  wire _14938 = _14900 ^ _14937;
  wire _14939 = uncoded_block[1299] ^ uncoded_block[1302];
  wire _14940 = _14939 ^ _2255;
  wire _14941 = _8991 ^ _8407;
  wire _14942 = _14940 ^ _14941;
  wire _14943 = _1483 ^ _2262;
  wire _14944 = _12287 ^ _3029;
  wire _14945 = _14943 ^ _14944;
  wire _14946 = _14942 ^ _14945;
  wire _14947 = _8998 ^ _8413;
  wire _14948 = _13396 ^ _14947;
  wire _14949 = _5259 ^ _2277;
  wire _14950 = uncoded_block[1342] ^ uncoded_block[1344];
  wire _14951 = _14950 ^ _3039;
  wire _14952 = _14949 ^ _14951;
  wire _14953 = _14948 ^ _14952;
  wire _14954 = _14946 ^ _14953;
  wire _14955 = _669 ^ _5938;
  wire _14956 = uncoded_block[1355] ^ uncoded_block[1358];
  wire _14957 = _14956 ^ _6588;
  wire _14958 = _14955 ^ _14957;
  wire _14959 = uncoded_block[1367] ^ uncoded_block[1372];
  wire _14960 = uncoded_block[1373] ^ uncoded_block[1375];
  wire _14961 = _14959 ^ _14960;
  wire _14962 = _11225 ^ _14961;
  wire _14963 = _14958 ^ _14962;
  wire _14964 = _7217 ^ _7219;
  wire _14965 = _3059 ^ _13412;
  wire _14966 = _14964 ^ _14965;
  wire _14967 = _13416 ^ _6600;
  wire _14968 = uncoded_block[1404] ^ uncoded_block[1406];
  wire _14969 = _9016 ^ _14968;
  wire _14970 = _14967 ^ _14969;
  wire _14971 = _14966 ^ _14970;
  wire _14972 = _14963 ^ _14971;
  wire _14973 = _14954 ^ _14972;
  wire _14974 = _4580 ^ _6607;
  wire _14975 = _3853 ^ _709;
  wire _14976 = _14974 ^ _14975;
  wire _14977 = uncoded_block[1427] ^ uncoded_block[1431];
  wire _14978 = uncoded_block[1435] ^ uncoded_block[1437];
  wire _14979 = _14977 ^ _14978;
  wire _14980 = _13432 ^ _6613;
  wire _14981 = _14979 ^ _14980;
  wire _14982 = _14976 ^ _14981;
  wire _14983 = uncoded_block[1448] ^ uncoded_block[1452];
  wire _14984 = _3084 ^ _14983;
  wire _14985 = uncoded_block[1457] ^ uncoded_block[1462];
  wire _14986 = _2328 ^ _14985;
  wire _14987 = _14984 ^ _14986;
  wire _14988 = _9602 ^ _7247;
  wire _14989 = uncoded_block[1473] ^ uncoded_block[1475];
  wire _14990 = _1551 ^ _14989;
  wire _14991 = _14988 ^ _14990;
  wire _14992 = _14987 ^ _14991;
  wire _14993 = _14982 ^ _14992;
  wire _14994 = _3884 ^ _12342;
  wire _14995 = uncoded_block[1487] ^ uncoded_block[1490];
  wire _14996 = _7861 ^ _14995;
  wire _14997 = _14994 ^ _14996;
  wire _14998 = _3890 ^ _6634;
  wire _14999 = _1571 ^ _3893;
  wire _15000 = _14998 ^ _14999;
  wire _15001 = _14997 ^ _15000;
  wire _15002 = uncoded_block[1509] ^ uncoded_block[1510];
  wire _15003 = _7262 ^ _15002;
  wire _15004 = uncoded_block[1519] ^ uncoded_block[1520];
  wire _15005 = _15004 ^ _3900;
  wire _15006 = _15003 ^ _15005;
  wire _15007 = uncoded_block[1528] ^ uncoded_block[1531];
  wire _15008 = _9626 ^ _15007;
  wire _15009 = uncoded_block[1536] ^ uncoded_block[1538];
  wire _15010 = _12914 ^ _15009;
  wire _15011 = _15008 ^ _15010;
  wire _15012 = _15006 ^ _15011;
  wire _15013 = _15001 ^ _15012;
  wire _15014 = _14993 ^ _15013;
  wire _15015 = _14973 ^ _15014;
  wire _15016 = _14938 ^ _15015;
  wire _15017 = _3128 ^ _1590;
  wire _15018 = _2367 ^ _6013;
  wire _15019 = _15017 ^ _15018;
  wire _15020 = uncoded_block[1551] ^ uncoded_block[1553];
  wire _15021 = _15020 ^ _1596;
  wire _15022 = uncoded_block[1559] ^ uncoded_block[1562];
  wire _15023 = _15022 ^ _776;
  wire _15024 = _15021 ^ _15023;
  wire _15025 = _15019 ^ _15024;
  wire _15026 = uncoded_block[1571] ^ uncoded_block[1572];
  wire _15027 = _1606 ^ _15026;
  wire _15028 = _4647 ^ _3920;
  wire _15029 = _15027 ^ _15028;
  wire _15030 = _2383 ^ _6031;
  wire _15031 = uncoded_block[1586] ^ uncoded_block[1588];
  wire _15032 = _15031 ^ _12934;
  wire _15033 = _15030 ^ _15032;
  wire _15034 = _15029 ^ _15033;
  wire _15035 = _15025 ^ _15034;
  wire _15036 = _791 ^ _1620;
  wire _15037 = _1621 ^ _3936;
  wire _15038 = _15036 ^ _15037;
  wire _15039 = _3153 ^ _7908;
  wire _15040 = uncoded_block[1614] ^ uncoded_block[1620];
  wire _15041 = _15040 ^ _7912;
  wire _15042 = _15039 ^ _15041;
  wire _15043 = _15038 ^ _15042;
  wire _15044 = _10185 ^ _4667;
  wire _15045 = _4668 ^ _7308;
  wire _15046 = _15044 ^ _15045;
  wire _15047 = _1646 ^ _1649;
  wire _15048 = uncoded_block[1658] ^ uncoded_block[1661];
  wire _15049 = _13506 ^ _15048;
  wire _15050 = _15047 ^ _15049;
  wire _15051 = _15046 ^ _15050;
  wire _15052 = _15043 ^ _15051;
  wire _15053 = _15035 ^ _15052;
  wire _15054 = _6058 ^ _8521;
  wire _15055 = uncoded_block[1673] ^ uncoded_block[1677];
  wire _15056 = _15055 ^ _6061;
  wire _15057 = _15054 ^ _15056;
  wire _15058 = uncoded_block[1691] ^ uncoded_block[1696];
  wire _15059 = _3967 ^ _15058;
  wire _15060 = _14544 ^ _15059;
  wire _15061 = _15057 ^ _15060;
  wire _15062 = _5409 ^ _3975;
  wire _15063 = uncoded_block[1705] ^ uncoded_block[1706];
  wire _15064 = _15063 ^ _848;
  wire _15065 = _15062 ^ _15064;
  wire _15066 = _11879 ^ _2443;
  wire _15067 = _15066 ^ uncoded_block[1722];
  wire _15068 = _15065 ^ _15067;
  wire _15069 = _15061 ^ _15068;
  wire _15070 = _15053 ^ _15069;
  wire _15071 = _15016 ^ _15070;
  wire _15072 = _14865 ^ _15071;
  wire _15073 = uncoded_block[6] ^ uncoded_block[10];
  wire _15074 = _3210 ^ _15073;
  wire _15075 = uncoded_block[12] ^ uncoded_block[14];
  wire _15076 = uncoded_block[19] ^ uncoded_block[22];
  wire _15077 = _15075 ^ _15076;
  wire _15078 = _15074 ^ _15077;
  wire _15079 = _11343 ^ _1693;
  wire _15080 = uncoded_block[32] ^ uncoded_block[34];
  wire _15081 = _15080 ^ _2466;
  wire _15082 = _15079 ^ _15081;
  wire _15083 = _15078 ^ _15082;
  wire _15084 = _3230 ^ _6736;
  wire _15085 = _8554 ^ _4726;
  wire _15086 = _15084 ^ _15085;
  wire _15087 = uncoded_block[57] ^ uncoded_block[58];
  wire _15088 = _10238 ^ _15087;
  wire _15089 = _11355 ^ _1706;
  wire _15090 = _15088 ^ _15089;
  wire _15091 = _15086 ^ _15090;
  wire _15092 = _15083 ^ _15091;
  wire _15093 = _1711 ^ _39;
  wire _15094 = _11363 ^ _2483;
  wire _15095 = _15093 ^ _15094;
  wire _15096 = _9713 ^ _903;
  wire _15097 = uncoded_block[100] ^ uncoded_block[101];
  wire _15098 = _9715 ^ _15097;
  wire _15099 = _15096 ^ _15098;
  wire _15100 = _15095 ^ _15099;
  wire _15101 = uncoded_block[102] ^ uncoded_block[103];
  wire _15102 = _15101 ^ _2490;
  wire _15103 = uncoded_block[109] ^ uncoded_block[112];
  wire _15104 = _1722 ^ _15103;
  wire _15105 = _15102 ^ _15104;
  wire _15106 = _54 ^ _13016;
  wire _15107 = _917 ^ _1735;
  wire _15108 = _15106 ^ _15107;
  wire _15109 = _15105 ^ _15108;
  wire _15110 = _15100 ^ _15109;
  wire _15111 = _15092 ^ _15110;
  wire _15112 = uncoded_block[133] ^ uncoded_block[135];
  wire _15113 = _15112 ^ _9729;
  wire _15114 = uncoded_block[142] ^ uncoded_block[143];
  wire _15115 = _15114 ^ _5463;
  wire _15116 = _15113 ^ _15115;
  wire _15117 = _3268 ^ _8003;
  wire _15118 = uncoded_block[159] ^ uncoded_block[160];
  wire _15119 = _5470 ^ _15118;
  wire _15120 = _15117 ^ _15119;
  wire _15121 = _15116 ^ _15120;
  wire _15122 = _4053 ^ _6787;
  wire _15123 = uncoded_block[171] ^ uncoded_block[173];
  wire _15124 = _7399 ^ _15123;
  wire _15125 = _15122 ^ _15124;
  wire _15126 = uncoded_block[175] ^ uncoded_block[177];
  wire _15127 = _15126 ^ _7403;
  wire _15128 = _13583 ^ _2528;
  wire _15129 = _15127 ^ _15128;
  wire _15130 = _15125 ^ _15129;
  wire _15131 = _15121 ^ _15130;
  wire _15132 = _4062 ^ _7409;
  wire _15133 = _4776 ^ _3284;
  wire _15134 = _15132 ^ _15133;
  wire _15135 = uncoded_block[197] ^ uncoded_block[200];
  wire _15136 = _15135 ^ _4070;
  wire _15137 = _8600 ^ _3292;
  wire _15138 = _15136 ^ _15137;
  wire _15139 = _15134 ^ _15138;
  wire _15140 = _1767 ^ _8606;
  wire _15141 = _3298 ^ _2545;
  wire _15142 = _15140 ^ _15141;
  wire _15143 = _6168 ^ _4081;
  wire _15144 = uncoded_block[240] ^ uncoded_block[243];
  wire _15145 = _2552 ^ _15144;
  wire _15146 = _15143 ^ _15145;
  wire _15147 = _15142 ^ _15146;
  wire _15148 = _15139 ^ _15147;
  wire _15149 = _15131 ^ _15148;
  wire _15150 = _15111 ^ _15149;
  wire _15151 = _6180 ^ _13053;
  wire _15152 = _14117 ^ _13055;
  wire _15153 = _15151 ^ _15152;
  wire _15154 = uncoded_block[265] ^ uncoded_block[268];
  wire _15155 = _15154 ^ _1793;
  wire _15156 = _15155 ^ _5514;
  wire _15157 = _15153 ^ _15156;
  wire _15158 = _11967 ^ _8632;
  wire _15159 = uncoded_block[287] ^ uncoded_block[290];
  wire _15160 = _15159 ^ _2573;
  wire _15161 = _15158 ^ _15160;
  wire _15162 = _10312 ^ _8636;
  wire _15163 = uncoded_block[303] ^ uncoded_block[309];
  wire _15164 = _15163 ^ _3338;
  wire _15165 = _15162 ^ _15164;
  wire _15166 = _15161 ^ _15165;
  wire _15167 = _15157 ^ _15166;
  wire _15168 = uncoded_block[314] ^ uncoded_block[317];
  wire _15169 = _15168 ^ _1008;
  wire _15170 = _3346 ^ _11444;
  wire _15171 = _15169 ^ _15170;
  wire _15172 = uncoded_block[330] ^ uncoded_block[333];
  wire _15173 = uncoded_block[334] ^ uncoded_block[338];
  wire _15174 = _15172 ^ _15173;
  wire _15175 = _4840 ^ _6859;
  wire _15176 = _15174 ^ _15175;
  wire _15177 = _15171 ^ _15176;
  wire _15178 = uncoded_block[347] ^ uncoded_block[350];
  wire _15179 = uncoded_block[351] ^ uncoded_block[353];
  wire _15180 = _15178 ^ _15179;
  wire _15181 = _6221 ^ _1031;
  wire _15182 = _15180 ^ _15181;
  wire _15183 = uncoded_block[366] ^ uncoded_block[368];
  wire _15184 = _15183 ^ _169;
  wire _15185 = _15184 ^ _13641;
  wire _15186 = _15182 ^ _15185;
  wire _15187 = _15177 ^ _15186;
  wire _15188 = _15167 ^ _15187;
  wire _15189 = _1039 ^ _1045;
  wire _15190 = _3383 ^ _6881;
  wire _15191 = _15189 ^ _15190;
  wire _15192 = uncoded_block[401] ^ uncoded_block[406];
  wire _15193 = _2622 ^ _15192;
  wire _15194 = _190 ^ _5564;
  wire _15195 = _15193 ^ _15194;
  wire _15196 = _15191 ^ _15195;
  wire _15197 = uncoded_block[418] ^ uncoded_block[420];
  wire _15198 = _3396 ^ _15197;
  wire _15199 = _1062 ^ _6894;
  wire _15200 = _15198 ^ _15199;
  wire _15201 = uncoded_block[430] ^ uncoded_block[434];
  wire _15202 = _15201 ^ _7497;
  wire _15203 = _205 ^ _3409;
  wire _15204 = _15202 ^ _15203;
  wire _15205 = _15200 ^ _15204;
  wire _15206 = _15196 ^ _15205;
  wire _15207 = uncoded_block[458] ^ uncoded_block[464];
  wire _15208 = _212 ^ _15207;
  wire _15209 = _14171 ^ _15208;
  wire _15210 = _1874 ^ _3418;
  wire _15211 = uncoded_block[478] ^ uncoded_block[482];
  wire _15212 = uncoded_block[483] ^ uncoded_block[484];
  wire _15213 = _15211 ^ _15212;
  wire _15214 = _15210 ^ _15213;
  wire _15215 = _15209 ^ _15214;
  wire _15216 = _224 ^ _9832;
  wire _15217 = _4902 ^ _1097;
  wire _15218 = _15216 ^ _15217;
  wire _15219 = _2671 ^ _231;
  wire _15220 = uncoded_block[512] ^ uncoded_block[514];
  wire _15221 = _15220 ^ _9840;
  wire _15222 = _15219 ^ _15221;
  wire _15223 = _15218 ^ _15222;
  wire _15224 = _15215 ^ _15223;
  wire _15225 = _15206 ^ _15224;
  wire _15226 = _15188 ^ _15225;
  wire _15227 = _15150 ^ _15226;
  wire _15228 = _6289 ^ _1900;
  wire _15229 = _8130 ^ _15228;
  wire _15230 = uncoded_block[530] ^ uncoded_block[534];
  wire _15231 = _15230 ^ _6932;
  wire _15232 = _5619 ^ _9854;
  wire _15233 = _15231 ^ _15232;
  wire _15234 = _15229 ^ _15233;
  wire _15235 = _1909 ^ _1912;
  wire _15236 = uncoded_block[552] ^ uncoded_block[554];
  wire _15237 = _15236 ^ _12051;
  wire _15238 = _15235 ^ _15237;
  wire _15239 = uncoded_block[564] ^ uncoded_block[570];
  wire _15240 = _15239 ^ _262;
  wire _15241 = _13695 ^ _15240;
  wire _15242 = _15238 ^ _15241;
  wire _15243 = _15234 ^ _15242;
  wire _15244 = _6947 ^ _1933;
  wire _15245 = _1932 ^ _15244;
  wire _15246 = _270 ^ _4950;
  wire _15247 = uncoded_block[594] ^ uncoded_block[595];
  wire _15248 = _9330 ^ _15247;
  wire _15249 = _15246 ^ _15248;
  wire _15250 = _15245 ^ _15249;
  wire _15251 = _8149 ^ _3486;
  wire _15252 = uncoded_block[600] ^ uncoded_block[603];
  wire _15253 = _15252 ^ _8152;
  wire _15254 = _15251 ^ _15253;
  wire _15255 = _1942 ^ _6957;
  wire _15256 = _15255 ^ _5654;
  wire _15257 = _15254 ^ _15256;
  wire _15258 = _15250 ^ _15257;
  wire _15259 = _15243 ^ _15258;
  wire _15260 = _4243 ^ _3495;
  wire _15261 = uncoded_block[624] ^ uncoded_block[627];
  wire _15262 = uncoded_block[629] ^ uncoded_block[634];
  wire _15263 = _15261 ^ _15262;
  wire _15264 = _15260 ^ _15263;
  wire _15265 = _4249 ^ _12624;
  wire _15266 = _6338 ^ _14234;
  wire _15267 = _15265 ^ _15266;
  wire _15268 = _15264 ^ _15267;
  wire _15269 = _4975 ^ _3508;
  wire _15270 = uncoded_block[661] ^ uncoded_block[663];
  wire _15271 = _3513 ^ _15270;
  wire _15272 = _15269 ^ _15271;
  wire _15273 = uncoded_block[664] ^ uncoded_block[666];
  wire _15274 = _15273 ^ _10990;
  wire _15275 = uncoded_block[669] ^ uncoded_block[673];
  wire _15276 = _15275 ^ _2748;
  wire _15277 = _15274 ^ _15276;
  wire _15278 = _15272 ^ _15277;
  wire _15279 = _15268 ^ _15278;
  wire _15280 = uncoded_block[679] ^ uncoded_block[682];
  wire _15281 = uncoded_block[685] ^ uncoded_block[686];
  wire _15282 = _15280 ^ _15281;
  wire _15283 = _2754 ^ _4272;
  wire _15284 = _15282 ^ _15283;
  wire _15285 = _328 ^ _6360;
  wire _15286 = _333 ^ _14250;
  wire _15287 = _15285 ^ _15286;
  wire _15288 = _15284 ^ _15287;
  wire _15289 = uncoded_block[713] ^ uncoded_block[718];
  wire _15290 = _15289 ^ _341;
  wire _15291 = _1193 ^ _15290;
  wire _15292 = uncoded_block[722] ^ uncoded_block[726];
  wire _15293 = _15292 ^ _4286;
  wire _15294 = _5005 ^ _1995;
  wire _15295 = _15293 ^ _15294;
  wire _15296 = _15291 ^ _15295;
  wire _15297 = _15288 ^ _15296;
  wire _15298 = _15279 ^ _15297;
  wire _15299 = _15259 ^ _15298;
  wire _15300 = uncoded_block[738] ^ uncoded_block[742];
  wire _15301 = uncoded_block[743] ^ uncoded_block[748];
  wire _15302 = _15300 ^ _15301;
  wire _15303 = _14266 ^ _12663;
  wire _15304 = _15302 ^ _15303;
  wire _15305 = uncoded_block[756] ^ uncoded_block[757];
  wire _15306 = _15305 ^ _5019;
  wire _15307 = _364 ^ _1218;
  wire _15308 = _15306 ^ _15307;
  wire _15309 = _15304 ^ _15308;
  wire _15310 = uncoded_block[771] ^ uncoded_block[775];
  wire _15311 = _15310 ^ _2014;
  wire _15312 = _15311 ^ _2020;
  wire _15313 = _382 ^ _2022;
  wire _15314 = _386 ^ _8793;
  wire _15315 = _15313 ^ _15314;
  wire _15316 = _15312 ^ _15315;
  wire _15317 = _15309 ^ _15316;
  wire _15318 = uncoded_block[811] ^ uncoded_block[813];
  wire _15319 = _392 ^ _15318;
  wire _15320 = uncoded_block[820] ^ uncoded_block[823];
  wire _15321 = _11597 ^ _15320;
  wire _15322 = _15319 ^ _15321;
  wire _15323 = _1246 ^ _8800;
  wire _15324 = uncoded_block[832] ^ uncoded_block[834];
  wire _15325 = _15324 ^ _1253;
  wire _15326 = _15323 ^ _15325;
  wire _15327 = _15322 ^ _15326;
  wire _15328 = _2815 ^ _3597;
  wire _15329 = uncoded_block[846] ^ uncoded_block[853];
  wire _15330 = uncoded_block[855] ^ uncoded_block[857];
  wire _15331 = _15329 ^ _15330;
  wire _15332 = _15328 ^ _15331;
  wire _15333 = _2827 ^ _12150;
  wire _15334 = _11615 ^ _15333;
  wire _15335 = _15332 ^ _15334;
  wire _15336 = _15327 ^ _15335;
  wire _15337 = _15317 ^ _15336;
  wire _15338 = _2831 ^ _420;
  wire _15339 = uncoded_block[884] ^ uncoded_block[888];
  wire _15340 = _7062 ^ _15339;
  wire _15341 = _15338 ^ _15340;
  wire _15342 = uncoded_block[889] ^ uncoded_block[891];
  wire _15343 = uncoded_block[893] ^ uncoded_block[897];
  wire _15344 = _15342 ^ _15343;
  wire _15345 = uncoded_block[904] ^ uncoded_block[906];
  wire _15346 = _10508 ^ _15345;
  wire _15347 = _15344 ^ _15346;
  wire _15348 = _15341 ^ _15347;
  wire _15349 = _6428 ^ _12708;
  wire _15350 = uncoded_block[918] ^ uncoded_block[919];
  wire _15351 = _2852 ^ _15350;
  wire _15352 = _15349 ^ _15351;
  wire _15353 = _3632 ^ _1295;
  wire _15354 = uncoded_block[928] ^ uncoded_block[934];
  wire _15355 = uncoded_block[936] ^ uncoded_block[941];
  wire _15356 = _15354 ^ _15355;
  wire _15357 = _15353 ^ _15356;
  wire _15358 = _15352 ^ _15357;
  wire _15359 = _15348 ^ _15358;
  wire _15360 = _2086 ^ _8274;
  wire _15361 = _461 ^ _1307;
  wire _15362 = _15360 ^ _15361;
  wire _15363 = uncoded_block[966] ^ uncoded_block[970];
  wire _15364 = _12179 ^ _15363;
  wire _15365 = _468 ^ _5789;
  wire _15366 = _15364 ^ _15365;
  wire _15367 = _15362 ^ _15366;
  wire _15368 = _2100 ^ _8287;
  wire _15369 = uncoded_block[987] ^ uncoded_block[989];
  wire _15370 = _15369 ^ _4401;
  wire _15371 = _15368 ^ _15370;
  wire _15372 = uncoded_block[994] ^ uncoded_block[999];
  wire _15373 = uncoded_block[1000] ^ uncoded_block[1005];
  wire _15374 = _15372 ^ _15373;
  wire _15375 = _1327 ^ _4410;
  wire _15376 = _15374 ^ _15375;
  wire _15377 = _15371 ^ _15376;
  wire _15378 = _15367 ^ _15377;
  wire _15379 = _15359 ^ _15378;
  wire _15380 = _15337 ^ _15379;
  wire _15381 = _15299 ^ _15380;
  wire _15382 = _15227 ^ _15381;
  wire _15383 = _2117 ^ _5134;
  wire _15384 = _8871 ^ _8301;
  wire _15385 = _15383 ^ _15384;
  wire _15386 = _1339 ^ _4418;
  wire _15387 = uncoded_block[1039] ^ uncoded_block[1042];
  wire _15388 = _6474 ^ _15387;
  wire _15389 = _15386 ^ _15388;
  wire _15390 = _15385 ^ _15389;
  wire _15391 = _2133 ^ _5147;
  wire _15392 = uncoded_block[1058] ^ uncoded_block[1062];
  wire _15393 = _8311 ^ _15392;
  wire _15394 = _15391 ^ _15393;
  wire _15395 = uncoded_block[1064] ^ uncoded_block[1067];
  wire _15396 = uncoded_block[1070] ^ uncoded_block[1073];
  wire _15397 = _15395 ^ _15396;
  wire _15398 = _15397 ^ _12773;
  wire _15399 = _15394 ^ _15398;
  wire _15400 = _15390 ^ _15399;
  wire _15401 = uncoded_block[1084] ^ uncoded_block[1087];
  wire _15402 = _15401 ^ _8906;
  wire _15403 = _11137 ^ _10026;
  wire _15404 = _15402 ^ _15403;
  wire _15405 = uncoded_block[1101] ^ uncoded_block[1104];
  wire _15406 = _5846 ^ _15405;
  wire _15407 = uncoded_block[1111] ^ uncoded_block[1114];
  wire _15408 = _14372 ^ _15407;
  wire _15409 = _15406 ^ _15408;
  wire _15410 = _15404 ^ _15409;
  wire _15411 = _13322 ^ _8920;
  wire _15412 = _4455 ^ _12789;
  wire _15413 = _15411 ^ _15412;
  wire _15414 = _1393 ^ _10591;
  wire _15415 = _6500 ^ _15414;
  wire _15416 = _15413 ^ _15415;
  wire _15417 = _15410 ^ _15416;
  wire _15418 = _15400 ^ _15417;
  wire _15419 = _8929 ^ _3721;
  wire _15420 = uncoded_block[1148] ^ uncoded_block[1152];
  wire _15421 = _10597 ^ _15420;
  wire _15422 = _15419 ^ _15421;
  wire _15423 = _6507 ^ _9502;
  wire _15424 = _5193 ^ _1408;
  wire _15425 = _15423 ^ _15424;
  wire _15426 = _15422 ^ _15425;
  wire _15427 = _8362 ^ _5200;
  wire _15428 = uncoded_block[1187] ^ uncoded_block[1192];
  wire _15429 = _3746 ^ _15428;
  wire _15430 = _15427 ^ _15429;
  wire _15431 = uncoded_block[1198] ^ uncoded_block[1202];
  wire _15432 = _1421 ^ _15431;
  wire _15433 = _2209 ^ _6530;
  wire _15434 = _15432 ^ _15433;
  wire _15435 = _15430 ^ _15434;
  wire _15436 = _15426 ^ _15435;
  wire _15437 = _11726 ^ _606;
  wire _15438 = _612 ^ _5894;
  wire _15439 = _15437 ^ _15438;
  wire _15440 = _1440 ^ _11181;
  wire _15441 = uncoded_block[1239] ^ uncoded_block[1240];
  wire _15442 = _15441 ^ _10627;
  wire _15443 = _15440 ^ _15442;
  wire _15444 = _15439 ^ _15443;
  wire _15445 = _11734 ^ _1449;
  wire _15446 = _1451 ^ _7778;
  wire _15447 = _15445 ^ _15446;
  wire _15448 = _3786 ^ _1459;
  wire _15449 = _13370 ^ _15448;
  wire _15450 = _15447 ^ _15449;
  wire _15451 = _15444 ^ _15450;
  wire _15452 = _15436 ^ _15451;
  wire _15453 = _15418 ^ _15452;
  wire _15454 = _5905 ^ _2247;
  wire _15455 = uncoded_block[1281] ^ uncoded_block[1286];
  wire _15456 = uncoded_block[1287] ^ uncoded_block[1293];
  wire _15457 = _15455 ^ _15456;
  wire _15458 = _15454 ^ _15457;
  wire _15459 = _6564 ^ _4536;
  wire _15460 = _11198 ^ _15459;
  wire _15461 = _15458 ^ _15460;
  wire _15462 = uncoded_block[1304] ^ uncoded_block[1307];
  wire _15463 = _15462 ^ _1480;
  wire _15464 = _1482 ^ _2261;
  wire _15465 = _15463 ^ _15464;
  wire _15466 = _2262 ^ _3029;
  wire _15467 = uncoded_block[1326] ^ uncoded_block[1331];
  wire _15468 = _4543 ^ _15467;
  wire _15469 = _15466 ^ _15468;
  wire _15470 = _15465 ^ _15469;
  wire _15471 = _15461 ^ _15470;
  wire _15472 = _7815 ^ _7206;
  wire _15473 = uncoded_block[1351] ^ uncoded_block[1354];
  wire _15474 = _11218 ^ _15473;
  wire _15475 = _15472 ^ _15474;
  wire _15476 = _12853 ^ _15475;
  wire _15477 = uncoded_block[1356] ^ uncoded_block[1359];
  wire _15478 = _15477 ^ _3045;
  wire _15479 = uncoded_block[1366] ^ uncoded_block[1373];
  wire _15480 = _15479 ^ _3054;
  wire _15481 = _15478 ^ _15480;
  wire _15482 = _3055 ^ _7219;
  wire _15483 = uncoded_block[1383] ^ uncoded_block[1388];
  wire _15484 = _15483 ^ _4568;
  wire _15485 = _15482 ^ _15484;
  wire _15486 = _15481 ^ _15485;
  wire _15487 = _15476 ^ _15486;
  wire _15488 = _15471 ^ _15487;
  wire _15489 = uncoded_block[1407] ^ uncoded_block[1410];
  wire _15490 = _3847 ^ _15489;
  wire _15491 = _4573 ^ _15490;
  wire _15492 = uncoded_block[1413] ^ uncoded_block[1415];
  wire _15493 = _15492 ^ _10118;
  wire _15494 = uncoded_block[1422] ^ uncoded_block[1426];
  wire _15495 = _9021 ^ _15494;
  wire _15496 = _15493 ^ _15495;
  wire _15497 = _15491 ^ _15496;
  wire _15498 = uncoded_block[1429] ^ uncoded_block[1431];
  wire _15499 = _15498 ^ _1540;
  wire _15500 = uncoded_block[1440] ^ uncoded_block[1446];
  wire _15501 = _15500 ^ _3864;
  wire _15502 = _15499 ^ _15501;
  wire _15503 = _11246 ^ _6622;
  wire _15504 = _15503 ^ _3090;
  wire _15505 = _15502 ^ _15504;
  wire _15506 = _15497 ^ _15505;
  wire _15507 = uncoded_block[1470] ^ uncoded_block[1477];
  wire _15508 = _13440 ^ _15507;
  wire _15509 = _15508 ^ _1560;
  wire _15510 = uncoded_block[1488] ^ uncoded_block[1493];
  wire _15511 = _5988 ^ _15510;
  wire _15512 = _3890 ^ _2352;
  wire _15513 = _15511 ^ _15512;
  wire _15514 = _15509 ^ _15513;
  wire _15515 = uncoded_block[1501] ^ uncoded_block[1505];
  wire _15516 = _747 ^ _15515;
  wire _15517 = _1578 ^ _15004;
  wire _15518 = _15516 ^ _15517;
  wire _15519 = _7269 ^ _3905;
  wire _15520 = _4632 ^ _7883;
  wire _15521 = _15519 ^ _15520;
  wire _15522 = _15518 ^ _15521;
  wire _15523 = _15514 ^ _15522;
  wire _15524 = _15506 ^ _15523;
  wire _15525 = _15488 ^ _15524;
  wire _15526 = _15453 ^ _15525;
  wire _15527 = _5355 ^ _13471;
  wire _15528 = uncoded_block[1554] ^ uncoded_block[1557];
  wire _15529 = _15020 ^ _15528;
  wire _15530 = _15527 ^ _15529;
  wire _15531 = _773 ^ _7889;
  wire _15532 = _11284 ^ _9080;
  wire _15533 = _15531 ^ _15532;
  wire _15534 = _15530 ^ _15533;
  wire _15535 = uncoded_block[1576] ^ uncoded_block[1578];
  wire _15536 = _15535 ^ _2383;
  wire _15537 = uncoded_block[1583] ^ uncoded_block[1585];
  wire _15538 = uncoded_block[1587] ^ uncoded_block[1590];
  wire _15539 = _15537 ^ _15538;
  wire _15540 = _15536 ^ _15539;
  wire _15541 = uncoded_block[1593] ^ uncoded_block[1597];
  wire _15542 = _3146 ^ _15541;
  wire _15543 = _11295 ^ _3936;
  wire _15544 = _15542 ^ _15543;
  wire _15545 = _15540 ^ _15544;
  wire _15546 = _15534 ^ _15545;
  wire _15547 = _7906 ^ _6679;
  wire _15548 = _9094 ^ _7912;
  wire _15549 = _15547 ^ _15548;
  wire _15550 = _3941 ^ _807;
  wire _15551 = uncoded_block[1629] ^ uncoded_block[1632];
  wire _15552 = _14525 ^ _15551;
  wire _15553 = _15550 ^ _15552;
  wire _15554 = _15549 ^ _15553;
  wire _15555 = uncoded_block[1638] ^ uncoded_block[1640];
  wire _15556 = _7306 ^ _15555;
  wire _15557 = _2408 ^ _1647;
  wire _15558 = _15556 ^ _15557;
  wire _15559 = uncoded_block[1651] ^ uncoded_block[1654];
  wire _15560 = _9661 ^ _15559;
  wire _15561 = _3174 ^ _12960;
  wire _15562 = _15560 ^ _15561;
  wire _15563 = _15558 ^ _15562;
  wire _15564 = _15554 ^ _15563;
  wire _15565 = _15546 ^ _15564;
  wire _15566 = uncoded_block[1665] ^ uncoded_block[1669];
  wire _15567 = _15566 ^ _3182;
  wire _15568 = _15567 ^ _6702;
  wire _15569 = _10766 ^ _13519;
  wire _15570 = _6707 ^ _5409;
  wire _15571 = _15569 ^ _15570;
  wire _15572 = _15568 ^ _15571;
  wire _15573 = _2435 ^ _11879;
  wire _15574 = _3977 ^ _15573;
  wire _15575 = _3200 ^ _12976;
  wire _15576 = _15575 ^ uncoded_block[1722];
  wire _15577 = _15574 ^ _15576;
  wire _15578 = _15572 ^ _15577;
  wire _15579 = _15565 ^ _15578;
  wire _15580 = _15526 ^ _15579;
  wire _15581 = _15382 ^ _15580;
  wire _15582 = uncoded_block[2] ^ uncoded_block[7];
  wire _15583 = _15582 ^ _3995;
  wire _15584 = _4713 ^ _868;
  wire _15585 = _15583 ^ _15584;
  wire _15586 = _871 ^ _3217;
  wire _15587 = _15586 ^ _4002;
  wire _15588 = _15585 ^ _15587;
  wire _15589 = _11890 ^ _3225;
  wire _15590 = uncoded_block[36] ^ uncoded_block[38];
  wire _15591 = uncoded_block[41] ^ uncoded_block[44];
  wire _15592 = _15590 ^ _15591;
  wire _15593 = _15589 ^ _15592;
  wire _15594 = uncoded_block[45] ^ uncoded_block[47];
  wire _15595 = _15594 ^ _1699;
  wire _15596 = _10238 ^ _11899;
  wire _15597 = _15595 ^ _15596;
  wire _15598 = _15593 ^ _15597;
  wire _15599 = _15588 ^ _15598;
  wire _15600 = _32 ^ _12436;
  wire _15601 = _10244 ^ _901;
  wire _15602 = _15600 ^ _15601;
  wire _15603 = uncoded_block[89] ^ uncoded_block[90];
  wire _15604 = _11905 ^ _15603;
  wire _15605 = _8567 ^ _12443;
  wire _15606 = _15604 ^ _15605;
  wire _15607 = _15602 ^ _15606;
  wire _15608 = _4745 ^ _49;
  wire _15609 = uncoded_block[108] ^ uncoded_block[112];
  wire _15610 = _2490 ^ _15609;
  wire _15611 = _15608 ^ _15610;
  wire _15612 = _3253 ^ _54;
  wire _15613 = _1729 ^ _10821;
  wire _15614 = _15612 ^ _15613;
  wire _15615 = _15611 ^ _15614;
  wire _15616 = _15607 ^ _15615;
  wire _15617 = _15599 ^ _15616;
  wire _15618 = _1730 ^ _6774;
  wire _15619 = _15618 ^ _10260;
  wire _15620 = uncoded_block[139] ^ uncoded_block[143];
  wire _15621 = _15620 ^ _1742;
  wire _15622 = uncoded_block[148] ^ uncoded_block[150];
  wire _15623 = uncoded_block[151] ^ uncoded_block[153];
  wire _15624 = _15622 ^ _15623;
  wire _15625 = _15621 ^ _15624;
  wire _15626 = _15619 ^ _15625;
  wire _15627 = uncoded_block[159] ^ uncoded_block[165];
  wire _15628 = _15627 ^ _79;
  wire _15629 = _7398 ^ _15628;
  wire _15630 = _82 ^ _85;
  wire _15631 = uncoded_block[185] ^ uncoded_block[189];
  wire _15632 = _5479 ^ _15631;
  wire _15633 = _15630 ^ _15632;
  wire _15634 = _15629 ^ _15633;
  wire _15635 = _15626 ^ _15634;
  wire _15636 = _5483 ^ _6800;
  wire _15637 = _6801 ^ _95;
  wire _15638 = _15636 ^ _15637;
  wire _15639 = _12479 ^ _1764;
  wire _15640 = _11405 ^ _959;
  wire _15641 = _15639 ^ _15640;
  wire _15642 = _15638 ^ _15641;
  wire _15643 = _3296 ^ _1772;
  wire _15644 = uncoded_block[220] ^ uncoded_block[223];
  wire _15645 = uncoded_block[224] ^ uncoded_block[229];
  wire _15646 = _15644 ^ _15645;
  wire _15647 = _15643 ^ _15646;
  wire _15648 = _7422 ^ _112;
  wire _15649 = uncoded_block[246] ^ uncoded_block[252];
  wire _15650 = _6179 ^ _15649;
  wire _15651 = _15648 ^ _15650;
  wire _15652 = _15647 ^ _15651;
  wire _15653 = _15642 ^ _15652;
  wire _15654 = _15635 ^ _15653;
  wire _15655 = _15617 ^ _15654;
  wire _15656 = uncoded_block[253] ^ uncoded_block[256];
  wire _15657 = uncoded_block[257] ^ uncoded_block[262];
  wire _15658 = _15656 ^ _15657;
  wire _15659 = _984 ^ _7441;
  wire _15660 = _15658 ^ _15659;
  wire _15661 = _5513 ^ _5515;
  wire _15662 = _11428 ^ _992;
  wire _15663 = _15661 ^ _15662;
  wire _15664 = _15660 ^ _15663;
  wire _15665 = uncoded_block[292] ^ uncoded_block[295];
  wire _15666 = _10876 ^ _15665;
  wire _15667 = _15666 ^ _15162;
  wire _15668 = uncoded_block[307] ^ uncoded_block[309];
  wire _15669 = _4826 ^ _15668;
  wire _15670 = uncoded_block[311] ^ uncoded_block[312];
  wire _15671 = uncoded_block[313] ^ uncoded_block[315];
  wire _15672 = _15670 ^ _15671;
  wire _15673 = _15669 ^ _15672;
  wire _15674 = _15667 ^ _15673;
  wire _15675 = _15664 ^ _15674;
  wire _15676 = _4830 ^ _1008;
  wire _15677 = uncoded_block[322] ^ uncoded_block[324];
  wire _15678 = _15677 ^ _152;
  wire _15679 = _15676 ^ _15678;
  wire _15680 = _8063 ^ _13629;
  wire _15681 = _9242 ^ _6859;
  wire _15682 = _15680 ^ _15681;
  wire _15683 = _15679 ^ _15682;
  wire _15684 = uncoded_block[352] ^ uncoded_block[355];
  wire _15685 = _9790 ^ _15684;
  wire _15686 = uncoded_block[357] ^ uncoded_block[362];
  wire _15687 = _15686 ^ _7470;
  wire _15688 = _15685 ^ _15687;
  wire _15689 = _8076 ^ _7474;
  wire _15690 = _1841 ^ _4858;
  wire _15691 = _15689 ^ _15690;
  wire _15692 = _15688 ^ _15691;
  wire _15693 = _15683 ^ _15692;
  wire _15694 = _15675 ^ _15693;
  wire _15695 = _12541 ^ _3384;
  wire _15696 = uncoded_block[397] ^ uncoded_block[401];
  wire _15697 = uncoded_block[403] ^ uncoded_block[405];
  wire _15698 = _15696 ^ _15697;
  wire _15699 = _15695 ^ _15698;
  wire _15700 = _184 ^ _1055;
  wire _15701 = _1854 ^ _4874;
  wire _15702 = _15700 ^ _15701;
  wire _15703 = _15699 ^ _15702;
  wire _15704 = uncoded_block[430] ^ uncoded_block[432];
  wire _15705 = _197 ^ _15704;
  wire _15706 = uncoded_block[436] ^ uncoded_block[441];
  wire _15707 = _10352 ^ _15706;
  wire _15708 = _15705 ^ _15707;
  wire _15709 = uncoded_block[442] ^ uncoded_block[447];
  wire _15710 = _15709 ^ _4176;
  wire _15711 = _212 ^ _1871;
  wire _15712 = _15710 ^ _15711;
  wire _15713 = _15708 ^ _15712;
  wire _15714 = _15703 ^ _15713;
  wire _15715 = uncoded_block[461] ^ uncoded_block[463];
  wire _15716 = _15715 ^ _8683;
  wire _15717 = _9283 ^ _221;
  wire _15718 = _15716 ^ _15717;
  wire _15719 = uncoded_block[476] ^ uncoded_block[480];
  wire _15720 = _15719 ^ _4895;
  wire _15721 = uncoded_block[483] ^ uncoded_block[494];
  wire _15722 = _15721 ^ _13139;
  wire _15723 = _15720 ^ _15722;
  wire _15724 = _15718 ^ _15723;
  wire _15725 = uncoded_block[501] ^ uncoded_block[507];
  wire _15726 = _228 ^ _15725;
  wire _15727 = _15726 ^ _7532;
  wire _15728 = _9840 ^ _8708;
  wire _15729 = _10948 ^ _14716;
  wire _15730 = _15728 ^ _15729;
  wire _15731 = _15727 ^ _15730;
  wire _15732 = _15724 ^ _15731;
  wire _15733 = _15714 ^ _15732;
  wire _15734 = _15694 ^ _15733;
  wire _15735 = _15655 ^ _15734;
  wire _15736 = _1111 ^ _4926;
  wire _15737 = _7536 ^ _6298;
  wire _15738 = _15736 ^ _15737;
  wire _15739 = _4931 ^ _4933;
  wire _15740 = uncoded_block[555] ^ uncoded_block[557];
  wire _15741 = _15236 ^ _15740;
  wire _15742 = _15739 ^ _15741;
  wire _15743 = _15738 ^ _15742;
  wire _15744 = _3461 ^ _3465;
  wire _15745 = _259 ^ _1931;
  wire _15746 = _15744 ^ _15745;
  wire _15747 = uncoded_block[579] ^ uncoded_block[580];
  wire _15748 = _263 ^ _15747;
  wire _15749 = _5641 ^ _1139;
  wire _15750 = _15748 ^ _15749;
  wire _15751 = _15746 ^ _15750;
  wire _15752 = _15743 ^ _15751;
  wire _15753 = _271 ^ _1938;
  wire _15754 = uncoded_block[595] ^ uncoded_block[600];
  wire _15755 = _15754 ^ _5646;
  wire _15756 = _15753 ^ _15755;
  wire _15757 = uncoded_block[604] ^ uncoded_block[608];
  wire _15758 = uncoded_block[612] ^ uncoded_block[615];
  wire _15759 = _15757 ^ _15758;
  wire _15760 = _4243 ^ _10418;
  wire _15761 = _15759 ^ _15760;
  wire _15762 = _15756 ^ _15761;
  wire _15763 = _8161 ^ _12075;
  wire _15764 = _11543 ^ _296;
  wire _15765 = _15763 ^ _15764;
  wire _15766 = uncoded_block[647] ^ uncoded_block[649];
  wire _15767 = _15766 ^ _1170;
  wire _15768 = uncoded_block[661] ^ uncoded_block[662];
  wire _15769 = _2738 ^ _15768;
  wire _15770 = _15767 ^ _15769;
  wire _15771 = _15765 ^ _15770;
  wire _15772 = _15762 ^ _15771;
  wire _15773 = _15752 ^ _15772;
  wire _15774 = uncoded_block[663] ^ uncoded_block[669];
  wire _15775 = uncoded_block[672] ^ uncoded_block[674];
  wire _15776 = _15774 ^ _15775;
  wire _15777 = _15281 ^ _2751;
  wire _15778 = _15776 ^ _15777;
  wire _15779 = _2754 ^ _3529;
  wire _15780 = _3532 ^ _14250;
  wire _15781 = _15779 ^ _15780;
  wire _15782 = _15778 ^ _15781;
  wire _15783 = uncoded_block[706] ^ uncoded_block[709];
  wire _15784 = _15783 ^ _1192;
  wire _15785 = uncoded_block[713] ^ uncoded_block[720];
  wire _15786 = _15785 ^ _1988;
  wire _15787 = _15784 ^ _15786;
  wire _15788 = uncoded_block[733] ^ uncoded_block[736];
  wire _15789 = _8200 ^ _15788;
  wire _15790 = _7005 ^ _5699;
  wire _15791 = _15789 ^ _15790;
  wire _15792 = _15787 ^ _15791;
  wire _15793 = _15782 ^ _15792;
  wire _15794 = _5702 ^ _8209;
  wire _15795 = uncoded_block[757] ^ uncoded_block[761];
  wire _15796 = _11012 ^ _15795;
  wire _15797 = _15794 ^ _15796;
  wire _15798 = _13762 ^ _10470;
  wire _15799 = uncoded_block[772] ^ uncoded_block[774];
  wire _15800 = _1218 ^ _15799;
  wire _15801 = _15798 ^ _15800;
  wire _15802 = _15797 ^ _15801;
  wire _15803 = _9382 ^ _9384;
  wire _15804 = _4309 ^ _6388;
  wire _15805 = _15803 ^ _15804;
  wire _15806 = _2019 ^ _1232;
  wire _15807 = _6391 ^ _8223;
  wire _15808 = _15806 ^ _15807;
  wire _15809 = _15805 ^ _15808;
  wire _15810 = _15802 ^ _15809;
  wire _15811 = _15793 ^ _15810;
  wire _15812 = _15773 ^ _15811;
  wire _15813 = _7029 ^ _4317;
  wire _15814 = uncoded_block[807] ^ uncoded_block[809];
  wire _15815 = _3577 ^ _15814;
  wire _15816 = _15813 ^ _15815;
  wire _15817 = _11596 ^ _5046;
  wire _15818 = _15320 ^ _5052;
  wire _15819 = _15817 ^ _15818;
  wire _15820 = _15816 ^ _15819;
  wire _15821 = _1253 ^ _5057;
  wire _15822 = _1262 ^ _3600;
  wire _15823 = _15821 ^ _15822;
  wire _15824 = uncoded_block[859] ^ uncoded_block[863];
  wire _15825 = _15824 ^ _1266;
  wire _15826 = uncoded_block[872] ^ uncoded_block[875];
  wire _15827 = _5072 ^ _15826;
  wire _15828 = _15825 ^ _15827;
  wire _15829 = _15823 ^ _15828;
  wire _15830 = _15820 ^ _15829;
  wire _15831 = _420 ^ _2836;
  wire _15832 = _423 ^ _2059;
  wire _15833 = _15831 ^ _15832;
  wire _15834 = _12704 ^ _4355;
  wire _15835 = _15834 ^ _7067;
  wire _15836 = _15833 ^ _15835;
  wire _15837 = _15345 ^ _4361;
  wire _15838 = _1287 ^ _10513;
  wire _15839 = _15837 ^ _15838;
  wire _15840 = uncoded_block[920] ^ uncoded_block[923];
  wire _15841 = uncoded_block[925] ^ uncoded_block[928];
  wire _15842 = _15840 ^ _15841;
  wire _15843 = _1296 ^ _2078;
  wire _15844 = _15842 ^ _15843;
  wire _15845 = _15839 ^ _15844;
  wire _15846 = _15836 ^ _15845;
  wire _15847 = _15830 ^ _15846;
  wire _15848 = uncoded_block[936] ^ uncoded_block[938];
  wire _15849 = _15848 ^ _8271;
  wire _15850 = _15849 ^ _9436;
  wire _15851 = _11646 ^ _11649;
  wire _15852 = _7681 ^ _15851;
  wire _15853 = _15850 ^ _15852;
  wire _15854 = uncoded_block[975] ^ uncoded_block[980];
  wire _15855 = _15854 ^ _8287;
  wire _15856 = _10543 ^ _4402;
  wire _15857 = _15855 ^ _15856;
  wire _15858 = uncoded_block[999] ^ uncoded_block[1003];
  wire _15859 = _15858 ^ _2886;
  wire _15860 = uncoded_block[1008] ^ uncoded_block[1011];
  wire _15861 = _15860 ^ _8296;
  wire _15862 = _15859 ^ _15861;
  wire _15863 = _15857 ^ _15862;
  wire _15864 = _15853 ^ _15863;
  wire _15865 = _12750 ^ _9454;
  wire _15866 = _8874 ^ _4417;
  wire _15867 = _15865 ^ _15866;
  wire _15868 = _10555 ^ _1348;
  wire _15869 = _15867 ^ _15868;
  wire _15870 = _3681 ^ _1357;
  wire _15871 = uncoded_block[1051] ^ uncoded_block[1055];
  wire _15872 = _15871 ^ _5816;
  wire _15873 = _15870 ^ _15872;
  wire _15874 = _3689 ^ _2143;
  wire _15875 = _5827 ^ _15874;
  wire _15876 = _15873 ^ _15875;
  wire _15877 = _15869 ^ _15876;
  wire _15878 = _15864 ^ _15877;
  wire _15879 = _15847 ^ _15878;
  wire _15880 = _15812 ^ _15879;
  wire _15881 = _15735 ^ _15880;
  wire _15882 = _5831 ^ _6486;
  wire _15883 = uncoded_block[1078] ^ uncoded_block[1083];
  wire _15884 = _15883 ^ _1373;
  wire _15885 = _15882 ^ _15884;
  wire _15886 = _1374 ^ _10021;
  wire _15887 = _542 ^ _3708;
  wire _15888 = _15886 ^ _15887;
  wire _15889 = _15885 ^ _15888;
  wire _15890 = uncoded_block[1112] ^ uncoded_block[1116];
  wire _15891 = _7132 ^ _15890;
  wire _15892 = _5853 ^ _8342;
  wire _15893 = _15891 ^ _15892;
  wire _15894 = uncoded_block[1127] ^ uncoded_block[1128];
  wire _15895 = _15894 ^ _8343;
  wire _15896 = uncoded_block[1133] ^ uncoded_block[1134];
  wire _15897 = _15896 ^ _9496;
  wire _15898 = _15895 ^ _15897;
  wire _15899 = _15893 ^ _15898;
  wire _15900 = _15889 ^ _15899;
  wire _15901 = _5859 ^ _2953;
  wire _15902 = uncoded_block[1148] ^ uncoded_block[1151];
  wire _15903 = _15902 ^ _4468;
  wire _15904 = _15901 ^ _15903;
  wire _15905 = uncoded_block[1154] ^ uncoded_block[1162];
  wire _15906 = _15905 ^ _6511;
  wire _15907 = uncoded_block[1166] ^ uncoded_block[1168];
  wire _15908 = _15907 ^ _7154;
  wire _15909 = _15906 ^ _15908;
  wire _15910 = _15904 ^ _15909;
  wire _15911 = _2967 ^ _2193;
  wire _15912 = _2195 ^ _5200;
  wire _15913 = _15911 ^ _15912;
  wire _15914 = _2200 ^ _4488;
  wire _15915 = _5883 ^ _5209;
  wire _15916 = _15914 ^ _15915;
  wire _15917 = _15913 ^ _15916;
  wire _15918 = _15910 ^ _15917;
  wire _15919 = _15900 ^ _15918;
  wire _15920 = _10617 ^ _3762;
  wire _15921 = uncoded_block[1217] ^ uncoded_block[1221];
  wire _15922 = _2219 ^ _15921;
  wire _15923 = _15920 ^ _15922;
  wire _15924 = uncoded_block[1222] ^ uncoded_block[1226];
  wire _15925 = _15924 ^ _5894;
  wire _15926 = uncoded_block[1231] ^ uncoded_block[1234];
  wire _15927 = uncoded_block[1235] ^ uncoded_block[1237];
  wire _15928 = _15926 ^ _15927;
  wire _15929 = _15925 ^ _15928;
  wire _15930 = _15923 ^ _15929;
  wire _15931 = _2230 ^ _2995;
  wire _15932 = _3777 ^ _4511;
  wire _15933 = _15931 ^ _15932;
  wire _15934 = uncoded_block[1254] ^ uncoded_block[1257];
  wire _15935 = _7778 ^ _15934;
  wire _15936 = _12825 ^ _5235;
  wire _15937 = _15935 ^ _15936;
  wire _15938 = _15933 ^ _15937;
  wire _15939 = _15930 ^ _15938;
  wire _15940 = _6550 ^ _11188;
  wire _15941 = _9538 ^ _630;
  wire _15942 = _15940 ^ _15941;
  wire _15943 = _6556 ^ _4526;
  wire _15944 = _8980 ^ _3800;
  wire _15945 = _15943 ^ _15944;
  wire _15946 = _15942 ^ _15945;
  wire _15947 = _3801 ^ _1471;
  wire _15948 = _1472 ^ _3025;
  wire _15949 = _15947 ^ _15948;
  wire _15950 = _5919 ^ _2262;
  wire _15951 = uncoded_block[1318] ^ uncoded_block[1322];
  wire _15952 = _15951 ^ _8411;
  wire _15953 = _15950 ^ _15952;
  wire _15954 = _15949 ^ _15953;
  wire _15955 = _15946 ^ _15954;
  wire _15956 = _15939 ^ _15955;
  wire _15957 = _15919 ^ _15956;
  wire _15958 = uncoded_block[1329] ^ uncoded_block[1339];
  wire _15959 = _15958 ^ _5262;
  wire _15960 = _15473 ^ _12300;
  wire _15961 = _15959 ^ _15960;
  wire _15962 = uncoded_block[1363] ^ uncoded_block[1366];
  wire _15963 = _15962 ^ _12302;
  wire _15964 = _15963 ^ _3053;
  wire _15965 = _15961 ^ _15964;
  wire _15966 = uncoded_block[1375] ^ uncoded_block[1378];
  wire _15967 = _15966 ^ _13410;
  wire _15968 = _5950 ^ _1513;
  wire _15969 = _15967 ^ _15968;
  wire _15970 = uncoded_block[1393] ^ uncoded_block[1400];
  wire _15971 = _15970 ^ _1519;
  wire _15972 = uncoded_block[1412] ^ uncoded_block[1415];
  wire _15973 = _5961 ^ _15972;
  wire _15974 = _15971 ^ _15973;
  wire _15975 = _15969 ^ _15974;
  wire _15976 = _15965 ^ _15975;
  wire _15977 = _705 ^ _10120;
  wire _15978 = _9588 ^ _2311;
  wire _15979 = _15977 ^ _15978;
  wire _15980 = uncoded_block[1429] ^ uncoded_block[1432];
  wire _15981 = _15980 ^ _1534;
  wire _15982 = uncoded_block[1436] ^ uncoded_block[1440];
  wire _15983 = _15982 ^ _12330;
  wire _15984 = _15981 ^ _15983;
  wire _15985 = _15979 ^ _15984;
  wire _15986 = _2325 ^ _2328;
  wire _15987 = _9037 ^ _3870;
  wire _15988 = _15986 ^ _15987;
  wire _15989 = _3094 ^ _2338;
  wire _15990 = _15989 ^ _11803;
  wire _15991 = _15988 ^ _15990;
  wire _15992 = _15985 ^ _15991;
  wire _15993 = _15976 ^ _15992;
  wire _15994 = uncoded_block[1480] ^ uncoded_block[1483];
  wire _15995 = _15994 ^ _2349;
  wire _15996 = uncoded_block[1489] ^ uncoded_block[1493];
  wire _15997 = _15996 ^ _12898;
  wire _15998 = _15995 ^ _15997;
  wire _15999 = uncoded_block[1501] ^ uncoded_block[1507];
  wire _16000 = _747 ^ _15999;
  wire _16001 = _750 ^ _9053;
  wire _16002 = _16000 ^ _16001;
  wire _16003 = _15998 ^ _16002;
  wire _16004 = uncoded_block[1514] ^ uncoded_block[1516];
  wire _16005 = _16004 ^ _15004;
  wire _16006 = _755 ^ _2360;
  wire _16007 = _16005 ^ _16006;
  wire _16008 = uncoded_block[1532] ^ uncoded_block[1535];
  wire _16009 = _16008 ^ _15009;
  wire _16010 = uncoded_block[1539] ^ uncoded_block[1542];
  wire _16011 = _16010 ^ _5355;
  wire _16012 = _16009 ^ _16011;
  wire _16013 = _16007 ^ _16012;
  wire _16014 = _16003 ^ _16013;
  wire _16015 = _7275 ^ _767;
  wire _16016 = uncoded_block[1554] ^ uncoded_block[1558];
  wire _16017 = _16016 ^ _4640;
  wire _16018 = _16015 ^ _16017;
  wire _16019 = uncoded_block[1563] ^ uncoded_block[1567];
  wire _16020 = uncoded_block[1570] ^ uncoded_block[1573];
  wire _16021 = _16019 ^ _16020;
  wire _16022 = _2383 ^ _12369;
  wire _16023 = _16021 ^ _16022;
  wire _16024 = _16018 ^ _16023;
  wire _16025 = uncoded_block[1585] ^ uncoded_block[1591];
  wire _16026 = uncoded_block[1592] ^ uncoded_block[1598];
  wire _16027 = _16025 ^ _16026;
  wire _16028 = _5373 ^ _12373;
  wire _16029 = _16027 ^ _16028;
  wire _16030 = _2396 ^ _5380;
  wire _16031 = uncoded_block[1611] ^ uncoded_block[1614];
  wire _16032 = uncoded_block[1616] ^ uncoded_block[1617];
  wire _16033 = _16031 ^ _16032;
  wire _16034 = _16030 ^ _16033;
  wire _16035 = _16029 ^ _16034;
  wire _16036 = _16024 ^ _16035;
  wire _16037 = _16014 ^ _16036;
  wire _16038 = _15993 ^ _16037;
  wire _16039 = _15957 ^ _16038;
  wire _16040 = _6684 ^ _14525;
  wire _16041 = _2404 ^ _9099;
  wire _16042 = _16040 ^ _16041;
  wire _16043 = _6689 ^ _13500;
  wire _16044 = _5394 ^ _12386;
  wire _16045 = _16043 ^ _16044;
  wire _16046 = _16042 ^ _16045;
  wire _16047 = uncoded_block[1648] ^ uncoded_block[1655];
  wire _16048 = _16047 ^ _13508;
  wire _16049 = uncoded_block[1662] ^ uncoded_block[1664];
  wire _16050 = _4680 ^ _16049;
  wire _16051 = _16048 ^ _16050;
  wire _16052 = uncoded_block[1668] ^ uncoded_block[1670];
  wire _16053 = _7319 ^ _16052;
  wire _16054 = _6700 ^ _5406;
  wire _16055 = _16053 ^ _16054;
  wire _16056 = _16051 ^ _16055;
  wire _16057 = _16046 ^ _16056;
  wire _16058 = uncoded_block[1683] ^ uncoded_block[1686];
  wire _16059 = _16058 ^ _3189;
  wire _16060 = uncoded_block[1691] ^ uncoded_block[1694];
  wire _16061 = uncoded_block[1698] ^ uncoded_block[1704];
  wire _16062 = _16060 ^ _16061;
  wire _16063 = _16059 ^ _16062;
  wire _16064 = uncoded_block[1706] ^ uncoded_block[1710];
  wire _16065 = uncoded_block[1712] ^ uncoded_block[1718];
  wire _16066 = _16064 ^ _16065;
  wire _16067 = _16066 ^ uncoded_block[1719];
  wire _16068 = _16063 ^ _16067;
  wire _16069 = _16057 ^ _16068;
  wire _16070 = _16039 ^ _16069;
  wire _16071 = _15881 ^ _16070;
  wire _16072 = _3993 ^ _4;
  wire _16073 = _7953 ^ _16072;
  wire _16074 = _4716 ^ _1690;
  wire _16075 = _5424 ^ _16074;
  wire _16076 = _16073 ^ _16075;
  wire _16077 = _6728 ^ _3225;
  wire _16078 = _11347 ^ _19;
  wire _16079 = _16077 ^ _16078;
  wire _16080 = _4008 ^ _10234;
  wire _16081 = _16080 ^ _10236;
  wire _16082 = _16079 ^ _16081;
  wire _16083 = _16076 ^ _16082;
  wire _16084 = uncoded_block[54] ^ uncoded_block[64];
  wire _16085 = uncoded_block[66] ^ uncoded_block[69];
  wire _16086 = _16084 ^ _16085;
  wire _16087 = _7976 ^ _900;
  wire _16088 = _16086 ^ _16087;
  wire _16089 = uncoded_block[79] ^ uncoded_block[86];
  wire _16090 = _901 ^ _16089;
  wire _16091 = uncoded_block[90] ^ uncoded_block[97];
  wire _16092 = _16091 ^ _11909;
  wire _16093 = _16090 ^ _16092;
  wire _16094 = _16088 ^ _16093;
  wire _16095 = _1726 ^ _6769;
  wire _16096 = _1723 ^ _16095;
  wire _16097 = uncoded_block[122] ^ uncoded_block[126];
  wire _16098 = _9721 ^ _16097;
  wire _16099 = _6774 ^ _1735;
  wire _16100 = _16098 ^ _16099;
  wire _16101 = _16096 ^ _16100;
  wire _16102 = _16094 ^ _16101;
  wire _16103 = _16083 ^ _16102;
  wire _16104 = uncoded_block[139] ^ uncoded_block[148];
  wire _16105 = _16104 ^ _1744;
  wire _16106 = _10260 ^ _16105;
  wire _16107 = _15623 ^ _3271;
  wire _16108 = _6785 ^ _4054;
  wire _16109 = _16107 ^ _16108;
  wire _16110 = _16106 ^ _16109;
  wire _16111 = _2522 ^ _82;
  wire _16112 = _7403 ^ _10843;
  wire _16113 = _16111 ^ _16112;
  wire _16114 = uncoded_block[185] ^ uncoded_block[188];
  wire _16115 = _16114 ^ _6155;
  wire _16116 = uncoded_block[197] ^ uncoded_block[198];
  wire _16117 = _16116 ^ _2537;
  wire _16118 = _16115 ^ _16117;
  wire _16119 = _16113 ^ _16118;
  wire _16120 = _16110 ^ _16119;
  wire _16121 = _8021 ^ _1766;
  wire _16122 = _959 ^ _3296;
  wire _16123 = _16121 ^ _16122;
  wire _16124 = _4787 ^ _5498;
  wire _16125 = uncoded_block[229] ^ uncoded_block[232];
  wire _16126 = _16125 ^ _2550;
  wire _16127 = _16124 ^ _16126;
  wire _16128 = _16123 ^ _16127;
  wire _16129 = uncoded_block[244] ^ uncoded_block[248];
  wire _16130 = _16129 ^ _11954;
  wire _16131 = _15145 ^ _16130;
  wire _16132 = _4803 ^ _4088;
  wire _16133 = _14641 ^ _984;
  wire _16134 = _16132 ^ _16133;
  wire _16135 = _16131 ^ _16134;
  wire _16136 = _16128 ^ _16135;
  wire _16137 = _16120 ^ _16136;
  wire _16138 = _16103 ^ _16137;
  wire _16139 = _14642 ^ _10872;
  wire _16140 = _2568 ^ _7445;
  wire _16141 = _16139 ^ _16140;
  wire _16142 = uncoded_block[281] ^ uncoded_block[285];
  wire _16143 = _16142 ^ _992;
  wire _16144 = uncoded_block[291] ^ uncoded_block[294];
  wire _16145 = _16144 ^ _137;
  wire _16146 = _16143 ^ _16145;
  wire _16147 = _16141 ^ _16146;
  wire _16148 = _1810 ^ _4826;
  wire _16149 = uncoded_block[314] ^ uncoded_block[318];
  wire _16150 = _6845 ^ _16149;
  wire _16151 = _16148 ^ _16150;
  wire _16152 = _1818 ^ _3347;
  wire _16153 = _11444 ^ _11983;
  wire _16154 = _16152 ^ _16153;
  wire _16155 = _16151 ^ _16154;
  wire _16156 = _16147 ^ _16155;
  wire _16157 = _4838 ^ _1825;
  wire _16158 = uncoded_block[343] ^ uncoded_block[345];
  wire _16159 = _6217 ^ _16158;
  wire _16160 = _16157 ^ _16159;
  wire _16161 = uncoded_block[346] ^ uncoded_block[349];
  wire _16162 = _16161 ^ _1028;
  wire _16163 = _3361 ^ _6227;
  wire _16164 = _16162 ^ _16163;
  wire _16165 = _16160 ^ _16164;
  wire _16166 = _7470 ^ _169;
  wire _16167 = _4141 ^ _12538;
  wire _16168 = _16166 ^ _16167;
  wire _16169 = uncoded_block[383] ^ uncoded_block[387];
  wire _16170 = _16169 ^ _6239;
  wire _16171 = _5554 ^ _177;
  wire _16172 = _16170 ^ _16171;
  wire _16173 = _16168 ^ _16172;
  wire _16174 = _16165 ^ _16173;
  wire _16175 = _16156 ^ _16174;
  wire _16176 = _10910 ^ _4155;
  wire _16177 = uncoded_block[404] ^ uncoded_block[407];
  wire _16178 = _16177 ^ _10344;
  wire _16179 = _16176 ^ _16178;
  wire _16180 = _2630 ^ _3396;
  wire _16181 = _4872 ^ _4874;
  wire _16182 = _16180 ^ _16181;
  wire _16183 = _16179 ^ _16182;
  wire _16184 = uncoded_block[428] ^ uncoded_block[431];
  wire _16185 = _1062 ^ _16184;
  wire _16186 = uncoded_block[432] ^ uncoded_block[436];
  wire _16187 = uncoded_block[437] ^ uncoded_block[439];
  wire _16188 = _16186 ^ _16187;
  wire _16189 = _16185 ^ _16188;
  wire _16190 = uncoded_block[441] ^ uncoded_block[444];
  wire _16191 = uncoded_block[445] ^ uncoded_block[448];
  wire _16192 = _16190 ^ _16191;
  wire _16193 = _213 ^ _15715;
  wire _16194 = _16192 ^ _16193;
  wire _16195 = _16189 ^ _16194;
  wire _16196 = _16183 ^ _16195;
  wire _16197 = _4890 ^ _9283;
  wire _16198 = _11494 ^ _5593;
  wire _16199 = _16197 ^ _16198;
  wire _16200 = uncoded_block[484] ^ uncoded_block[489];
  wire _16201 = _1086 ^ _16200;
  wire _16202 = _16201 ^ _9836;
  wire _16203 = _16199 ^ _16202;
  wire _16204 = _9837 ^ _3434;
  wire _16205 = _16204 ^ _7530;
  wire _16206 = uncoded_block[517] ^ uncoded_block[524];
  wire _16207 = _8706 ^ _16206;
  wire _16208 = _14192 ^ _16207;
  wire _16209 = _16205 ^ _16208;
  wire _16210 = _16203 ^ _16209;
  wire _16211 = _16196 ^ _16210;
  wire _16212 = _16175 ^ _16211;
  wire _16213 = _16138 ^ _16212;
  wire _16214 = _1900 ^ _6929;
  wire _16215 = uncoded_block[533] ^ uncoded_block[534];
  wire _16216 = _1111 ^ _16215;
  wire _16217 = _16214 ^ _16216;
  wire _16218 = _10961 ^ _15236;
  wire _16219 = _1910 ^ _16218;
  wire _16220 = _16217 ^ _16219;
  wire _16221 = _15740 ^ _8139;
  wire _16222 = _9319 ^ _4940;
  wire _16223 = _16221 ^ _16222;
  wire _16224 = _6942 ^ _14209;
  wire _16225 = _10400 ^ _9325;
  wire _16226 = _16224 ^ _16225;
  wire _16227 = _16223 ^ _16226;
  wire _16228 = _16220 ^ _16227;
  wire _16229 = _1139 ^ _4950;
  wire _16230 = _4234 ^ _1938;
  wire _16231 = _16229 ^ _16230;
  wire _16232 = _8149 ^ _15252;
  wire _16233 = uncoded_block[607] ^ uncoded_block[609];
  wire _16234 = _8152 ^ _16233;
  wire _16235 = _16232 ^ _16234;
  wire _16236 = _16231 ^ _16235;
  wire _16237 = _8154 ^ _7563;
  wire _16238 = uncoded_block[615] ^ uncoded_block[619];
  wire _16239 = _16238 ^ _4246;
  wire _16240 = _16237 ^ _16239;
  wire _16241 = uncoded_block[640] ^ uncoded_block[643];
  wire _16242 = _16241 ^ _296;
  wire _16243 = _7578 ^ _16242;
  wire _16244 = _16240 ^ _16243;
  wire _16245 = _16236 ^ _16244;
  wire _16246 = _16228 ^ _16245;
  wire _16247 = uncoded_block[647] ^ uncoded_block[651];
  wire _16248 = _16247 ^ _302;
  wire _16249 = uncoded_block[655] ^ uncoded_block[656];
  wire _16250 = _16249 ^ _2739;
  wire _16251 = _16248 ^ _16250;
  wire _16252 = uncoded_block[662] ^ uncoded_block[668];
  wire _16253 = _16252 ^ _311;
  wire _16254 = _312 ^ _8760;
  wire _16255 = _16253 ^ _16254;
  wire _16256 = _16251 ^ _16255;
  wire _16257 = _13731 ^ _6352;
  wire _16258 = uncoded_block[681] ^ uncoded_block[689];
  wire _16259 = _16258 ^ _4272;
  wire _16260 = _16257 ^ _16259;
  wire _16261 = _11557 ^ _11562;
  wire _16262 = uncoded_block[703] ^ uncoded_block[709];
  wire _16263 = _6992 ^ _16262;
  wire _16264 = _16261 ^ _16263;
  wire _16265 = _16260 ^ _16264;
  wire _16266 = _16256 ^ _16265;
  wire _16267 = _1192 ^ _5002;
  wire _16268 = _16267 ^ _1989;
  wire _16269 = _10457 ^ _349;
  wire _16270 = _1995 ^ _13208;
  wire _16271 = _16269 ^ _16270;
  wire _16272 = _16268 ^ _16271;
  wire _16273 = uncoded_block[747] ^ uncoded_block[754];
  wire _16274 = _16273 ^ _15795;
  wire _16275 = _16274 ^ _15798;
  wire _16276 = _11019 ^ _13216;
  wire _16277 = _3562 ^ _3567;
  wire _16278 = _16276 ^ _16277;
  wire _16279 = _16275 ^ _16278;
  wire _16280 = _16272 ^ _16279;
  wire _16281 = _16266 ^ _16280;
  wire _16282 = _16246 ^ _16281;
  wire _16283 = _3570 ^ _8790;
  wire _16284 = _7626 ^ _2799;
  wire _16285 = _16283 ^ _16284;
  wire _16286 = _6391 ^ _7029;
  wire _16287 = _1235 ^ _390;
  wire _16288 = _16286 ^ _16287;
  wire _16289 = _16285 ^ _16288;
  wire _16290 = _2026 ^ _6398;
  wire _16291 = _7037 ^ _1247;
  wire _16292 = _16290 ^ _16291;
  wire _16293 = uncoded_block[834] ^ uncoded_block[837];
  wire _16294 = _16293 ^ _4339;
  wire _16295 = uncoded_block[849] ^ uncoded_block[855];
  wire _16296 = _405 ^ _16295;
  wire _16297 = _16294 ^ _16296;
  wire _16298 = _16292 ^ _16297;
  wire _16299 = _16289 ^ _16298;
  wire _16300 = uncoded_block[860] ^ uncoded_block[866];
  wire _16301 = _8812 ^ _16300;
  wire _16302 = _16301 ^ _14306;
  wire _16303 = uncoded_block[874] ^ uncoded_block[878];
  wire _16304 = uncoded_block[879] ^ uncoded_block[880];
  wire _16305 = _16303 ^ _16304;
  wire _16306 = _423 ^ _2061;
  wire _16307 = _16305 ^ _16306;
  wire _16308 = _16302 ^ _16307;
  wire _16309 = _2841 ^ _6424;
  wire _16310 = _1281 ^ _1284;
  wire _16311 = _16309 ^ _16310;
  wire _16312 = uncoded_block[909] ^ uncoded_block[912];
  wire _16313 = uncoded_block[913] ^ uncoded_block[916];
  wire _16314 = _16312 ^ _16313;
  wire _16315 = uncoded_block[922] ^ uncoded_block[925];
  wire _16316 = _438 ^ _16315;
  wire _16317 = _16314 ^ _16316;
  wire _16318 = _16311 ^ _16317;
  wire _16319 = _16308 ^ _16318;
  wire _16320 = _16299 ^ _16319;
  wire _16321 = uncoded_block[929] ^ uncoded_block[934];
  wire _16322 = _16321 ^ _5101;
  wire _16323 = _6439 ^ _455;
  wire _16324 = _16322 ^ _16323;
  wire _16325 = _456 ^ _5777;
  wire _16326 = uncoded_block[953] ^ uncoded_block[958];
  wire _16327 = _16326 ^ _1308;
  wire _16328 = _16325 ^ _16327;
  wire _16329 = _16324 ^ _16328;
  wire _16330 = _10529 ^ _12179;
  wire _16331 = _11087 ^ _1314;
  wire _16332 = _16330 ^ _16331;
  wire _16333 = _1315 ^ _5789;
  wire _16334 = _2100 ^ _8855;
  wire _16335 = _16333 ^ _16334;
  wire _16336 = _16332 ^ _16335;
  wire _16337 = _16329 ^ _16336;
  wire _16338 = uncoded_block[989] ^ uncoded_block[990];
  wire _16339 = _1317 ^ _16338;
  wire _16340 = _1323 ^ _10543;
  wire _16341 = _16339 ^ _16340;
  wire _16342 = _11101 ^ _7691;
  wire _16343 = uncoded_block[1003] ^ uncoded_block[1006];
  wire _16344 = _16343 ^ _4405;
  wire _16345 = _16342 ^ _16344;
  wire _16346 = _16341 ^ _16345;
  wire _16347 = _4410 ^ _10547;
  wire _16348 = _1334 ^ _8301;
  wire _16349 = _16347 ^ _16348;
  wire _16350 = _5806 ^ _2127;
  wire _16351 = _502 ^ _511;
  wire _16352 = _16350 ^ _16351;
  wire _16353 = _16349 ^ _16352;
  wire _16354 = _16346 ^ _16353;
  wire _16355 = _16337 ^ _16354;
  wire _16356 = _16320 ^ _16355;
  wire _16357 = _16282 ^ _16356;
  wire _16358 = _16213 ^ _16357;
  wire _16359 = _2133 ^ _13844;
  wire _16360 = uncoded_block[1057] ^ uncoded_block[1065];
  wire _16361 = _3682 ^ _16360;
  wire _16362 = _16359 ^ _16361;
  wire _16363 = _9475 ^ _1366;
  wire _16364 = _16363 ^ _5833;
  wire _16365 = _16362 ^ _16364;
  wire _16366 = _13311 ^ _10021;
  wire _16367 = _8905 ^ _16366;
  wire _16368 = uncoded_block[1092] ^ uncoded_block[1097];
  wire _16369 = _16368 ^ _5169;
  wire _16370 = _7731 ^ _8914;
  wire _16371 = _16369 ^ _16370;
  wire _16372 = _16367 ^ _16371;
  wire _16373 = _16365 ^ _16372;
  wire _16374 = uncoded_block[1110] ^ uncoded_block[1113];
  wire _16375 = _16374 ^ _3713;
  wire _16376 = uncoded_block[1120] ^ uncoded_block[1124];
  wire _16377 = _11147 ^ _16376;
  wire _16378 = _16375 ^ _16377;
  wire _16379 = _6499 ^ _5856;
  wire _16380 = uncoded_block[1140] ^ uncoded_block[1143];
  wire _16381 = _8346 ^ _16380;
  wire _16382 = _16379 ^ _16381;
  wire _16383 = _16378 ^ _16382;
  wire _16384 = _15902 ^ _3727;
  wire _16385 = _14389 ^ _6511;
  wire _16386 = _16384 ^ _16385;
  wire _16387 = _4476 ^ _11161;
  wire _16388 = _1410 ^ _2967;
  wire _16389 = _16387 ^ _16388;
  wire _16390 = _16386 ^ _16389;
  wire _16391 = _16383 ^ _16390;
  wire _16392 = _16373 ^ _16391;
  wire _16393 = uncoded_block[1179] ^ uncoded_block[1182];
  wire _16394 = _589 ^ _16393;
  wire _16395 = _4486 ^ _2971;
  wire _16396 = _16394 ^ _16395;
  wire _16397 = uncoded_block[1192] ^ uncoded_block[1198];
  wire _16398 = _16397 ^ _7162;
  wire _16399 = uncoded_block[1204] ^ uncoded_block[1207];
  wire _16400 = _16399 ^ _7765;
  wire _16401 = _16398 ^ _16400;
  wire _16402 = _16396 ^ _16401;
  wire _16403 = uncoded_block[1212] ^ uncoded_block[1215];
  wire _16404 = _16403 ^ _2220;
  wire _16405 = _4502 ^ _609;
  wire _16406 = _16404 ^ _16405;
  wire _16407 = _12819 ^ _14919;
  wire _16408 = uncoded_block[1241] ^ uncoded_block[1244];
  wire _16409 = _2989 ^ _16408;
  wire _16410 = _16407 ^ _16409;
  wire _16411 = _16406 ^ _16410;
  wire _16412 = _16402 ^ _16411;
  wire _16413 = _3780 ^ _1455;
  wire _16414 = _5900 ^ _16413;
  wire _16415 = _5234 ^ _8391;
  wire _16416 = _7179 ^ _9538;
  wire _16417 = _16415 ^ _16416;
  wire _16418 = _16414 ^ _16417;
  wire _16419 = uncoded_block[1274] ^ uncoded_block[1275];
  wire _16420 = _16419 ^ _631;
  wire _16421 = _6560 ^ _639;
  wire _16422 = _16420 ^ _16421;
  wire _16423 = _4529 ^ _1469;
  wire _16424 = uncoded_block[1301] ^ uncoded_block[1302];
  wire _16425 = _6563 ^ _16424;
  wire _16426 = _16423 ^ _16425;
  wire _16427 = _16422 ^ _16426;
  wire _16428 = _16418 ^ _16427;
  wire _16429 = _16412 ^ _16428;
  wire _16430 = _16392 ^ _16429;
  wire _16431 = uncoded_block[1303] ^ uncoded_block[1306];
  wire _16432 = _16431 ^ _14430;
  wire _16433 = _14432 ^ _4540;
  wire _16434 = _16432 ^ _16433;
  wire _16435 = uncoded_block[1327] ^ uncoded_block[1331];
  wire _16436 = _3032 ^ _16435;
  wire _16437 = uncoded_block[1335] ^ uncoded_block[1338];
  wire _16438 = _3820 ^ _16437;
  wire _16439 = _16436 ^ _16438;
  wire _16440 = _16434 ^ _16439;
  wire _16441 = _669 ^ _1502;
  wire _16442 = _13928 ^ _16441;
  wire _16443 = _5940 ^ _6588;
  wire _16444 = uncoded_block[1361] ^ uncoded_block[1364];
  wire _16445 = _16444 ^ _3052;
  wire _16446 = _16443 ^ _16445;
  wire _16447 = _16442 ^ _16446;
  wire _16448 = _16440 ^ _16447;
  wire _16449 = uncoded_block[1371] ^ uncoded_block[1374];
  wire _16450 = _16449 ^ _12305;
  wire _16451 = uncoded_block[1380] ^ uncoded_block[1382];
  wire _16452 = _2290 ^ _16451;
  wire _16453 = _16450 ^ _16452;
  wire _16454 = _3061 ^ _7222;
  wire _16455 = _691 ^ _5952;
  wire _16456 = _16454 ^ _16455;
  wire _16457 = _16453 ^ _16456;
  wire _16458 = uncoded_block[1399] ^ uncoded_block[1402];
  wire _16459 = uncoded_block[1403] ^ uncoded_block[1407];
  wire _16460 = _16458 ^ _16459;
  wire _16461 = _7226 ^ _16460;
  wire _16462 = _5957 ^ _12877;
  wire _16463 = uncoded_block[1420] ^ uncoded_block[1421];
  wire _16464 = _12322 ^ _16463;
  wire _16465 = _16462 ^ _16464;
  wire _16466 = _16461 ^ _16465;
  wire _16467 = _16457 ^ _16466;
  wire _16468 = _16448 ^ _16467;
  wire _16469 = uncoded_block[1422] ^ uncoded_block[1427];
  wire _16470 = _16469 ^ _9590;
  wire _16471 = _15982 ^ _2321;
  wire _16472 = _16470 ^ _16471;
  wire _16473 = uncoded_block[1445] ^ uncoded_block[1449];
  wire _16474 = uncoded_block[1452] ^ uncoded_block[1455];
  wire _16475 = _16473 ^ _16474;
  wire _16476 = _3088 ^ _7243;
  wire _16477 = _16475 ^ _16476;
  wire _16478 = _16472 ^ _16477;
  wire _16479 = uncoded_block[1473] ^ uncoded_block[1478];
  wire _16480 = _7247 ^ _16479;
  wire _16481 = _11807 ^ _2349;
  wire _16482 = _16480 ^ _16481;
  wire _16483 = _4610 ^ _13967;
  wire _16484 = _2352 ^ _15515;
  wire _16485 = _16483 ^ _16484;
  wire _16486 = _16482 ^ _16485;
  wire _16487 = _16478 ^ _16486;
  wire _16488 = uncoded_block[1510] ^ uncoded_block[1512];
  wire _16489 = _3112 ^ _16488;
  wire _16490 = _16489 ^ _5338;
  wire _16491 = _754 ^ _9059;
  wire _16492 = _8473 ^ _4623;
  wire _16493 = _16491 ^ _16492;
  wire _16494 = _16490 ^ _16493;
  wire _16495 = _2360 ^ _9631;
  wire _16496 = uncoded_block[1533] ^ uncoded_block[1537];
  wire _16497 = _16496 ^ _6651;
  wire _16498 = _16495 ^ _16497;
  wire _16499 = uncoded_block[1543] ^ uncoded_block[1546];
  wire _16500 = _1589 ^ _16499;
  wire _16501 = uncoded_block[1550] ^ uncoded_block[1553];
  wire _16502 = _7275 ^ _16501;
  wire _16503 = _16500 ^ _16502;
  wire _16504 = _16498 ^ _16503;
  wire _16505 = _16494 ^ _16504;
  wire _16506 = _16487 ^ _16505;
  wire _16507 = _16468 ^ _16506;
  wire _16508 = _16430 ^ _16507;
  wire _16509 = _3131 ^ _6016;
  wire _16510 = uncoded_block[1567] ^ uncoded_block[1570];
  wire _16511 = _3139 ^ _16510;
  wire _16512 = _16509 ^ _16511;
  wire _16513 = uncoded_block[1578] ^ uncoded_block[1582];
  wire _16514 = _1608 ^ _16513;
  wire _16515 = uncoded_block[1586] ^ uncoded_block[1590];
  wire _16516 = _15537 ^ _16515;
  wire _16517 = _16514 ^ _16516;
  wire _16518 = _16512 ^ _16517;
  wire _16519 = _12935 ^ _11847;
  wire _16520 = uncoded_block[1603] ^ uncoded_block[1608];
  wire _16521 = _16520 ^ _7906;
  wire _16522 = _16519 ^ _16521;
  wire _16523 = _5382 ^ _804;
  wire _16524 = _9095 ^ _7300;
  wire _16525 = _16523 ^ _16524;
  wire _16526 = _16522 ^ _16525;
  wire _16527 = _16518 ^ _16526;
  wire _16528 = _807 ^ _2404;
  wire _16529 = uncoded_block[1632] ^ uncoded_block[1635];
  wire _16530 = _16529 ^ _10754;
  wire _16531 = _16528 ^ _16530;
  wire _16532 = _6689 ^ _815;
  wire _16533 = _7312 ^ _9661;
  wire _16534 = _16532 ^ _16533;
  wire _16535 = _16531 ^ _16534;
  wire _16536 = _15559 ^ _5398;
  wire _16537 = uncoded_block[1662] ^ uncoded_block[1665];
  wire _16538 = _16537 ^ _2422;
  wire _16539 = _16536 ^ _16538;
  wire _16540 = _6700 ^ _5401;
  wire _16541 = uncoded_block[1679] ^ uncoded_block[1682];
  wire _16542 = _16541 ^ _4693;
  wire _16543 = _16540 ^ _16542;
  wire _16544 = _16539 ^ _16543;
  wire _16545 = _16535 ^ _16544;
  wire _16546 = _16527 ^ _16545;
  wire _16547 = _14543 ^ _13519;
  wire _16548 = _11325 ^ _844;
  wire _16549 = _16547 ^ _16548;
  wire _16550 = _6068 ^ _4700;
  wire _16551 = uncoded_block[1704] ^ uncoded_block[1708];
  wire _16552 = _16551 ^ _10778;
  wire _16553 = _16550 ^ _16552;
  wire _16554 = _16549 ^ _16553;
  wire _16555 = _14553 ^ uncoded_block[1720];
  wire _16556 = _16554 ^ _16555;
  wire _16557 = _16546 ^ _16556;
  wire _16558 = _16508 ^ _16557;
  wire _16559 = _16358 ^ _16558;
  wire _16560 = uncoded_block[0] ^ uncoded_block[4];
  wire _16561 = _16560 ^ _4712;
  wire _16562 = _6724 ^ _4;
  wire _16563 = _16561 ^ _16562;
  wire _16564 = uncoded_block[13] ^ uncoded_block[16];
  wire _16565 = _7 ^ _16564;
  wire _16566 = _16565 ^ _9695;
  wire _16567 = _16563 ^ _16566;
  wire _16568 = _11344 ^ _875;
  wire _16569 = _6095 ^ _18;
  wire _16570 = _16568 ^ _16569;
  wire _16571 = _19 ^ _10234;
  wire _16572 = uncoded_block[55] ^ uncoded_block[57];
  wire _16573 = _6101 ^ _16572;
  wire _16574 = _16571 ^ _16573;
  wire _16575 = _16570 ^ _16574;
  wire _16576 = _16567 ^ _16575;
  wire _16577 = uncoded_block[64] ^ uncoded_block[69];
  wire _16578 = _2472 ^ _16577;
  wire _16579 = uncoded_block[72] ^ uncoded_block[80];
  wire _16580 = uncoded_block[82] ^ uncoded_block[86];
  wire _16581 = _16579 ^ _16580;
  wire _16582 = _16578 ^ _16581;
  wire _16583 = _6755 ^ _903;
  wire _16584 = uncoded_block[93] ^ uncoded_block[97];
  wire _16585 = _16584 ^ _11909;
  wire _16586 = _16583 ^ _16585;
  wire _16587 = _16582 ^ _16586;
  wire _16588 = _3250 ^ _1722;
  wire _16589 = uncoded_block[113] ^ uncoded_block[116];
  wire _16590 = _15103 ^ _16589;
  wire _16591 = _16588 ^ _16590;
  wire _16592 = uncoded_block[117] ^ uncoded_block[120];
  wire _16593 = _16592 ^ _10256;
  wire _16594 = _1730 ^ _4754;
  wire _16595 = _16593 ^ _16594;
  wire _16596 = _16591 ^ _16595;
  wire _16597 = _16587 ^ _16596;
  wire _16598 = _16576 ^ _16597;
  wire _16599 = uncoded_block[132] ^ uncoded_block[140];
  wire _16600 = uncoded_block[142] ^ uncoded_block[144];
  wire _16601 = _16599 ^ _16600;
  wire _16602 = _6780 ^ _5470;
  wire _16603 = _16601 ^ _16602;
  wire _16604 = uncoded_block[165] ^ uncoded_block[168];
  wire _16605 = _15118 ^ _16604;
  wire _16606 = _15123 ^ _11933;
  wire _16607 = _16605 ^ _16606;
  wire _16608 = _16603 ^ _16607;
  wire _16609 = _5479 ^ _10275;
  wire _16610 = _947 ^ _1763;
  wire _16611 = _16609 ^ _16610;
  wire _16612 = _15135 ^ _10278;
  wire _16613 = _14101 ^ _955;
  wire _16614 = _16612 ^ _16613;
  wire _16615 = _16611 ^ _16614;
  wire _16616 = _16608 ^ _16615;
  wire _16617 = _2540 ^ _4787;
  wire _16618 = uncoded_block[220] ^ uncoded_block[225];
  wire _16619 = _16618 ^ _109;
  wire _16620 = _16617 ^ _16619;
  wire _16621 = _1774 ^ _967;
  wire _16622 = uncoded_block[239] ^ uncoded_block[242];
  wire _16623 = _968 ^ _16622;
  wire _16624 = _16621 ^ _16623;
  wire _16625 = _16620 ^ _16624;
  wire _16626 = uncoded_block[246] ^ uncoded_block[248];
  wire _16627 = _4085 ^ _16626;
  wire _16628 = _14116 ^ _117;
  wire _16629 = _16627 ^ _16628;
  wire _16630 = _13055 ^ _7438;
  wire _16631 = _16630 ^ _4805;
  wire _16632 = _16629 ^ _16631;
  wire _16633 = _16625 ^ _16632;
  wire _16634 = _16616 ^ _16633;
  wire _16635 = _16598 ^ _16634;
  wire _16636 = uncoded_block[269] ^ uncoded_block[271];
  wire _16637 = _11421 ^ _16636;
  wire _16638 = _2568 ^ _5515;
  wire _16639 = _16637 ^ _16638;
  wire _16640 = _11424 ^ _1803;
  wire _16641 = _5522 ^ _6838;
  wire _16642 = _16640 ^ _16641;
  wire _16643 = _16639 ^ _16642;
  wire _16644 = _4820 ^ _10312;
  wire _16645 = uncoded_block[300] ^ uncoded_block[304];
  wire _16646 = _16645 ^ _4114;
  wire _16647 = _16644 ^ _16646;
  wire _16648 = uncoded_block[311] ^ uncoded_block[314];
  wire _16649 = _3337 ^ _16648;
  wire _16650 = _6208 ^ _8642;
  wire _16651 = _16649 ^ _16650;
  wire _16652 = _16647 ^ _16651;
  wire _16653 = _16643 ^ _16652;
  wire _16654 = _1819 ^ _2587;
  wire _16655 = _16654 ^ _6858;
  wire _16656 = _1021 ^ _4844;
  wire _16657 = _3359 ^ _4132;
  wire _16658 = _16656 ^ _16657;
  wire _16659 = _16655 ^ _16658;
  wire _16660 = _2606 ^ _5548;
  wire _16661 = _4136 ^ _16660;
  wire _16662 = uncoded_block[367] ^ uncoded_block[369];
  wire _16663 = _7470 ^ _16662;
  wire _16664 = uncoded_block[370] ^ uncoded_block[375];
  wire _16665 = _16664 ^ _4854;
  wire _16666 = _16663 ^ _16665;
  wire _16667 = _16661 ^ _16666;
  wire _16668 = _16659 ^ _16667;
  wire _16669 = _16653 ^ _16668;
  wire _16670 = _11999 ^ _176;
  wire _16671 = uncoded_block[391] ^ uncoded_block[395];
  wire _16672 = _16671 ^ _5559;
  wire _16673 = _16670 ^ _16672;
  wire _16674 = _15697 ^ _184;
  wire _16675 = _10344 ^ _14682;
  wire _16676 = _16674 ^ _16675;
  wire _16677 = _16673 ^ _16676;
  wire _16678 = _11477 ^ _12551;
  wire _16679 = _9816 ^ _10352;
  wire _16680 = _16678 ^ _16679;
  wire _16681 = _2641 ^ _205;
  wire _16682 = _10356 ^ _3411;
  wire _16683 = _16681 ^ _16682;
  wire _16684 = _16680 ^ _16683;
  wire _16685 = _16677 ^ _16684;
  wire _16686 = _12562 ^ _5584;
  wire _16687 = uncoded_block[460] ^ uncoded_block[464];
  wire _16688 = _3415 ^ _16687;
  wire _16689 = _16686 ^ _16688;
  wire _16690 = uncoded_block[465] ^ uncoded_block[468];
  wire _16691 = _16690 ^ _4186;
  wire _16692 = uncoded_block[471] ^ uncoded_block[475];
  wire _16693 = uncoded_block[479] ^ uncoded_block[481];
  wire _16694 = _16692 ^ _16693;
  wire _16695 = _16691 ^ _16694;
  wire _16696 = _16689 ^ _16695;
  wire _16697 = _4897 ^ _4194;
  wire _16698 = _8117 ^ _13139;
  wire _16699 = _16697 ^ _16698;
  wire _16700 = uncoded_block[499] ^ uncoded_block[508];
  wire _16701 = _16700 ^ _7531;
  wire _16702 = _13676 ^ _8706;
  wire _16703 = _16701 ^ _16702;
  wire _16704 = _16699 ^ _16703;
  wire _16705 = _16696 ^ _16704;
  wire _16706 = _16685 ^ _16705;
  wire _16707 = _16669 ^ _16706;
  wire _16708 = _16635 ^ _16707;
  wire _16709 = uncoded_block[523] ^ uncoded_block[525];
  wire _16710 = _1107 ^ _16709;
  wire _16711 = uncoded_block[527] ^ uncoded_block[530];
  wire _16712 = _16711 ^ _6931;
  wire _16713 = _16710 ^ _16712;
  wire _16714 = _1905 ^ _14721;
  wire _16715 = uncoded_block[544] ^ uncoded_block[546];
  wire _16716 = _16715 ^ _12592;
  wire _16717 = _16714 ^ _16716;
  wire _16718 = _16713 ^ _16717;
  wire _16719 = _1913 ^ _1915;
  wire _16720 = _12051 ^ _1924;
  wire _16721 = _16719 ^ _16720;
  wire _16722 = _1126 ^ _6309;
  wire _16723 = _4941 ^ _1132;
  wire _16724 = _16722 ^ _16723;
  wire _16725 = _16721 ^ _16724;
  wire _16726 = _16718 ^ _16725;
  wire _16727 = uncoded_block[578] ^ uncoded_block[582];
  wire _16728 = _16727 ^ _1933;
  wire _16729 = _9864 ^ _2700;
  wire _16730 = _16728 ^ _16729;
  wire _16731 = _6316 ^ _10408;
  wire _16732 = _16731 ^ _10410;
  wire _16733 = _16730 ^ _16732;
  wire _16734 = uncoded_block[609] ^ uncoded_block[611];
  wire _16735 = _277 ^ _16734;
  wire _16736 = _6325 ^ _4243;
  wire _16737 = _16735 ^ _16736;
  wire _16738 = uncoded_block[620] ^ uncoded_block[623];
  wire _16739 = _16738 ^ _8161;
  wire _16740 = uncoded_block[635] ^ uncoded_block[640];
  wire _16741 = _16740 ^ _294;
  wire _16742 = _16739 ^ _16741;
  wire _16743 = _16737 ^ _16742;
  wire _16744 = _16733 ^ _16743;
  wire _16745 = _16726 ^ _16744;
  wire _16746 = _6973 ^ _302;
  wire _16747 = uncoded_block[656] ^ uncoded_block[659];
  wire _16748 = _304 ^ _16747;
  wire _16749 = _16746 ^ _16748;
  wire _16750 = _2739 ^ _12630;
  wire _16751 = uncoded_block[666] ^ uncoded_block[670];
  wire _16752 = uncoded_block[671] ^ uncoded_block[673];
  wire _16753 = _16751 ^ _16752;
  wire _16754 = _16750 ^ _16753;
  wire _16755 = _16749 ^ _16754;
  wire _16756 = _13731 ^ _6353;
  wire _16757 = uncoded_block[689] ^ uncoded_block[695];
  wire _16758 = _6983 ^ _16757;
  wire _16759 = _16756 ^ _16758;
  wire _16760 = _3529 ^ _14249;
  wire _16761 = uncoded_block[708] ^ uncoded_block[710];
  wire _16762 = _7595 ^ _16761;
  wire _16763 = _16760 ^ _16762;
  wire _16764 = _16759 ^ _16763;
  wire _16765 = _16755 ^ _16764;
  wire _16766 = _2762 ^ _4999;
  wire _16767 = _5002 ^ _341;
  wire _16768 = _16766 ^ _16767;
  wire _16769 = uncoded_block[725] ^ uncoded_block[730];
  wire _16770 = _6374 ^ _16769;
  wire _16771 = _3547 ^ _2770;
  wire _16772 = _16770 ^ _16771;
  wire _16773 = _16768 ^ _16772;
  wire _16774 = _5702 ^ _3554;
  wire _16775 = uncoded_block[749] ^ uncoded_block[752];
  wire _16776 = uncoded_block[753] ^ uncoded_block[758];
  wire _16777 = _16775 ^ _16776;
  wire _16778 = _16774 ^ _16777;
  wire _16779 = _2006 ^ _4301;
  wire _16780 = _6382 ^ _2794;
  wire _16781 = _16779 ^ _16780;
  wire _16782 = _16778 ^ _16781;
  wire _16783 = _16773 ^ _16782;
  wire _16784 = _16765 ^ _16783;
  wire _16785 = _16745 ^ _16784;
  wire _16786 = uncoded_block[783] ^ uncoded_block[786];
  wire _16787 = _16786 ^ _8790;
  wire _16788 = _2799 ^ _382;
  wire _16789 = _16787 ^ _16788;
  wire _16790 = uncoded_block[799] ^ uncoded_block[803];
  wire _16791 = uncoded_block[806] ^ uncoded_block[807];
  wire _16792 = _16790 ^ _16791;
  wire _16793 = uncoded_block[808] ^ uncoded_block[810];
  wire _16794 = _16793 ^ _10483;
  wire _16795 = _16792 ^ _16794;
  wire _16796 = _16789 ^ _16795;
  wire _16797 = uncoded_block[817] ^ uncoded_block[823];
  wire _16798 = _4324 ^ _16797;
  wire _16799 = _1246 ^ _6401;
  wire _16800 = _16798 ^ _16799;
  wire _16801 = uncoded_block[834] ^ uncoded_block[835];
  wire _16802 = _7039 ^ _16801;
  wire _16803 = _11043 ^ _7640;
  wire _16804 = _16802 ^ _16803;
  wire _16805 = _16800 ^ _16804;
  wire _16806 = _16796 ^ _16805;
  wire _16807 = _405 ^ _7643;
  wire _16808 = uncoded_block[855] ^ uncoded_block[862];
  wire _16809 = _8237 ^ _16808;
  wire _16810 = _16807 ^ _16809;
  wire _16811 = uncoded_block[867] ^ uncoded_block[870];
  wire _16812 = _14302 ^ _16811;
  wire _16813 = _16812 ^ _418;
  wire _16814 = _16810 ^ _16813;
  wire _16815 = uncoded_block[877] ^ uncoded_block[878];
  wire _16816 = _16815 ^ _5079;
  wire _16817 = _2838 ^ _11059;
  wire _16818 = _16816 ^ _16817;
  wire _16819 = uncoded_block[890] ^ uncoded_block[892];
  wire _16820 = _16819 ^ _2843;
  wire _16821 = uncoded_block[905] ^ uncoded_block[908];
  wire _16822 = _2844 ^ _16821;
  wire _16823 = _16820 ^ _16822;
  wire _16824 = _16818 ^ _16823;
  wire _16825 = _16814 ^ _16824;
  wire _16826 = _16806 ^ _16825;
  wire _16827 = uncoded_block[926] ^ uncoded_block[927];
  wire _16828 = _439 ^ _16827;
  wire _16829 = _1296 ^ _5096;
  wire _16830 = _16828 ^ _16829;
  wire _16831 = _15352 ^ _16830;
  wire _16832 = uncoded_block[939] ^ uncoded_block[942];
  wire _16833 = _2079 ^ _16832;
  wire _16834 = _2865 ^ _2086;
  wire _16835 = _16833 ^ _16834;
  wire _16836 = _14329 ^ _11642;
  wire _16837 = _13267 ^ _16836;
  wire _16838 = _16835 ^ _16837;
  wire _16839 = _16831 ^ _16838;
  wire _16840 = _2871 ^ _12179;
  wire _16841 = uncoded_block[975] ^ uncoded_block[978];
  wire _16842 = _11087 ^ _16841;
  wire _16843 = _16840 ^ _16842;
  wire _16844 = uncoded_block[982] ^ uncoded_block[987];
  wire _16845 = _5790 ^ _16844;
  wire _16846 = _12737 ^ _2883;
  wire _16847 = _16845 ^ _16846;
  wire _16848 = _16843 ^ _16847;
  wire _16849 = _2107 ^ _2112;
  wire _16850 = _6459 ^ _5129;
  wire _16851 = _16849 ^ _16850;
  wire _16852 = uncoded_block[1010] ^ uncoded_block[1017];
  wire _16853 = uncoded_block[1018] ^ uncoded_block[1020];
  wire _16854 = _16852 ^ _16853;
  wire _16855 = _5137 ^ _8874;
  wire _16856 = _16854 ^ _16855;
  wire _16857 = _16851 ^ _16856;
  wire _16858 = _16848 ^ _16857;
  wire _16859 = _16839 ^ _16858;
  wire _16860 = _16826 ^ _16859;
  wire _16861 = _16785 ^ _16860;
  wire _16862 = _16708 ^ _16861;
  wire _16863 = _13289 ^ _8881;
  wire _16864 = uncoded_block[1042] ^ uncoded_block[1045];
  wire _16865 = _16864 ^ _2914;
  wire _16866 = _519 ^ _3684;
  wire _16867 = _16865 ^ _16866;
  wire _16868 = _16863 ^ _16867;
  wire _16869 = uncoded_block[1064] ^ uncoded_block[1069];
  wire _16870 = _16869 ^ _2143;
  wire _16871 = _5831 ^ _2924;
  wire _16872 = _16870 ^ _16871;
  wire _16873 = _530 ^ _1371;
  wire _16874 = _1373 ^ _2930;
  wire _16875 = _16873 ^ _16874;
  wire _16876 = _16872 ^ _16875;
  wire _16877 = _16868 ^ _16876;
  wire _16878 = uncoded_block[1095] ^ uncoded_block[1098];
  wire _16879 = _16878 ^ _5169;
  wire _16880 = uncoded_block[1101] ^ uncoded_block[1106];
  wire _16881 = uncoded_block[1108] ^ uncoded_block[1113];
  wire _16882 = _16880 ^ _16881;
  wire _16883 = _16879 ^ _16882;
  wire _16884 = _3713 ^ _1388;
  wire _16885 = _2941 ^ _558;
  wire _16886 = _16884 ^ _16885;
  wire _16887 = _16883 ^ _16886;
  wire _16888 = _9494 ^ _5181;
  wire _16889 = _3721 ^ _574;
  wire _16890 = _16888 ^ _16889;
  wire _16891 = _7143 ^ _3728;
  wire _16892 = _578 ^ _2958;
  wire _16893 = _16891 ^ _16892;
  wire _16894 = _16890 ^ _16893;
  wire _16895 = _16887 ^ _16894;
  wire _16896 = _16877 ^ _16895;
  wire _16897 = _2964 ^ _7151;
  wire _16898 = uncoded_block[1175] ^ uncoded_block[1179];
  wire _16899 = _3739 ^ _16898;
  wire _16900 = _16897 ^ _16899;
  wire _16901 = uncoded_block[1183] ^ uncoded_block[1185];
  wire _16902 = _2195 ^ _16901;
  wire _16903 = _5201 ^ _4488;
  wire _16904 = _16902 ^ _16903;
  wire _16905 = _16900 ^ _16904;
  wire _16906 = _7758 ^ _2974;
  wire _16907 = uncoded_block[1207] ^ uncoded_block[1214];
  wire _16908 = _2210 ^ _16907;
  wire _16909 = _16906 ^ _16908;
  wire _16910 = _2219 ^ _606;
  wire _16911 = _4502 ^ _9522;
  wire _16912 = _16910 ^ _16911;
  wire _16913 = _16909 ^ _16912;
  wire _16914 = _16905 ^ _16913;
  wire _16915 = uncoded_block[1237] ^ uncoded_block[1240];
  wire _16916 = _3769 ^ _16915;
  wire _16917 = _3779 ^ _2235;
  wire _16918 = _16916 ^ _16917;
  wire _16919 = uncoded_block[1262] ^ uncoded_block[1266];
  wire _16920 = _16919 ^ _7179;
  wire _16921 = _6549 ^ _16920;
  wire _16922 = _16918 ^ _16921;
  wire _16923 = _628 ^ _630;
  wire _16924 = uncoded_block[1282] ^ uncoded_block[1286];
  wire _16925 = _6556 ^ _16924;
  wire _16926 = _16923 ^ _16925;
  wire _16927 = _641 ^ _1469;
  wire _16928 = _4531 ^ _6564;
  wire _16929 = _16927 ^ _16928;
  wire _16930 = _16926 ^ _16929;
  wire _16931 = _16922 ^ _16930;
  wire _16932 = _16914 ^ _16931;
  wire _16933 = _16896 ^ _16932;
  wire _16934 = _14430 ^ _3811;
  wire _16935 = _650 ^ _16934;
  wire _16936 = uncoded_block[1318] ^ uncoded_block[1332];
  wire _16937 = _16936 ^ _3034;
  wire _16938 = uncoded_block[1339] ^ uncoded_block[1343];
  wire _16939 = _16938 ^ _664;
  wire _16940 = _16937 ^ _16939;
  wire _16941 = _16935 ^ _16940;
  wire _16942 = uncoded_block[1354] ^ uncoded_block[1356];
  wire _16943 = _16942 ^ _5940;
  wire _16944 = _14955 ^ _16943;
  wire _16945 = _3047 ^ _11226;
  wire _16946 = _678 ^ _16945;
  wire _16947 = _16944 ^ _16946;
  wire _16948 = _16941 ^ _16947;
  wire _16949 = _10669 ^ _5285;
  wire _16950 = _3834 ^ _3061;
  wire _16951 = _16949 ^ _16950;
  wire _16952 = uncoded_block[1388] ^ uncoded_block[1392];
  wire _16953 = _16952 ^ _4569;
  wire _16954 = uncoded_block[1405] ^ uncoded_block[1407];
  wire _16955 = _16458 ^ _16954;
  wire _16956 = _16953 ^ _16955;
  wire _16957 = _16951 ^ _16956;
  wire _16958 = _8436 ^ _702;
  wire _16959 = _5964 ^ _3074;
  wire _16960 = _16958 ^ _16959;
  wire _16961 = _2308 ^ _9590;
  wire _16962 = uncoded_block[1432] ^ uncoded_block[1435];
  wire _16963 = _16962 ^ _3857;
  wire _16964 = _16961 ^ _16963;
  wire _16965 = _16960 ^ _16964;
  wire _16966 = _16957 ^ _16965;
  wire _16967 = _16948 ^ _16966;
  wire _16968 = _3083 ^ _6613;
  wire _16969 = uncoded_block[1444] ^ uncoded_block[1449];
  wire _16970 = uncoded_block[1450] ^ uncoded_block[1453];
  wire _16971 = _16969 ^ _16970;
  wire _16972 = _16968 ^ _16971;
  wire _16973 = _6622 ^ _4596;
  wire _16974 = _3871 ^ _1550;
  wire _16975 = _16973 ^ _16974;
  wire _16976 = _16972 ^ _16975;
  wire _16977 = uncoded_block[1470] ^ uncoded_block[1473];
  wire _16978 = _16977 ^ _733;
  wire _16979 = _13963 ^ _739;
  wire _16980 = _16978 ^ _16979;
  wire _16981 = uncoded_block[1488] ^ uncoded_block[1490];
  wire _16982 = _16981 ^ _9614;
  wire _16983 = _12898 ^ _6634;
  wire _16984 = _16982 ^ _16983;
  wire _16985 = _16980 ^ _16984;
  wire _16986 = _16976 ^ _16985;
  wire _16987 = _4616 ^ _5334;
  wire _16988 = uncoded_block[1521] ^ uncoded_block[1523];
  wire _16989 = _15004 ^ _16988;
  wire _16990 = _16987 ^ _16989;
  wire _16991 = _8473 ^ _1582;
  wire _16992 = _16008 ^ _6651;
  wire _16993 = _16991 ^ _16992;
  wire _16994 = _16990 ^ _16993;
  wire _16995 = uncoded_block[1545] ^ uncoded_block[1548];
  wire _16996 = _7883 ^ _16995;
  wire _16997 = _6657 ^ _9070;
  wire _16998 = _16996 ^ _16997;
  wire _16999 = _1596 ^ _10160;
  wire _17000 = _1605 ^ _9072;
  wire _17001 = _16999 ^ _17000;
  wire _17002 = _16998 ^ _17001;
  wire _17003 = _16994 ^ _17002;
  wire _17004 = _16986 ^ _17003;
  wire _17005 = _16967 ^ _17004;
  wire _17006 = _16933 ^ _17005;
  wire _17007 = uncoded_block[1572] ^ uncoded_block[1574];
  wire _17008 = _17007 ^ _4648;
  wire _17009 = uncoded_block[1583] ^ uncoded_block[1586];
  wire _17010 = _4651 ^ _17009;
  wire _17011 = _17008 ^ _17010;
  wire _17012 = _5368 ^ _12934;
  wire _17013 = uncoded_block[1594] ^ uncoded_block[1598];
  wire _17014 = _791 ^ _17013;
  wire _17015 = _17012 ^ _17014;
  wire _17016 = _17011 ^ _17015;
  wire _17017 = _798 ^ _1625;
  wire _17018 = _3154 ^ _801;
  wire _17019 = _17017 ^ _17018;
  wire _17020 = uncoded_block[1614] ^ uncoded_block[1616];
  wire _17021 = _17020 ^ _7911;
  wire _17022 = uncoded_block[1626] ^ uncoded_block[1634];
  wire _17023 = _3941 ^ _17022;
  wire _17024 = _17021 ^ _17023;
  wire _17025 = _17019 ^ _17024;
  wire _17026 = _17016 ^ _17025;
  wire _17027 = uncoded_block[1637] ^ uncoded_block[1644];
  wire _17028 = _17027 ^ _7312;
  wire _17029 = _10757 ^ _4677;
  wire _17030 = _17028 ^ _17029;
  wire _17031 = _14011 ^ _3174;
  wire _17032 = uncoded_block[1663] ^ uncoded_block[1666];
  wire _17033 = _10196 ^ _17032;
  wire _17034 = _17031 ^ _17033;
  wire _17035 = _17030 ^ _17034;
  wire _17036 = _16052 ^ _8521;
  wire _17037 = _7323 ^ _3183;
  wire _17038 = _17036 ^ _17037;
  wire _17039 = _11321 ^ _10766;
  wire _17040 = uncoded_block[1682] ^ uncoded_block[1683];
  wire _17041 = uncoded_block[1685] ^ uncoded_block[1690];
  wire _17042 = _17040 ^ _17041;
  wire _17043 = _17039 ^ _17042;
  wire _17044 = _17038 ^ _17043;
  wire _17045 = _17035 ^ _17044;
  wire _17046 = _17026 ^ _17045;
  wire _17047 = _4700 ^ _847;
  wire _17048 = _14026 ^ _17047;
  wire _17049 = _7944 ^ _2443;
  wire _17050 = _13524 ^ _17049;
  wire _17051 = _17048 ^ _17050;
  wire _17052 = _17051 ^ uncoded_block[1720];
  wire _17053 = _17046 ^ _17052;
  wire _17054 = _17006 ^ _17053;
  wire _17055 = _16862 ^ _17054;
  wire _17056 = _6080 ^ _6082;
  wire _17057 = _3211 ^ _17056;
  wire _17058 = uncoded_block[10] ^ uncoded_block[12];
  wire _17059 = _17058 ^ _871;
  wire _17060 = uncoded_block[19] ^ uncoded_block[24];
  wire _17061 = _17060 ^ _13539;
  wire _17062 = _17059 ^ _17061;
  wire _17063 = _17057 ^ _17062;
  wire _17064 = _15589 ^ _10797;
  wire _17065 = uncoded_block[42] ^ uncoded_block[45];
  wire _17066 = _17065 ^ _6099;
  wire _17067 = uncoded_block[49] ^ uncoded_block[52];
  wire _17068 = _17067 ^ _5436;
  wire _17069 = _17066 ^ _17068;
  wire _17070 = _17064 ^ _17069;
  wire _17071 = _17063 ^ _17070;
  wire _17072 = _1703 ^ _26;
  wire _17073 = uncoded_block[68] ^ uncoded_block[76];
  wire _17074 = _32 ^ _17073;
  wire _17075 = _17072 ^ _17074;
  wire _17076 = _901 ^ _6749;
  wire _17077 = uncoded_block[84] ^ uncoded_block[86];
  wire _17078 = _6750 ^ _17077;
  wire _17079 = _17076 ^ _17078;
  wire _17080 = _17075 ^ _17079;
  wire _17081 = _15603 ^ _14591;
  wire _17082 = _17081 ^ _14069;
  wire _17083 = _15097 ^ _15101;
  wire _17084 = _6120 ^ _1722;
  wire _17085 = _17083 ^ _17084;
  wire _17086 = _17082 ^ _17085;
  wire _17087 = _17080 ^ _17086;
  wire _17088 = _17071 ^ _17087;
  wire _17089 = _4034 ^ _16589;
  wire _17090 = _6128 ^ _56;
  wire _17091 = _17089 ^ _17090;
  wire _17092 = _2502 ^ _1733;
  wire _17093 = _926 ^ _64;
  wire _17094 = _17092 ^ _17093;
  wire _17095 = _17091 ^ _17094;
  wire _17096 = _5461 ^ _6138;
  wire _17097 = uncoded_block[145] ^ uncoded_block[147];
  wire _17098 = _17097 ^ _8000;
  wire _17099 = _17096 ^ _17098;
  wire _17100 = uncoded_block[154] ^ uncoded_block[159];
  wire _17101 = _3269 ^ _17100;
  wire _17102 = _17101 ^ _14087;
  wire _17103 = _17099 ^ _17102;
  wire _17104 = _17095 ^ _17103;
  wire _17105 = uncoded_block[177] ^ uncoded_block[181];
  wire _17106 = uncoded_block[184] ^ uncoded_block[186];
  wire _17107 = _17105 ^ _17106;
  wire _17108 = _7402 ^ _17107;
  wire _17109 = _6798 ^ _89;
  wire _17110 = _11397 ^ _17109;
  wire _17111 = _17108 ^ _17110;
  wire _17112 = uncoded_block[198] ^ uncoded_block[200];
  wire _17113 = _17112 ^ _14622;
  wire _17114 = _8021 ^ _98;
  wire _17115 = _17113 ^ _17114;
  wire _17116 = uncoded_block[215] ^ uncoded_block[218];
  wire _17117 = _959 ^ _17116;
  wire _17118 = uncoded_block[225] ^ uncoded_block[228];
  wire _17119 = _4076 ^ _17118;
  wire _17120 = _17117 ^ _17119;
  wire _17121 = _17115 ^ _17120;
  wire _17122 = _17111 ^ _17121;
  wire _17123 = _17104 ^ _17122;
  wire _17124 = _17088 ^ _17123;
  wire _17125 = _970 ^ _9756;
  wire _17126 = _6823 ^ _17125;
  wire _17127 = uncoded_block[242] ^ uncoded_block[245];
  wire _17128 = _17127 ^ _116;
  wire _17129 = _7434 ^ _11419;
  wire _17130 = _17128 ^ _17129;
  wire _17131 = _17126 ^ _17130;
  wire _17132 = _3311 ^ _14639;
  wire _17133 = _17132 ^ _4097;
  wire _17134 = uncoded_block[269] ^ uncoded_block[273];
  wire _17135 = _7440 ^ _17134;
  wire _17136 = _6833 ^ _10304;
  wire _17137 = _17135 ^ _17136;
  wire _17138 = _17133 ^ _17137;
  wire _17139 = _17131 ^ _17138;
  wire _17140 = _4105 ^ _134;
  wire _17141 = _17140 ^ _13614;
  wire _17142 = uncoded_block[297] ^ uncoded_block[299];
  wire _17143 = _4820 ^ _17142;
  wire _17144 = uncoded_block[301] ^ uncoded_block[303];
  wire _17145 = uncoded_block[305] ^ uncoded_block[310];
  wire _17146 = _17144 ^ _17145;
  wire _17147 = _17143 ^ _17146;
  wire _17148 = _17141 ^ _17147;
  wire _17149 = _16648 ^ _146;
  wire _17150 = _4118 ^ _3346;
  wire _17151 = _17149 ^ _17150;
  wire _17152 = _2583 ^ _11444;
  wire _17153 = _9235 ^ _8063;
  wire _17154 = _17152 ^ _17153;
  wire _17155 = _17151 ^ _17154;
  wire _17156 = _17148 ^ _17155;
  wire _17157 = _17139 ^ _17156;
  wire _17158 = _5536 ^ _11984;
  wire _17159 = _2595 ^ _7465;
  wire _17160 = _17158 ^ _17159;
  wire _17161 = _16657 ^ _8070;
  wire _17162 = _17160 ^ _17161;
  wire _17163 = uncoded_block[366] ^ uncoded_block[367];
  wire _17164 = _12530 ^ _17163;
  wire _17165 = uncoded_block[368] ^ uncoded_block[370];
  wire _17166 = _17165 ^ _10895;
  wire _17167 = _17164 ^ _17166;
  wire _17168 = _10335 ^ _2615;
  wire _17169 = _4152 ^ _3388;
  wire _17170 = _17168 ^ _17169;
  wire _17171 = _17167 ^ _17170;
  wire _17172 = _17162 ^ _17171;
  wire _17173 = _1850 ^ _190;
  wire _17174 = _9266 ^ _5565;
  wire _17175 = _17173 ^ _17174;
  wire _17176 = _194 ^ _2633;
  wire _17177 = uncoded_block[426] ^ uncoded_block[429];
  wire _17178 = _17177 ^ _7495;
  wire _17179 = _17176 ^ _17178;
  wire _17180 = _17175 ^ _17179;
  wire _17181 = uncoded_block[440] ^ uncoded_block[444];
  wire _17182 = _2640 ^ _17181;
  wire _17183 = _10356 ^ _208;
  wire _17184 = _17182 ^ _17183;
  wire _17185 = uncoded_block[454] ^ uncoded_block[457];
  wire _17186 = _2645 ^ _17185;
  wire _17187 = _2653 ^ _1079;
  wire _17188 = _17186 ^ _17187;
  wire _17189 = _17184 ^ _17188;
  wire _17190 = _17180 ^ _17189;
  wire _17191 = _17172 ^ _17190;
  wire _17192 = _17157 ^ _17191;
  wire _17193 = _17124 ^ _17192;
  wire _17194 = _1879 ^ _5590;
  wire _17195 = _7513 ^ _12028;
  wire _17196 = _17194 ^ _17195;
  wire _17197 = _4897 ^ _7515;
  wire _17198 = uncoded_block[489] ^ uncoded_block[492];
  wire _17199 = _17198 ^ _3432;
  wire _17200 = _17197 ^ _17199;
  wire _17201 = _17196 ^ _17200;
  wire _17202 = _6919 ^ _4905;
  wire _17203 = _1887 ^ _7529;
  wire _17204 = _17202 ^ _17203;
  wire _17205 = uncoded_block[515] ^ uncoded_block[518];
  wire _17206 = _17205 ^ _3444;
  wire _17207 = _13149 ^ _17206;
  wire _17208 = _17204 ^ _17207;
  wire _17209 = _17201 ^ _17208;
  wire _17210 = _1108 ^ _14716;
  wire _17211 = _10384 ^ _16215;
  wire _17212 = _17210 ^ _17211;
  wire _17213 = _6932 ^ _7536;
  wire _17214 = _8132 ^ _16715;
  wire _17215 = _17213 ^ _17214;
  wire _17216 = _17212 ^ _17215;
  wire _17217 = _1913 ^ _15740;
  wire _17218 = uncoded_block[559] ^ uncoded_block[565];
  wire _17219 = _17218 ^ _1927;
  wire _17220 = _17217 ^ _17219;
  wire _17221 = uncoded_block[571] ^ uncoded_block[572];
  wire _17222 = _17221 ^ _263;
  wire _17223 = _9325 ^ _1934;
  wire _17224 = _17222 ^ _17223;
  wire _17225 = _17220 ^ _17224;
  wire _17226 = _17216 ^ _17225;
  wire _17227 = _17209 ^ _17226;
  wire _17228 = uncoded_block[594] ^ uncoded_block[598];
  wire _17229 = _9330 ^ _17228;
  wire _17230 = _2707 ^ _1146;
  wire _17231 = _17229 ^ _17230;
  wire _17232 = uncoded_block[611] ^ uncoded_block[612];
  wire _17233 = _278 ^ _17232;
  wire _17234 = _14223 ^ _3495;
  wire _17235 = _17233 ^ _17234;
  wire _17236 = _17231 ^ _17235;
  wire _17237 = _12618 ^ _4964;
  wire _17238 = uncoded_block[627] ^ uncoded_block[629];
  wire _17239 = _17238 ^ _14745;
  wire _17240 = _17237 ^ _17239;
  wire _17241 = _5661 ^ _11543;
  wire _17242 = uncoded_block[643] ^ uncoded_block[646];
  wire _17243 = _2727 ^ _17242;
  wire _17244 = _17241 ^ _17243;
  wire _17245 = _17240 ^ _17244;
  wire _17246 = _17236 ^ _17245;
  wire _17247 = _3507 ^ _16249;
  wire _17248 = uncoded_block[658] ^ uncoded_block[664];
  wire _17249 = _17248 ^ _16751;
  wire _17250 = _17247 ^ _17249;
  wire _17251 = _312 ^ _3519;
  wire _17252 = _8179 ^ _3526;
  wire _17253 = _17251 ^ _17252;
  wire _17254 = _17250 ^ _17253;
  wire _17255 = _3527 ^ _13735;
  wire _17256 = _3529 ^ _6360;
  wire _17257 = _17255 ^ _17256;
  wire _17258 = uncoded_block[700] ^ uncoded_block[702];
  wire _17259 = _17258 ^ _10447;
  wire _17260 = _10448 ^ _337;
  wire _17261 = _17259 ^ _17260;
  wire _17262 = _17257 ^ _17261;
  wire _17263 = _17254 ^ _17262;
  wire _17264 = _17246 ^ _17263;
  wire _17265 = _17227 ^ _17264;
  wire _17266 = uncoded_block[715] ^ uncoded_block[717];
  wire _17267 = _17266 ^ _9369;
  wire _17268 = uncoded_block[723] ^ uncoded_block[730];
  wire _17269 = _17268 ^ _7002;
  wire _17270 = _17267 ^ _17269;
  wire _17271 = _1995 ^ _7005;
  wire _17272 = uncoded_block[741] ^ uncoded_block[745];
  wire _17273 = _17272 ^ _5013;
  wire _17274 = _17271 ^ _17273;
  wire _17275 = _17270 ^ _17274;
  wire _17276 = _2002 ^ _1214;
  wire _17277 = _2778 ^ _15795;
  wire _17278 = _17276 ^ _17277;
  wire _17279 = _5020 ^ _1218;
  wire _17280 = _8787 ^ _9382;
  wire _17281 = _17279 ^ _17280;
  wire _17282 = _17278 ^ _17281;
  wire _17283 = _17275 ^ _17282;
  wire _17284 = uncoded_block[779] ^ uncoded_block[781];
  wire _17285 = uncoded_block[783] ^ uncoded_block[785];
  wire _17286 = _17284 ^ _17285;
  wire _17287 = _17286 ^ _5034;
  wire _17288 = _8791 ^ _8223;
  wire _17289 = _17288 ^ _15815;
  wire _17290 = _17287 ^ _17289;
  wire _17291 = _7632 ^ _5046;
  wire _17292 = _2028 ^ _14290;
  wire _17293 = _17291 ^ _17292;
  wire _17294 = uncoded_block[826] ^ uncoded_block[831];
  wire _17295 = _17294 ^ _4331;
  wire _17296 = _12138 ^ _4337;
  wire _17297 = _17295 ^ _17296;
  wire _17298 = _17293 ^ _17297;
  wire _17299 = _17290 ^ _17298;
  wire _17300 = _17283 ^ _17299;
  wire _17301 = _5737 ^ _8808;
  wire _17302 = _17301 ^ _14298;
  wire _17303 = _6406 ^ _8237;
  wire _17304 = uncoded_block[863] ^ uncoded_block[867];
  wire _17305 = _408 ^ _17304;
  wire _17306 = _17303 ^ _17305;
  wire _17307 = _17302 ^ _17306;
  wire _17308 = _3608 ^ _11056;
  wire _17309 = _13792 ^ _17308;
  wire _17310 = _11059 ^ _10506;
  wire _17311 = _5758 ^ _3617;
  wire _17312 = _17310 ^ _17311;
  wire _17313 = _17309 ^ _17312;
  wire _17314 = _17307 ^ _17313;
  wire _17315 = _9960 ^ _15345;
  wire _17316 = _6428 ^ _3625;
  wire _17317 = _17315 ^ _17316;
  wire _17318 = uncoded_block[917] ^ uncoded_block[921];
  wire _17319 = _17318 ^ _445;
  wire _17320 = _1295 ^ _448;
  wire _17321 = _17319 ^ _17320;
  wire _17322 = _17317 ^ _17321;
  wire _17323 = _2862 ^ _2083;
  wire _17324 = _12723 ^ _460;
  wire _17325 = _17323 ^ _17324;
  wire _17326 = _8277 ^ _4385;
  wire _17327 = _9977 ^ _17326;
  wire _17328 = _17325 ^ _17327;
  wire _17329 = _17322 ^ _17328;
  wire _17330 = _17314 ^ _17329;
  wire _17331 = _17300 ^ _17330;
  wire _17332 = _17265 ^ _17331;
  wire _17333 = _17193 ^ _17332;
  wire _17334 = _11646 ^ _11648;
  wire _17335 = _2877 ^ _3657;
  wire _17336 = _17334 ^ _17335;
  wire _17337 = _2100 ^ _5792;
  wire _17338 = _17337 ^ _8289;
  wire _17339 = _17336 ^ _17338;
  wire _17340 = uncoded_block[993] ^ uncoded_block[996];
  wire _17341 = _17340 ^ _11101;
  wire _17342 = _2111 ^ _486;
  wire _17343 = _17341 ^ _17342;
  wire _17344 = uncoded_block[1010] ^ uncoded_block[1014];
  wire _17345 = _17344 ^ _9996;
  wire _17346 = _2893 ^ _14855;
  wire _17347 = _17345 ^ _17346;
  wire _17348 = _17343 ^ _17347;
  wire _17349 = _17339 ^ _17348;
  wire _17350 = _8301 ^ _1339;
  wire _17351 = uncoded_block[1031] ^ uncoded_block[1035];
  wire _17352 = _17351 ^ _12198;
  wire _17353 = _17350 ^ _17352;
  wire _17354 = _12199 ^ _8309;
  wire _17355 = _1357 ^ _2136;
  wire _17356 = _17354 ^ _17355;
  wire _17357 = _17353 ^ _17356;
  wire _17358 = _1359 ^ _7117;
  wire _17359 = _5153 ^ _10569;
  wire _17360 = _17358 ^ _17359;
  wire _17361 = _2143 ^ _8893;
  wire _17362 = uncoded_block[1077] ^ uncoded_block[1081];
  wire _17363 = uncoded_block[1083] ^ uncoded_block[1086];
  wire _17364 = _17362 ^ _17363;
  wire _17365 = _17361 ^ _17364;
  wire _17366 = _17360 ^ _17365;
  wire _17367 = _17357 ^ _17366;
  wire _17368 = _17349 ^ _17367;
  wire _17369 = uncoded_block[1089] ^ uncoded_block[1096];
  wire _17370 = _2149 ^ _17369;
  wire _17371 = _543 ^ _8910;
  wire _17372 = _17370 ^ _17371;
  wire _17373 = uncoded_block[1110] ^ uncoded_block[1114];
  wire _17374 = _17373 ^ _553;
  wire _17375 = _10028 ^ _17374;
  wire _17376 = _17372 ^ _17375;
  wire _17377 = _10587 ^ _2944;
  wire _17378 = _6499 ^ _13866;
  wire _17379 = _17377 ^ _17378;
  wire _17380 = _5856 ^ _565;
  wire _17381 = _16380 ^ _574;
  wire _17382 = _17380 ^ _17381;
  wire _17383 = _17379 ^ _17382;
  wire _17384 = _17376 ^ _17383;
  wire _17385 = _4465 ^ _2956;
  wire _17386 = uncoded_block[1151] ^ uncoded_block[1155];
  wire _17387 = _17386 ^ _578;
  wire _17388 = _17385 ^ _17387;
  wire _17389 = uncoded_block[1161] ^ uncoded_block[1164];
  wire _17390 = uncoded_block[1165] ^ uncoded_block[1167];
  wire _17391 = _17389 ^ _17390;
  wire _17392 = uncoded_block[1172] ^ uncoded_block[1174];
  wire _17393 = _10046 ^ _17392;
  wire _17394 = _17391 ^ _17393;
  wire _17395 = _17388 ^ _17394;
  wire _17396 = uncoded_block[1175] ^ uncoded_block[1177];
  wire _17397 = uncoded_block[1180] ^ uncoded_block[1183];
  wire _17398 = _17396 ^ _17397;
  wire _17399 = _17398 ^ _11167;
  wire _17400 = uncoded_block[1199] ^ uncoded_block[1202];
  wire _17401 = _11719 ^ _17400;
  wire _17402 = _5204 ^ _17401;
  wire _17403 = _17399 ^ _17402;
  wire _17404 = _17395 ^ _17403;
  wire _17405 = _17384 ^ _17404;
  wire _17406 = _17368 ^ _17405;
  wire _17407 = uncoded_block[1207] ^ uncoded_block[1213];
  wire _17408 = _2209 ^ _17407;
  wire _17409 = _2982 ^ _605;
  wire _17410 = _17408 ^ _17409;
  wire _17411 = uncoded_block[1227] ^ uncoded_block[1232];
  wire _17412 = uncoded_block[1233] ^ uncoded_block[1236];
  wire _17413 = _17411 ^ _17412;
  wire _17414 = _16405 ^ _17413;
  wire _17415 = _17410 ^ _17414;
  wire _17416 = uncoded_block[1237] ^ uncoded_block[1241];
  wire _17417 = _17416 ^ _2995;
  wire _17418 = _2997 ^ _6543;
  wire _17419 = _17417 ^ _17418;
  wire _17420 = _1455 ^ _2238;
  wire _17421 = _1458 ^ _7788;
  wire _17422 = _17420 ^ _17421;
  wire _17423 = _17419 ^ _17422;
  wire _17424 = _17415 ^ _17423;
  wire _17425 = uncoded_block[1276] ^ uncoded_block[1282];
  wire _17426 = _9538 ^ _17425;
  wire _17427 = _3797 ^ _639;
  wire _17428 = _17426 ^ _17427;
  wire _17429 = uncoded_block[1288] ^ uncoded_block[1291];
  wire _17430 = _17429 ^ _10646;
  wire _17431 = uncoded_block[1298] ^ uncoded_block[1303];
  wire _17432 = _17431 ^ _2259;
  wire _17433 = _17430 ^ _17432;
  wire _17434 = _17428 ^ _17433;
  wire _17435 = uncoded_block[1309] ^ uncoded_block[1311];
  wire _17436 = _17435 ^ _2261;
  wire _17437 = _3812 ^ _3814;
  wire _17438 = _17436 ^ _17437;
  wire _17439 = _10655 ^ _4550;
  wire _17440 = uncoded_block[1338] ^ uncoded_block[1346];
  wire _17441 = _661 ^ _17440;
  wire _17442 = _17439 ^ _17441;
  wire _17443 = _17438 ^ _17442;
  wire _17444 = _17434 ^ _17443;
  wire _17445 = _17424 ^ _17444;
  wire _17446 = _5268 ^ _14442;
  wire _17447 = _672 ^ _4559;
  wire _17448 = _17446 ^ _17447;
  wire _17449 = _1504 ^ _10668;
  wire _17450 = _3832 ^ _3054;
  wire _17451 = _17449 ^ _17450;
  wire _17452 = _17448 ^ _17451;
  wire _17453 = _2290 ^ _10108;
  wire _17454 = _17453 ^ _12312;
  wire _17455 = _5952 ^ _13416;
  wire _17456 = _4572 ^ _5293;
  wire _17457 = _17455 ^ _17456;
  wire _17458 = _17454 ^ _17457;
  wire _17459 = _17452 ^ _17458;
  wire _17460 = _2300 ^ _5961;
  wire _17461 = uncoded_block[1412] ^ uncoded_block[1413];
  wire _17462 = _17461 ^ _8438;
  wire _17463 = _17460 ^ _17462;
  wire _17464 = _11792 ^ _3853;
  wire _17465 = _5967 ^ _10684;
  wire _17466 = _17464 ^ _17465;
  wire _17467 = _17463 ^ _17466;
  wire _17468 = uncoded_block[1430] ^ uncoded_block[1433];
  wire _17469 = _17468 ^ _1534;
  wire _17470 = uncoded_block[1437] ^ uncoded_block[1438];
  wire _17471 = _17470 ^ _2319;
  wire _17472 = _17469 ^ _17471;
  wire _17473 = _716 ^ _2325;
  wire _17474 = _6620 ^ _719;
  wire _17475 = _17473 ^ _17474;
  wire _17476 = _17472 ^ _17475;
  wire _17477 = _17467 ^ _17476;
  wire _17478 = _17459 ^ _17477;
  wire _17479 = _17445 ^ _17478;
  wire _17480 = _17406 ^ _17479;
  wire _17481 = _12335 ^ _726;
  wire _17482 = _17481 ^ _5982;
  wire _17483 = uncoded_block[1472] ^ uncoded_block[1474];
  wire _17484 = _5983 ^ _17483;
  wire _17485 = uncoded_block[1475] ^ uncoded_block[1479];
  wire _17486 = _17485 ^ _1558;
  wire _17487 = _17484 ^ _17486;
  wire _17488 = _17482 ^ _17487;
  wire _17489 = uncoded_block[1490] ^ uncoded_block[1492];
  wire _17490 = _17489 ^ _13967;
  wire _17491 = _743 ^ _7258;
  wire _17492 = _17490 ^ _17491;
  wire _17493 = _1572 ^ _11264;
  wire _17494 = _7875 ^ _3115;
  wire _17495 = _17493 ^ _17494;
  wire _17496 = _17492 ^ _17495;
  wire _17497 = _17488 ^ _17496;
  wire _17498 = _14488 ^ _12352;
  wire _17499 = uncoded_block[1525] ^ uncoded_block[1528];
  wire _17500 = _17499 ^ _8474;
  wire _17501 = _17498 ^ _17500;
  wire _17502 = _16496 ^ _1589;
  wire _17503 = _7274 ^ _9067;
  wire _17504 = _17502 ^ _17503;
  wire _17505 = _17501 ^ _17504;
  wire _17506 = uncoded_block[1555] ^ uncoded_block[1558];
  wire _17507 = _17506 ^ _2372;
  wire _17508 = _1606 ^ _9080;
  wire _17509 = _17507 ^ _17508;
  wire _17510 = _4648 ^ _784;
  wire _17511 = _6034 ^ _2394;
  wire _17512 = _17510 ^ _17511;
  wire _17513 = _17509 ^ _17512;
  wire _17514 = _17505 ^ _17513;
  wire _17515 = _17497 ^ _17514;
  wire _17516 = uncoded_block[1605] ^ uncoded_block[1610];
  wire _17517 = _3151 ^ _17516;
  wire _17518 = _1622 ^ _17517;
  wire _17519 = _3157 ^ _6679;
  wire _17520 = uncoded_block[1623] ^ uncoded_block[1628];
  wire _17521 = _5383 ^ _17520;
  wire _17522 = _17519 ^ _17521;
  wire _17523 = _17518 ^ _17522;
  wire _17524 = _4667 ^ _5388;
  wire _17525 = _3946 ^ _1642;
  wire _17526 = _17524 ^ _17525;
  wire _17527 = uncoded_block[1642] ^ uncoded_block[1647];
  wire _17528 = _6689 ^ _17527;
  wire _17529 = uncoded_block[1650] ^ uncoded_block[1653];
  wire _17530 = _17529 ^ _7925;
  wire _17531 = _17528 ^ _17530;
  wire _17532 = _17526 ^ _17531;
  wire _17533 = _17523 ^ _17532;
  wire _17534 = _1653 ^ _6055;
  wire _17535 = _7319 ^ _8521;
  wire _17536 = _17534 ^ _17535;
  wire _17537 = uncoded_block[1673] ^ uncoded_block[1676];
  wire _17538 = uncoded_block[1677] ^ uncoded_block[1680];
  wire _17539 = _17537 ^ _17538;
  wire _17540 = uncoded_block[1686] ^ uncoded_block[1690];
  wire _17541 = _3187 ^ _17540;
  wire _17542 = _17539 ^ _17541;
  wire _17543 = _17536 ^ _17542;
  wire _17544 = _11325 ^ _9118;
  wire _17545 = _3973 ^ _4700;
  wire _17546 = _17544 ^ _17545;
  wire _17547 = _10778 ^ _7944;
  wire _17548 = _849 ^ _17547;
  wire _17549 = _17546 ^ _17548;
  wire _17550 = _17543 ^ _17549;
  wire _17551 = _17533 ^ _17550;
  wire _17552 = _17515 ^ _17551;
  wire _17553 = uncoded_block[1718] ^ uncoded_block[1720];
  wire _17554 = _17553 ^ uncoded_block[1721];
  wire _17555 = _17552 ^ _17554;
  wire _17556 = _17480 ^ _17555;
  wire _17557 = _17333 ^ _17556;
  wire _17558 = _3209 ^ _3;
  wire _17559 = uncoded_block[8] ^ uncoded_block[12];
  wire _17560 = _17559 ^ _3998;
  wire _17561 = _17558 ^ _17560;
  wire _17562 = uncoded_block[26] ^ uncoded_block[30];
  wire _17563 = _13537 ^ _17562;
  wire _17564 = _14569 ^ _2466;
  wire _17565 = _17563 ^ _17564;
  wire _17566 = _17561 ^ _17565;
  wire _17567 = _3230 ^ _7965;
  wire _17568 = uncoded_block[46] ^ uncoded_block[50];
  wire _17569 = _12425 ^ _17568;
  wire _17570 = _17567 ^ _17569;
  wire _17571 = _12429 ^ _1703;
  wire _17572 = _10801 ^ _9705;
  wire _17573 = _17571 ^ _17572;
  wire _17574 = _17570 ^ _17573;
  wire _17575 = _17566 ^ _17574;
  wire _17576 = _7367 ^ _897;
  wire _17577 = _17576 ^ _6751;
  wire _17578 = uncoded_block[85] ^ uncoded_block[86];
  wire _17579 = _17578 ^ _14065;
  wire _17580 = _903 ^ _6115;
  wire _17581 = _17579 ^ _17580;
  wire _17582 = _17577 ^ _17581;
  wire _17583 = uncoded_block[101] ^ uncoded_block[104];
  wire _17584 = uncoded_block[105] ^ uncoded_block[106];
  wire _17585 = _17583 ^ _17584;
  wire _17586 = _14069 ^ _17585;
  wire _17587 = uncoded_block[108] ^ uncoded_block[117];
  wire _17588 = _17587 ^ _14602;
  wire _17589 = _3255 ^ _13017;
  wire _17590 = _17588 ^ _17589;
  wire _17591 = _17586 ^ _17590;
  wire _17592 = _17582 ^ _17591;
  wire _17593 = _17575 ^ _17592;
  wire _17594 = _1735 ^ _15112;
  wire _17595 = _9729 ^ _15114;
  wire _17596 = _17594 ^ _17595;
  wire _17597 = _4046 ^ _15622;
  wire _17598 = _15623 ^ _4048;
  wire _17599 = _17597 ^ _17598;
  wire _17600 = _17596 ^ _17599;
  wire _17601 = _4049 ^ _74;
  wire _17602 = _8591 ^ _1756;
  wire _17603 = _17601 ^ _17602;
  wire _17604 = _940 ^ _5479;
  wire _17605 = _7408 ^ _6798;
  wire _17606 = _17604 ^ _17605;
  wire _17607 = _17603 ^ _17606;
  wire _17608 = _17600 ^ _17607;
  wire _17609 = _2532 ^ _9745;
  wire _17610 = _6805 ^ _3291;
  wire _17611 = _17609 ^ _17610;
  wire _17612 = _8600 ^ _98;
  wire _17613 = uncoded_block[216] ^ uncoded_block[219];
  wire _17614 = _17613 ^ _5492;
  wire _17615 = _17612 ^ _17614;
  wire _17616 = _17611 ^ _17615;
  wire _17617 = uncoded_block[223] ^ uncoded_block[225];
  wire _17618 = _17617 ^ _4791;
  wire _17619 = _17618 ^ _11948;
  wire _17620 = _12495 ^ _5503;
  wire _17621 = uncoded_block[246] ^ uncoded_block[253];
  wire _17622 = _6179 ^ _17621;
  wire _17623 = _17620 ^ _17622;
  wire _17624 = _17619 ^ _17623;
  wire _17625 = _17616 ^ _17624;
  wire _17626 = _17608 ^ _17625;
  wire _17627 = _17593 ^ _17626;
  wire _17628 = uncoded_block[254] ^ uncoded_block[257];
  wire _17629 = uncoded_block[259] ^ uncoded_block[265];
  wire _17630 = _17628 ^ _17629;
  wire _17631 = uncoded_block[267] ^ uncoded_block[280];
  wire _17632 = _17631 ^ _11967;
  wire _17633 = _17630 ^ _17632;
  wire _17634 = _1803 ^ _994;
  wire _17635 = uncoded_block[295] ^ uncoded_block[297];
  wire _17636 = _995 ^ _17635;
  wire _17637 = _17634 ^ _17636;
  wire _17638 = _17633 ^ _17637;
  wire _17639 = uncoded_block[304] ^ uncoded_block[307];
  wire _17640 = _4111 ^ _17639;
  wire _17641 = _6203 ^ _17640;
  wire _17642 = uncoded_block[314] ^ uncoded_block[316];
  wire _17643 = _13619 ^ _17642;
  wire _17644 = _17643 ^ _15676;
  wire _17645 = _17641 ^ _17644;
  wire _17646 = _17638 ^ _17645;
  wire _17647 = _3347 ^ _9235;
  wire _17648 = _2587 ^ _13629;
  wire _17649 = _17647 ^ _17648;
  wire _17650 = _158 ^ _6218;
  wire _17651 = uncoded_block[349] ^ uncoded_block[354];
  wire _17652 = _1023 ^ _17651;
  wire _17653 = _17650 ^ _17652;
  wire _17654 = _17649 ^ _17653;
  wire _17655 = _9249 ^ _2606;
  wire _17656 = _11463 ^ _15183;
  wire _17657 = _17655 ^ _17656;
  wire _17658 = uncoded_block[369] ^ uncoded_block[372];
  wire _17659 = _17658 ^ _10895;
  wire _17660 = uncoded_block[376] ^ uncoded_block[381];
  wire _17661 = uncoded_block[382] ^ uncoded_block[386];
  wire _17662 = _17660 ^ _17661;
  wire _17663 = _17659 ^ _17662;
  wire _17664 = _17657 ^ _17663;
  wire _17665 = _17654 ^ _17664;
  wire _17666 = _17646 ^ _17665;
  wire _17667 = _3383 ^ _1847;
  wire _17668 = uncoded_block[399] ^ uncoded_block[402];
  wire _17669 = _10910 ^ _17668;
  wire _17670 = _17667 ^ _17669;
  wire _17671 = _15697 ^ _13106;
  wire _17672 = uncoded_block[415] ^ uncoded_block[419];
  wire _17673 = _1054 ^ _17672;
  wire _17674 = _17671 ^ _17673;
  wire _17675 = _17670 ^ _17674;
  wire _17676 = _11477 ^ _2633;
  wire _17677 = _17676 ^ _15199;
  wire _17678 = uncoded_block[431] ^ uncoded_block[437];
  wire _17679 = _17678 ^ _1863;
  wire _17680 = _12559 ^ _208;
  wire _17681 = _17679 ^ _17680;
  wire _17682 = _17677 ^ _17681;
  wire _17683 = _17675 ^ _17682;
  wire _17684 = _1075 ^ _7504;
  wire _17685 = _2653 ^ _9281;
  wire _17686 = _17684 ^ _17685;
  wire _17687 = _221 ^ _8688;
  wire _17688 = _12024 ^ _17687;
  wire _17689 = _17686 ^ _17688;
  wire _17690 = _1085 ^ _2659;
  wire _17691 = _1090 ^ _4194;
  wire _17692 = _17690 ^ _17691;
  wire _17693 = _9837 ^ _2668;
  wire _17694 = uncoded_block[510] ^ uncoded_block[512];
  wire _17695 = _9294 ^ _17694;
  wire _17696 = _17693 ^ _17695;
  wire _17697 = _17692 ^ _17696;
  wire _17698 = _17689 ^ _17697;
  wire _17699 = _17683 ^ _17698;
  wire _17700 = _17666 ^ _17699;
  wire _17701 = _17627 ^ _17700;
  wire _17702 = uncoded_block[513] ^ uncoded_block[518];
  wire _17703 = _17702 ^ _3444;
  wire _17704 = _17703 ^ _9302;
  wire _17705 = _6929 ^ _6931;
  wire _17706 = _243 ^ _9854;
  wire _17707 = _17705 ^ _17706;
  wire _17708 = _17704 ^ _17707;
  wire _17709 = _13689 ^ _8720;
  wire _17710 = uncoded_block[557] ^ uncoded_block[561];
  wire _17711 = _1915 ^ _17710;
  wire _17712 = _17709 ^ _17711;
  wire _17713 = _258 ^ _7550;
  wire _17714 = _4223 ^ _262;
  wire _17715 = _17713 ^ _17714;
  wire _17716 = _17712 ^ _17715;
  wire _17717 = _17708 ^ _17716;
  wire _17718 = uncoded_block[577] ^ uncoded_block[582];
  wire _17719 = _17718 ^ _266;
  wire _17720 = _17719 ^ _3479;
  wire _17721 = uncoded_block[594] ^ uncoded_block[597];
  wire _17722 = _17721 ^ _3486;
  wire _17723 = _5646 ^ _2710;
  wire _17724 = _17722 ^ _17723;
  wire _17725 = _17720 ^ _17724;
  wire _17726 = _8744 ^ _13713;
  wire _17727 = _17233 ^ _17726;
  wire _17728 = _7568 ^ _12618;
  wire _17729 = _4964 ^ _6966;
  wire _17730 = _17728 ^ _17729;
  wire _17731 = _17727 ^ _17730;
  wire _17732 = _17725 ^ _17731;
  wire _17733 = _17717 ^ _17732;
  wire _17734 = _12071 ^ _14228;
  wire _17735 = _290 ^ _4249;
  wire _17736 = _17734 ^ _17735;
  wire _17737 = _2727 ^ _2729;
  wire _17738 = _6973 ^ _4975;
  wire _17739 = _17737 ^ _17738;
  wire _17740 = _17736 ^ _17739;
  wire _17741 = _14755 ^ _5670;
  wire _17742 = uncoded_block[667] ^ uncoded_block[669];
  wire _17743 = _4978 ^ _17742;
  wire _17744 = _17741 ^ _17743;
  wire _17745 = uncoded_block[673] ^ uncoded_block[674];
  wire _17746 = _2744 ^ _17745;
  wire _17747 = uncoded_block[675] ^ uncoded_block[680];
  wire _17748 = _17747 ^ _6353;
  wire _17749 = _17746 ^ _17748;
  wire _17750 = _17744 ^ _17749;
  wire _17751 = _17740 ^ _17750;
  wire _17752 = _321 ^ _6983;
  wire _17753 = uncoded_block[689] ^ uncoded_block[692];
  wire _17754 = uncoded_block[694] ^ uncoded_block[699];
  wire _17755 = _17753 ^ _17754;
  wire _17756 = _17752 ^ _17755;
  wire _17757 = uncoded_block[704] ^ uncoded_block[708];
  wire _17758 = _17757 ^ _4996;
  wire _17759 = _15286 ^ _17758;
  wire _17760 = _17756 ^ _17759;
  wire _17761 = _10452 ^ _4999;
  wire _17762 = uncoded_block[717] ^ uncoded_block[719];
  wire _17763 = _17762 ^ _341;
  wire _17764 = _17761 ^ _17763;
  wire _17765 = _15292 ^ _7001;
  wire _17766 = _8200 ^ _5006;
  wire _17767 = _17765 ^ _17766;
  wire _17768 = _17764 ^ _17767;
  wire _17769 = _17760 ^ _17768;
  wire _17770 = _17751 ^ _17769;
  wire _17771 = _17733 ^ _17770;
  wire _17772 = _2775 ^ _1210;
  wire _17773 = _12656 ^ _17772;
  wire _17774 = uncoded_block[757] ^ uncoded_block[760];
  wire _17775 = _17774 ^ _13761;
  wire _17776 = uncoded_block[767] ^ uncoded_block[769];
  wire _17777 = _13762 ^ _17776;
  wire _17778 = _17775 ^ _17777;
  wire _17779 = _17773 ^ _17778;
  wire _17780 = _11019 ^ _1221;
  wire _17781 = _9382 ^ _12673;
  wire _17782 = _17780 ^ _17781;
  wire _17783 = uncoded_block[789] ^ uncoded_block[794];
  wire _17784 = _5032 ^ _17783;
  wire _17785 = _6391 ^ _383;
  wire _17786 = _17784 ^ _17785;
  wire _17787 = _17782 ^ _17786;
  wire _17788 = _17779 ^ _17787;
  wire _17789 = _385 ^ _389;
  wire _17790 = _14287 ^ _10483;
  wire _17791 = _17789 ^ _17790;
  wire _17792 = _10485 ^ _11597;
  wire _17793 = uncoded_block[825] ^ uncoded_block[828];
  wire _17794 = _5051 ^ _17793;
  wire _17795 = _17792 ^ _17794;
  wire _17796 = _17791 ^ _17795;
  wire _17797 = uncoded_block[829] ^ uncoded_block[832];
  wire _17798 = uncoded_block[836] ^ uncoded_block[841];
  wire _17799 = _17797 ^ _17798;
  wire _17800 = uncoded_block[845] ^ uncoded_block[850];
  wire _17801 = _5058 ^ _17800;
  wire _17802 = _17799 ^ _17801;
  wire _17803 = uncoded_block[860] ^ uncoded_block[862];
  wire _17804 = uncoded_block[863] ^ uncoded_block[866];
  wire _17805 = _17803 ^ _17804;
  wire _17806 = _12147 ^ _17805;
  wire _17807 = _17802 ^ _17806;
  wire _17808 = _17796 ^ _17807;
  wire _17809 = _17788 ^ _17808;
  wire _17810 = _8244 ^ _5078;
  wire _17811 = uncoded_block[885] ^ uncoded_block[890];
  wire _17812 = _2054 ^ _17811;
  wire _17813 = _17810 ^ _17812;
  wire _17814 = _2841 ^ _429;
  wire _17815 = _431 ^ _9424;
  wire _17816 = _17814 ^ _17815;
  wire _17817 = _17813 ^ _17816;
  wire _17818 = uncoded_block[914] ^ uncoded_block[915];
  wire _17819 = _17818 ^ _2852;
  wire _17820 = uncoded_block[919] ^ uncoded_block[921];
  wire _17821 = _17820 ^ _4368;
  wire _17822 = _17819 ^ _17821;
  wire _17823 = _1295 ^ _446;
  wire _17824 = _17823 ^ _16829;
  wire _17825 = _17822 ^ _17824;
  wire _17826 = _17817 ^ _17825;
  wire _17827 = _2083 ^ _6439;
  wire _17828 = uncoded_block[945] ^ uncoded_block[948];
  wire _17829 = _17828 ^ _13266;
  wire _17830 = _17827 ^ _17829;
  wire _17831 = _1303 ^ _6441;
  wire _17832 = _11086 ^ _5785;
  wire _17833 = _17831 ^ _17832;
  wire _17834 = _17830 ^ _17833;
  wire _17835 = _1315 ^ _3657;
  wire _17836 = uncoded_block[978] ^ uncoded_block[980];
  wire _17837 = uncoded_block[981] ^ uncoded_block[988];
  wire _17838 = _17836 ^ _17837;
  wire _17839 = _17835 ^ _17838;
  wire _17840 = uncoded_block[1006] ^ uncoded_block[1010];
  wire _17841 = _4404 ^ _17840;
  wire _17842 = _4403 ^ _17841;
  wire _17843 = _17839 ^ _17842;
  wire _17844 = _17834 ^ _17843;
  wire _17845 = _17826 ^ _17844;
  wire _17846 = _17809 ^ _17845;
  wire _17847 = _17771 ^ _17846;
  wire _17848 = _17701 ^ _17847;
  wire _17849 = _8296 ^ _1331;
  wire _17850 = _8871 ^ _2120;
  wire _17851 = _17849 ^ _17850;
  wire _17852 = _498 ^ _1341;
  wire _17853 = _17852 ^ _8881;
  wire _17854 = _17851 ^ _17853;
  wire _17855 = uncoded_block[1047] ^ uncoded_block[1050];
  wire _17856 = _2133 ^ _17855;
  wire _17857 = _11678 ^ _17856;
  wire _17858 = _8311 ^ _7117;
  wire _17859 = _12210 ^ _17858;
  wire _17860 = _17857 ^ _17859;
  wire _17861 = _17854 ^ _17860;
  wire _17862 = _6483 ^ _3685;
  wire _17863 = _3689 ^ _1366;
  wire _17864 = _17862 ^ _17863;
  wire _17865 = _11125 ^ _12219;
  wire _17866 = _2928 ^ _3696;
  wire _17867 = _17865 ^ _17866;
  wire _17868 = _17864 ^ _17867;
  wire _17869 = _1374 ^ _3698;
  wire _17870 = _17869 ^ _11140;
  wire _17871 = uncoded_block[1101] ^ uncoded_block[1110];
  wire _17872 = _17871 ^ _4451;
  wire _17873 = _5175 ^ _10587;
  wire _17874 = _17872 ^ _17873;
  wire _17875 = _17870 ^ _17874;
  wire _17876 = _17868 ^ _17875;
  wire _17877 = _17861 ^ _17876;
  wire _17878 = _2944 ^ _558;
  wire _17879 = _17878 ^ _5857;
  wire _17880 = uncoded_block[1137] ^ uncoded_block[1141];
  wire _17881 = _17880 ^ _1400;
  wire _17882 = uncoded_block[1150] ^ uncoded_block[1153];
  wire _17883 = _4465 ^ _17882;
  wire _17884 = _17881 ^ _17883;
  wire _17885 = _17879 ^ _17884;
  wire _17886 = uncoded_block[1156] ^ uncoded_block[1164];
  wire _17887 = _3727 ^ _17886;
  wire _17888 = _5193 ^ _11160;
  wire _17889 = _17887 ^ _17888;
  wire _17890 = uncoded_block[1174] ^ uncoded_block[1177];
  wire _17891 = _10602 ^ _17890;
  wire _17892 = uncoded_block[1178] ^ uncoded_block[1182];
  wire _17893 = _17892 ^ _4486;
  wire _17894 = _17891 ^ _17893;
  wire _17895 = _17889 ^ _17894;
  wire _17896 = _17885 ^ _17895;
  wire _17897 = _9508 ^ _2201;
  wire _17898 = uncoded_block[1195] ^ uncoded_block[1197];
  wire _17899 = _7159 ^ _17898;
  wire _17900 = _17897 ^ _17899;
  wire _17901 = _11721 ^ _2974;
  wire _17902 = _16399 ^ _7166;
  wire _17903 = _17901 ^ _17902;
  wire _17904 = _17900 ^ _17903;
  wire _17905 = _3762 ^ _2219;
  wire _17906 = _17905 ^ _14408;
  wire _17907 = uncoded_block[1224] ^ uncoded_block[1230];
  wire _17908 = uncoded_block[1231] ^ uncoded_block[1238];
  wire _17909 = _17907 ^ _17908;
  wire _17910 = uncoded_block[1240] ^ uncoded_block[1242];
  wire _17911 = uncoded_block[1245] ^ uncoded_block[1248];
  wire _17912 = _17910 ^ _17911;
  wire _17913 = _17909 ^ _17912;
  wire _17914 = _17906 ^ _17913;
  wire _17915 = _17904 ^ _17914;
  wire _17916 = _17896 ^ _17915;
  wire _17917 = _17877 ^ _17916;
  wire _17918 = _621 ^ _3001;
  wire _17919 = uncoded_block[1259] ^ uncoded_block[1263];
  wire _17920 = _7780 ^ _17919;
  wire _17921 = _17918 ^ _17920;
  wire _17922 = _3786 ^ _7179;
  wire _17923 = _17922 ^ _5909;
  wire _17924 = _17921 ^ _17923;
  wire _17925 = _631 ^ _638;
  wire _17926 = uncoded_block[1285] ^ uncoded_block[1297];
  wire _17927 = uncoded_block[1298] ^ uncoded_block[1300];
  wire _17928 = _17926 ^ _17927;
  wire _17929 = _17925 ^ _17928;
  wire _17930 = _2255 ^ _3807;
  wire _17931 = _4539 ^ _9552;
  wire _17932 = _17930 ^ _17931;
  wire _17933 = _17929 ^ _17932;
  wire _17934 = _17924 ^ _17933;
  wire _17935 = _8411 ^ _657;
  wire _17936 = _17935 ^ _14947;
  wire _17937 = _5259 ^ _1497;
  wire _17938 = uncoded_block[1343] ^ uncoded_block[1346];
  wire _17939 = uncoded_block[1347] ^ uncoded_block[1353];
  wire _17940 = _17938 ^ _17939;
  wire _17941 = _17937 ^ _17940;
  wire _17942 = _17936 ^ _17941;
  wire _17943 = _5272 ^ _12300;
  wire _17944 = _17943 ^ _2285;
  wire _17945 = uncoded_block[1371] ^ uncoded_block[1373];
  wire _17946 = _10668 ^ _17945;
  wire _17947 = _2289 ^ _5284;
  wire _17948 = _17946 ^ _17947;
  wire _17949 = _17944 ^ _17948;
  wire _17950 = _17942 ^ _17949;
  wire _17951 = _17934 ^ _17950;
  wire _17952 = _3058 ^ _3834;
  wire _17953 = uncoded_block[1385] ^ uncoded_block[1389];
  wire _17954 = _17953 ^ _2293;
  wire _17955 = _17952 ^ _17954;
  wire _17956 = _1517 ^ _2299;
  wire _17957 = _7226 ^ _17956;
  wire _17958 = _17955 ^ _17957;
  wire _17959 = _5957 ^ _4580;
  wire _17960 = uncoded_block[1418] ^ uncoded_block[1419];
  wire _17961 = _17960 ^ _16463;
  wire _17962 = _17959 ^ _17961;
  wire _17963 = uncoded_block[1425] ^ uncoded_block[1428];
  wire _17964 = _9022 ^ _17963;
  wire _17965 = _5299 ^ _10690;
  wire _17966 = _17964 ^ _17965;
  wire _17967 = _17962 ^ _17966;
  wire _17968 = _17958 ^ _17967;
  wire _17969 = _2318 ^ _5304;
  wire _17970 = _2321 ^ _1543;
  wire _17971 = _17969 ^ _17970;
  wire _17972 = _2328 ^ _2335;
  wire _17973 = _2336 ^ _3094;
  wire _17974 = _17972 ^ _17973;
  wire _17975 = _17971 ^ _17974;
  wire _17976 = uncoded_block[1469] ^ uncoded_block[1472];
  wire _17977 = _1550 ^ _17976;
  wire _17978 = _14989 ^ _2342;
  wire _17979 = _17977 ^ _17978;
  wire _17980 = uncoded_block[1486] ^ uncoded_block[1488];
  wire _17981 = _9042 ^ _17980;
  wire _17982 = _11809 ^ _12896;
  wire _17983 = _17981 ^ _17982;
  wire _17984 = _17979 ^ _17983;
  wire _17985 = _17975 ^ _17984;
  wire _17986 = _17968 ^ _17985;
  wire _17987 = _17951 ^ _17986;
  wire _17988 = _17917 ^ _17987;
  wire _17989 = _5993 ^ _1572;
  wire _17990 = _15512 ^ _17989;
  wire _17991 = _11264 ^ _6637;
  wire _17992 = _6642 ^ _5337;
  wire _17993 = _17991 ^ _17992;
  wire _17994 = _17990 ^ _17993;
  wire _17995 = _1582 ^ _11820;
  wire _17996 = _7879 ^ _17995;
  wire _17997 = _6650 ^ _16010;
  wire _17998 = uncoded_block[1544] ^ uncoded_block[1550];
  wire _17999 = _17998 ^ _767;
  wire _18000 = _17997 ^ _17999;
  wire _18001 = _17996 ^ _18000;
  wire _18002 = _17994 ^ _18001;
  wire _18003 = _3131 ^ _4638;
  wire _18004 = _4640 ^ _776;
  wire _18005 = _18003 ^ _18004;
  wire _18006 = _11284 ^ _5363;
  wire _18007 = _9080 ^ _1608;
  wire _18008 = _18006 ^ _18007;
  wire _18009 = _18005 ^ _18008;
  wire _18010 = uncoded_block[1583] ^ uncoded_block[1589];
  wire _18011 = _13479 ^ _18010;
  wire _18012 = _6673 ^ _11294;
  wire _18013 = _18011 ^ _18012;
  wire _18014 = _11295 ^ _3151;
  wire _18015 = _3153 ^ _2396;
  wire _18016 = _18014 ^ _18015;
  wire _18017 = _18013 ^ _18016;
  wire _18018 = _18009 ^ _18017;
  wire _18019 = _18002 ^ _18018;
  wire _18020 = uncoded_block[1618] ^ uncoded_block[1619];
  wire _18021 = _16032 ^ _18020;
  wire _18022 = _2399 ^ _18021;
  wire _18023 = uncoded_block[1620] ^ uncoded_block[1623];
  wire _18024 = _18023 ^ _6046;
  wire _18025 = _18024 ^ _1640;
  wire _18026 = _18022 ^ _18025;
  wire _18027 = _5392 ^ _13500;
  wire _18028 = _5394 ^ _2412;
  wire _18029 = _18027 ^ _18028;
  wire _18030 = uncoded_block[1652] ^ uncoded_block[1653];
  wire _18031 = _14530 ^ _18030;
  wire _18032 = _10760 ^ _822;
  wire _18033 = _18031 ^ _18032;
  wire _18034 = _18029 ^ _18033;
  wire _18035 = _18026 ^ _18034;
  wire _18036 = _6055 ^ _17032;
  wire _18037 = uncoded_block[1676] ^ uncoded_block[1680];
  wire _18038 = _1656 ^ _18037;
  wire _18039 = _18036 ^ _18038;
  wire _18040 = _3187 ^ _837;
  wire _18041 = uncoded_block[1693] ^ uncoded_block[1695];
  wire _18042 = _9115 ^ _18041;
  wire _18043 = _18040 ^ _18042;
  wire _18044 = _18039 ^ _18043;
  wire _18045 = uncoded_block[1697] ^ uncoded_block[1700];
  wire _18046 = _18045 ^ _14028;
  wire _18047 = _18046 ^ _3198;
  wire _18048 = _852 ^ _14552;
  wire _18049 = _18048 ^ _5416;
  wire _18050 = _18047 ^ _18049;
  wire _18051 = _18044 ^ _18050;
  wire _18052 = _18035 ^ _18051;
  wire _18053 = _18019 ^ _18052;
  wire _18054 = _17988 ^ _18053;
  wire _18055 = _17848 ^ _18054;
  wire _18056 = uncoded_block[0] ^ uncoded_block[6];
  wire _18057 = uncoded_block[8] ^ uncoded_block[10];
  wire _18058 = _18056 ^ _18057;
  wire _18059 = _7 ^ _7956;
  wire _18060 = _18058 ^ _18059;
  wire _18061 = _8545 ^ _2458;
  wire _18062 = _13539 ^ _15;
  wire _18063 = _18061 ^ _18062;
  wire _18064 = _18060 ^ _18063;
  wire _18065 = _879 ^ _2466;
  wire _18066 = _3230 ^ _17065;
  wire _18067 = _18065 ^ _18066;
  wire _18068 = _6099 ^ _1699;
  wire _18069 = _4014 ^ _5436;
  wire _18070 = _18068 ^ _18069;
  wire _18071 = _18067 ^ _18070;
  wire _18072 = _18064 ^ _18071;
  wire _18073 = _26 ^ _12435;
  wire _18074 = _18073 ^ _36;
  wire _18075 = _5442 ^ _3243;
  wire _18076 = uncoded_block[81] ^ uncoded_block[85];
  wire _18077 = uncoded_block[86] ^ uncoded_block[88];
  wire _18078 = _18076 ^ _18077;
  wire _18079 = _18075 ^ _18078;
  wire _18080 = _18074 ^ _18079;
  wire _18081 = _903 ^ _907;
  wire _18082 = _46 ^ _9718;
  wire _18083 = _18081 ^ _18082;
  wire _18084 = _15101 ^ _9166;
  wire _18085 = _2491 ^ _1726;
  wire _18086 = _18084 ^ _18085;
  wire _18087 = _18083 ^ _18086;
  wire _18088 = _18080 ^ _18087;
  wire _18089 = _18072 ^ _18088;
  wire _18090 = uncoded_block[116] ^ uncoded_block[119];
  wire _18091 = _10816 ^ _18090;
  wire _18092 = _12451 ^ _3255;
  wire _18093 = _18091 ^ _18092;
  wire _18094 = _9175 ^ _923;
  wire _18095 = uncoded_block[136] ^ uncoded_block[139];
  wire _18096 = _926 ^ _18095;
  wire _18097 = _18094 ^ _18096;
  wire _18098 = _18093 ^ _18097;
  wire _18099 = uncoded_block[141] ^ uncoded_block[147];
  wire _18100 = uncoded_block[148] ^ uncoded_block[152];
  wire _18101 = _18099 ^ _18100;
  wire _18102 = _7397 ^ _5470;
  wire _18103 = _18101 ^ _18102;
  wire _18104 = _6785 ^ _6787;
  wire _18105 = uncoded_block[170] ^ uncoded_block[177];
  wire _18106 = _18105 ^ _85;
  wire _18107 = _18104 ^ _18106;
  wire _18108 = _18103 ^ _18107;
  wire _18109 = _18098 ^ _18108;
  wire _18110 = uncoded_block[180] ^ uncoded_block[183];
  wire _18111 = uncoded_block[187] ^ uncoded_block[189];
  wire _18112 = _18110 ^ _18111;
  wire _18113 = uncoded_block[190] ^ uncoded_block[192];
  wire _18114 = _18113 ^ _2532;
  wire _18115 = _18112 ^ _18114;
  wire _18116 = _9745 ^ _4779;
  wire _18117 = _14101 ^ _98;
  wire _18118 = _18116 ^ _18117;
  wire _18119 = _18115 ^ _18118;
  wire _18120 = _4785 ^ _960;
  wire _18121 = _5492 ^ _9206;
  wire _18122 = _18120 ^ _18121;
  wire _18123 = uncoded_block[230] ^ uncoded_block[234];
  wire _18124 = _6168 ^ _18123;
  wire _18125 = uncoded_block[235] ^ uncoded_block[238];
  wire _18126 = _18125 ^ _15144;
  wire _18127 = _18124 ^ _18126;
  wire _18128 = _18122 ^ _18127;
  wire _18129 = _18119 ^ _18128;
  wire _18130 = _18109 ^ _18129;
  wire _18131 = _18089 ^ _18130;
  wire _18132 = _1781 ^ _9761;
  wire _18133 = _18132 ^ _14119;
  wire _18134 = uncoded_block[273] ^ uncoded_block[282];
  wire _18135 = _3320 ^ _18134;
  wire _18136 = _9768 ^ _18135;
  wire _18137 = _18133 ^ _18136;
  wire _18138 = _4105 ^ _5522;
  wire _18139 = _3328 ^ _17635;
  wire _18140 = _18138 ^ _18139;
  wire _18141 = _1807 ^ _17144;
  wire _18142 = _5528 ^ _145;
  wire _18143 = _18141 ^ _18142;
  wire _18144 = _18140 ^ _18143;
  wire _18145 = _18137 ^ _18144;
  wire _18146 = _146 ^ _1814;
  wire _18147 = uncoded_block[325] ^ uncoded_block[329];
  wire _18148 = _3347 ^ _18147;
  wire _18149 = _18146 ^ _18148;
  wire _18150 = _9240 ^ _1822;
  wire _18151 = uncoded_block[342] ^ uncoded_block[346];
  wire _18152 = _9242 ^ _18151;
  wire _18153 = _18150 ^ _18152;
  wire _18154 = _18149 ^ _18153;
  wire _18155 = _1023 ^ _5541;
  wire _18156 = _15179 ^ _3361;
  wire _18157 = _18155 ^ _18156;
  wire _18158 = uncoded_block[361] ^ uncoded_block[364];
  wire _18159 = _1029 ^ _18158;
  wire _18160 = uncoded_block[367] ^ uncoded_block[371];
  wire _18161 = _7470 ^ _18160;
  wire _18162 = _18159 ^ _18161;
  wire _18163 = _18157 ^ _18162;
  wire _18164 = _18154 ^ _18163;
  wire _18165 = _18145 ^ _18164;
  wire _18166 = _4853 ^ _7474;
  wire _18167 = uncoded_block[390] ^ uncoded_block[398];
  wire _18168 = _5552 ^ _18167;
  wire _18169 = _18166 ^ _18168;
  wire _18170 = uncoded_block[399] ^ uncoded_block[407];
  wire _18171 = _18170 ^ _1052;
  wire _18172 = _3394 ^ _14682;
  wire _18173 = _18171 ^ _18172;
  wire _18174 = _18169 ^ _18173;
  wire _18175 = uncoded_block[418] ^ uncoded_block[421];
  wire _18176 = _18175 ^ _2633;
  wire _18177 = _2637 ^ _1857;
  wire _18178 = _18176 ^ _18177;
  wire _18179 = _9274 ^ _207;
  wire _18180 = _18178 ^ _18179;
  wire _18181 = _18174 ^ _18180;
  wire _18182 = _16191 ^ _3411;
  wire _18183 = _4177 ^ _2650;
  wire _18184 = _18182 ^ _18183;
  wire _18185 = _3415 ^ _2653;
  wire _18186 = _9827 ^ _8683;
  wire _18187 = _18185 ^ _18186;
  wire _18188 = _18184 ^ _18187;
  wire _18189 = _1878 ^ _6266;
  wire _18190 = uncoded_block[479] ^ uncoded_block[483];
  wire _18191 = _5590 ^ _18190;
  wire _18192 = _18189 ^ _18191;
  wire _18193 = _3432 ^ _5603;
  wire _18194 = _7517 ^ _18193;
  wire _18195 = _18192 ^ _18194;
  wire _18196 = _18188 ^ _18195;
  wire _18197 = _18181 ^ _18196;
  wire _18198 = _18165 ^ _18197;
  wire _18199 = _18131 ^ _18198;
  wire _18200 = _5604 ^ _3434;
  wire _18201 = _6921 ^ _12034;
  wire _18202 = _18200 ^ _18201;
  wire _18203 = _5611 ^ _3437;
  wire _18204 = _18203 ^ _4911;
  wire _18205 = _18202 ^ _18204;
  wire _18206 = uncoded_block[518] ^ uncoded_block[522];
  wire _18207 = _18206 ^ _6289;
  wire _18208 = uncoded_block[531] ^ uncoded_block[534];
  wire _18209 = _14716 ^ _18208;
  wire _18210 = _18207 ^ _18209;
  wire _18211 = _6932 ^ _1115;
  wire _18212 = _244 ^ _1913;
  wire _18213 = _18211 ^ _18212;
  wire _18214 = _18210 ^ _18213;
  wire _18215 = _18205 ^ _18214;
  wire _18216 = uncoded_block[555] ^ uncoded_block[560];
  wire _18217 = _18216 ^ _5633;
  wire _18218 = _3465 ^ _13697;
  wire _18219 = _18217 ^ _18218;
  wire _18220 = _10398 ^ _1932;
  wire _18221 = _18219 ^ _18220;
  wire _18222 = uncoded_block[588] ^ uncoded_block[590];
  wire _18223 = _1139 ^ _18222;
  wire _18224 = _15244 ^ _18223;
  wire _18225 = uncoded_block[593] ^ uncoded_block[598];
  wire _18226 = _2700 ^ _18225;
  wire _18227 = _7558 ^ _8738;
  wire _18228 = _18226 ^ _18227;
  wire _18229 = _18224 ^ _18228;
  wire _18230 = _18221 ^ _18229;
  wire _18231 = _18215 ^ _18230;
  wire _18232 = uncoded_block[610] ^ uncoded_block[613];
  wire _18233 = _18232 ^ _4243;
  wire _18234 = _18233 ^ _17728;
  wire _18235 = uncoded_block[627] ^ uncoded_block[630];
  wire _18236 = _18235 ^ _4255;
  wire _18237 = _2727 ^ _1164;
  wire _18238 = _18236 ^ _18237;
  wire _18239 = _18234 ^ _18238;
  wire _18240 = uncoded_block[648] ^ uncoded_block[654];
  wire _18241 = _18240 ^ _3513;
  wire _18242 = _15768 ^ _309;
  wire _18243 = _18241 ^ _18242;
  wire _18244 = _13730 ^ _16257;
  wire _18245 = _18243 ^ _18244;
  wire _18246 = _18239 ^ _18245;
  wire _18247 = uncoded_block[681] ^ uncoded_block[683];
  wire _18248 = _18247 ^ _13194;
  wire _18249 = uncoded_block[687] ^ uncoded_block[689];
  wire _18250 = uncoded_block[691] ^ uncoded_block[695];
  wire _18251 = _18249 ^ _18250;
  wire _18252 = _18248 ^ _18251;
  wire _18253 = _333 ^ _10447;
  wire _18254 = _17256 ^ _18253;
  wire _18255 = _18252 ^ _18254;
  wire _18256 = _4995 ^ _8190;
  wire _18257 = _1983 ^ _6367;
  wire _18258 = _18256 ^ _18257;
  wire _18259 = uncoded_block[721] ^ uncoded_block[725];
  wire _18260 = _18259 ^ _9905;
  wire _18261 = _3547 ^ _8775;
  wire _18262 = _18260 ^ _18261;
  wire _18263 = _18258 ^ _18262;
  wire _18264 = _18255 ^ _18263;
  wire _18265 = _18246 ^ _18264;
  wire _18266 = _18231 ^ _18265;
  wire _18267 = _10464 ^ _2777;
  wire _18268 = _12656 ^ _18267;
  wire _18269 = _7013 ^ _1215;
  wire _18270 = _9914 ^ _2781;
  wire _18271 = _18269 ^ _18270;
  wire _18272 = _18268 ^ _18271;
  wire _18273 = _13762 ^ _13215;
  wire _18274 = uncoded_block[771] ^ uncoded_block[777];
  wire _18275 = _18274 ^ _368;
  wire _18276 = _18273 ^ _18275;
  wire _18277 = uncoded_block[782] ^ uncoded_block[785];
  wire _18278 = _12669 ^ _18277;
  wire _18279 = _1224 ^ _4311;
  wire _18280 = _18278 ^ _18279;
  wire _18281 = _18276 ^ _18280;
  wire _18282 = _18272 ^ _18281;
  wire _18283 = uncoded_block[790] ^ uncoded_block[793];
  wire _18284 = _18283 ^ _382;
  wire _18285 = _18284 ^ _15813;
  wire _18286 = uncoded_block[806] ^ uncoded_block[810];
  wire _18287 = _3577 ^ _18286;
  wire _18288 = uncoded_block[813] ^ uncoded_block[818];
  wire _18289 = uncoded_block[822] ^ uncoded_block[828];
  wire _18290 = _18288 ^ _18289;
  wire _18291 = _18287 ^ _18290;
  wire _18292 = _18285 ^ _18291;
  wire _18293 = _3590 ^ _4336;
  wire _18294 = _18293 ^ _5059;
  wire _18295 = _2043 ^ _8809;
  wire _18296 = uncoded_block[853] ^ uncoded_block[860];
  wire _18297 = _18296 ^ _9948;
  wire _18298 = _18295 ^ _18297;
  wire _18299 = _18294 ^ _18298;
  wire _18300 = _18292 ^ _18299;
  wire _18301 = _18282 ^ _18300;
  wire _18302 = uncoded_block[868] ^ uncoded_block[871];
  wire _18303 = _9949 ^ _18302;
  wire _18304 = uncoded_block[874] ^ uncoded_block[880];
  wire _18305 = _18304 ^ _2054;
  wire _18306 = _18303 ^ _18305;
  wire _18307 = uncoded_block[892] ^ uncoded_block[895];
  wire _18308 = _18307 ^ _429;
  wire _18309 = _5755 ^ _18308;
  wire _18310 = _18306 ^ _18309;
  wire _18311 = uncoded_block[903] ^ uncoded_block[905];
  wire _18312 = _18311 ^ _3623;
  wire _18313 = _16312 ^ _1287;
  wire _18314 = _18312 ^ _18313;
  wire _18315 = _15840 ^ _8834;
  wire _18316 = uncoded_block[929] ^ uncoded_block[932];
  wire _18317 = _18316 ^ _1299;
  wire _18318 = _18315 ^ _18317;
  wire _18319 = _18314 ^ _18318;
  wire _18320 = _18310 ^ _18319;
  wire _18321 = _452 ^ _10523;
  wire _18322 = _8274 ^ _2869;
  wire _18323 = _18321 ^ _18322;
  wire _18324 = uncoded_block[958] ^ uncoded_block[965];
  wire _18325 = _18324 ^ _9981;
  wire _18326 = _5112 ^ _3657;
  wire _18327 = _18325 ^ _18326;
  wire _18328 = _18323 ^ _18327;
  wire _18329 = uncoded_block[980] ^ uncoded_block[984];
  wire _18330 = _11092 ^ _18329;
  wire _18331 = _12186 ^ _8856;
  wire _18332 = _18330 ^ _18331;
  wire _18333 = uncoded_block[990] ^ uncoded_block[994];
  wire _18334 = _18333 ^ _13277;
  wire _18335 = _2107 ^ _2111;
  wire _18336 = _18334 ^ _18335;
  wire _18337 = _18332 ^ _18336;
  wire _18338 = _18328 ^ _18337;
  wire _18339 = _18320 ^ _18338;
  wire _18340 = _18301 ^ _18339;
  wire _18341 = _18266 ^ _18340;
  wire _18342 = _18199 ^ _18341;
  wire _18343 = _2114 ^ _1327;
  wire _18344 = uncoded_block[1013] ^ uncoded_block[1018];
  wire _18345 = _13283 ^ _18344;
  wire _18346 = _18343 ^ _18345;
  wire _18347 = _8299 ^ _495;
  wire _18348 = _8875 ^ _4417;
  wire _18349 = _18347 ^ _18348;
  wire _18350 = _18346 ^ _18349;
  wire _18351 = uncoded_block[1038] ^ uncoded_block[1045];
  wire _18352 = _18351 ^ _3681;
  wire _18353 = _2914 ^ _1363;
  wire _18354 = _18352 ^ _18353;
  wire _18355 = _2921 ^ _12213;
  wire _18356 = _3686 ^ _18355;
  wire _18357 = _18354 ^ _18356;
  wire _18358 = _18350 ^ _18357;
  wire _18359 = uncoded_block[1074] ^ uncoded_block[1078];
  wire _18360 = _12217 ^ _18359;
  wire _18361 = uncoded_block[1079] ^ uncoded_block[1084];
  wire _18362 = _18361 ^ _1373;
  wire _18363 = _18360 ^ _18362;
  wire _18364 = _1374 ^ _11137;
  wire _18365 = uncoded_block[1099] ^ uncoded_block[1101];
  wire _18366 = _5843 ^ _18365;
  wire _18367 = _18364 ^ _18366;
  wire _18368 = _18363 ^ _18367;
  wire _18369 = _4452 ^ _7735;
  wire _18370 = _1389 ^ _13327;
  wire _18371 = uncoded_block[1128] ^ uncoded_block[1130];
  wire _18372 = _18371 ^ _561;
  wire _18373 = _18370 ^ _18372;
  wire _18374 = _18369 ^ _18373;
  wire _18375 = _18368 ^ _18374;
  wire _18376 = _18358 ^ _18375;
  wire _18377 = uncoded_block[1141] ^ uncoded_block[1144];
  wire _18378 = _9496 ^ _18377;
  wire _18379 = _10597 ^ _3725;
  wire _18380 = _18378 ^ _18379;
  wire _18381 = _8351 ^ _3733;
  wire _18382 = uncoded_block[1168] ^ uncoded_block[1172];
  wire _18383 = _7749 ^ _18382;
  wire _18384 = _18381 ^ _18383;
  wire _18385 = _18380 ^ _18384;
  wire _18386 = _585 ^ _4481;
  wire _18387 = _18386 ^ _16902;
  wire _18388 = _13883 ^ _2971;
  wire _18389 = uncoded_block[1200] ^ uncoded_block[1203];
  wire _18390 = _3750 ^ _18389;
  wire _18391 = _18388 ^ _18390;
  wire _18392 = _18387 ^ _18391;
  wire _18393 = _18385 ^ _18392;
  wire _18394 = _2210 ^ _11171;
  wire _18395 = uncoded_block[1211] ^ uncoded_block[1213];
  wire _18396 = _18395 ^ _4498;
  wire _18397 = _18394 ^ _18396;
  wire _18398 = uncoded_block[1220] ^ uncoded_block[1225];
  wire _18399 = _606 ^ _18398;
  wire _18400 = uncoded_block[1230] ^ uncoded_block[1231];
  wire _18401 = _4504 ^ _18400;
  wire _18402 = _18399 ^ _18401;
  wire _18403 = _18397 ^ _18402;
  wire _18404 = uncoded_block[1232] ^ uncoded_block[1234];
  wire _18405 = _18404 ^ _3771;
  wire _18406 = _3772 ^ _8962;
  wire _18407 = _18405 ^ _18406;
  wire _18408 = uncoded_block[1249] ^ uncoded_block[1258];
  wire _18409 = _18408 ^ _3784;
  wire _18410 = _6539 ^ _18409;
  wire _18411 = _18407 ^ _18410;
  wire _18412 = _18403 ^ _18411;
  wire _18413 = _18393 ^ _18412;
  wire _18414 = _18376 ^ _18413;
  wire _18415 = _16919 ^ _3008;
  wire _18416 = _18415 ^ _11190;
  wire _18417 = uncoded_block[1286] ^ uncoded_block[1289];
  wire _18418 = _10077 ^ _18417;
  wire _18419 = uncoded_block[1293] ^ uncoded_block[1296];
  wire _18420 = _3800 ^ _18419;
  wire _18421 = _18418 ^ _18420;
  wire _18422 = _18416 ^ _18421;
  wire _18423 = uncoded_block[1308] ^ uncoded_block[1311];
  wire _18424 = _2255 ^ _18423;
  wire _18425 = _3019 ^ _18424;
  wire _18426 = uncoded_block[1317] ^ uncoded_block[1322];
  wire _18427 = _14430 ^ _18426;
  wire _18428 = _18427 ^ _4546;
  wire _18429 = _18425 ^ _18428;
  wire _18430 = _18422 ^ _18429;
  wire _18431 = uncoded_block[1332] ^ uncoded_block[1336];
  wire _18432 = _18431 ^ _7814;
  wire _18433 = _18432 ^ _5267;
  wire _18434 = uncoded_block[1350] ^ uncoded_block[1352];
  wire _18435 = _669 ^ _18434;
  wire _18436 = uncoded_block[1353] ^ uncoded_block[1354];
  wire _18437 = _18436 ^ _12857;
  wire _18438 = _18435 ^ _18437;
  wire _18439 = _18433 ^ _18438;
  wire _18440 = _7821 ^ _11224;
  wire _18441 = _7823 ^ _5284;
  wire _18442 = _18440 ^ _18441;
  wire _18443 = _2290 ^ _3834;
  wire _18444 = uncoded_block[1386] ^ uncoded_block[1388];
  wire _18445 = _18444 ^ _692;
  wire _18446 = _18443 ^ _18445;
  wire _18447 = _18442 ^ _18446;
  wire _18448 = _18439 ^ _18447;
  wire _18449 = _18430 ^ _18448;
  wire _18450 = _694 ^ _2296;
  wire _18451 = _18450 ^ _13418;
  wire _18452 = uncoded_block[1405] ^ uncoded_block[1408];
  wire _18453 = _18452 ^ _1523;
  wire _18454 = _18453 ^ _8439;
  wire _18455 = _18451 ^ _18454;
  wire _18456 = _10120 ^ _9588;
  wire _18457 = _709 ^ _14466;
  wire _18458 = _18456 ^ _18457;
  wire _18459 = uncoded_block[1432] ^ uncoded_block[1436];
  wire _18460 = _1531 ^ _18459;
  wire _18461 = _3083 ^ _6619;
  wire _18462 = _18460 ^ _18461;
  wire _18463 = _18458 ^ _18462;
  wire _18464 = _18455 ^ _18463;
  wire _18465 = uncoded_block[1451] ^ uncoded_block[1453];
  wire _18466 = _18465 ^ _5309;
  wire _18467 = _724 ^ _726;
  wire _18468 = _18466 ^ _18467;
  wire _18469 = uncoded_block[1464] ^ uncoded_block[1469];
  wire _18470 = uncoded_block[1471] ^ uncoded_block[1474];
  wire _18471 = _18469 ^ _18470;
  wire _18472 = _3881 ^ _3100;
  wire _18473 = _18471 ^ _18472;
  wire _18474 = _18468 ^ _18473;
  wire _18475 = _3101 ^ _739;
  wire _18476 = _3103 ^ _2352;
  wire _18477 = _18475 ^ _18476;
  wire _18478 = uncoded_block[1503] ^ uncoded_block[1505];
  wire _18479 = _18478 ^ _13973;
  wire _18480 = uncoded_block[1513] ^ uncoded_block[1517];
  wire _18481 = _18480 ^ _9058;
  wire _18482 = _18479 ^ _18481;
  wire _18483 = _18477 ^ _18482;
  wire _18484 = _18474 ^ _18483;
  wire _18485 = _18464 ^ _18484;
  wire _18486 = _18449 ^ _18485;
  wire _18487 = _18414 ^ _18486;
  wire _18488 = _8474 ^ _6005;
  wire _18489 = _6648 ^ _12917;
  wire _18490 = _18488 ^ _18489;
  wire _18491 = _1589 ^ _4634;
  wire _18492 = uncoded_block[1546] ^ uncoded_block[1549];
  wire _18493 = _18492 ^ _6015;
  wire _18494 = _18491 ^ _18493;
  wire _18495 = _18490 ^ _18494;
  wire _18496 = _6016 ^ _13991;
  wire _18497 = _3141 ^ _6028;
  wire _18498 = _18496 ^ _18497;
  wire _18499 = _6029 ^ _11838;
  wire _18500 = _15031 ^ _8496;
  wire _18501 = _18499 ^ _18500;
  wire _18502 = _18498 ^ _18501;
  wire _18503 = _18495 ^ _18502;
  wire _18504 = _13486 ^ _11295;
  wire _18505 = _11847 ^ _7902;
  wire _18506 = _18504 ^ _18505;
  wire _18507 = _4662 ^ _7908;
  wire _18508 = _6679 ^ _804;
  wire _18509 = _18507 ^ _18508;
  wire _18510 = _18506 ^ _18509;
  wire _18511 = uncoded_block[1626] ^ uncoded_block[1630];
  wire _18512 = _7911 ^ _18511;
  wire _18513 = uncoded_block[1638] ^ uncoded_block[1642];
  wire _18514 = _5388 ^ _18513;
  wire _18515 = _18512 ^ _18514;
  wire _18516 = uncoded_block[1644] ^ uncoded_block[1647];
  wire _18517 = _18516 ^ _1649;
  wire _18518 = _15559 ^ _2414;
  wire _18519 = _18517 ^ _18518;
  wire _18520 = _18515 ^ _18519;
  wire _18521 = _18510 ^ _18520;
  wire _18522 = _18503 ^ _18521;
  wire _18523 = uncoded_block[1665] ^ uncoded_block[1671];
  wire _18524 = _18523 ^ _17537;
  wire _18525 = _7318 ^ _18524;
  wire _18526 = _2426 ^ _3187;
  wire _18527 = _1665 ^ _9115;
  wire _18528 = _18526 ^ _18527;
  wire _18529 = _18525 ^ _18528;
  wire _18530 = _10771 ^ _847;
  wire _18531 = uncoded_block[1711] ^ uncoded_block[1719];
  wire _18532 = _10214 ^ _18531;
  wire _18533 = _18530 ^ _18532;
  wire _18534 = _18533 ^ uncoded_block[1722];
  wire _18535 = _18529 ^ _18534;
  wire _18536 = _18522 ^ _18535;
  wire _18537 = _18487 ^ _18536;
  wire _18538 = _18342 ^ _18537;
  wire _18539 = uncoded_block[1] ^ uncoded_block[3];
  wire _18540 = _18539 ^ _15073;
  wire _18541 = uncoded_block[12] ^ uncoded_block[16];
  wire _18542 = _18541 ^ _6087;
  wire _18543 = _18540 ^ _18542;
  wire _18544 = _3217 ^ _3219;
  wire _18545 = _11343 ^ _2461;
  wire _18546 = _18544 ^ _18545;
  wire _18547 = _18543 ^ _18546;
  wire _18548 = uncoded_block[33] ^ uncoded_block[35];
  wire _18549 = uncoded_block[36] ^ uncoded_block[39];
  wire _18550 = _18548 ^ _18549;
  wire _18551 = _882 ^ _3232;
  wire _18552 = _18550 ^ _18551;
  wire _18553 = _4726 ^ _4015;
  wire _18554 = _1706 ^ _5440;
  wire _18555 = _18553 ^ _18554;
  wire _18556 = _18552 ^ _18555;
  wire _18557 = _18547 ^ _18556;
  wire _18558 = uncoded_block[76] ^ uncoded_block[81];
  wire _18559 = _10244 ^ _18558;
  wire _18560 = _17578 ^ _46;
  wire _18561 = _18559 ^ _18560;
  wire _18562 = _1722 ^ _6123;
  wire _18563 = _9719 ^ _18562;
  wire _18564 = _18561 ^ _18563;
  wire _18565 = _7990 ^ _1727;
  wire _18566 = _18565 ^ _8577;
  wire _18567 = uncoded_block[130] ^ uncoded_block[137];
  wire _18568 = _3262 ^ _18567;
  wire _18569 = _11918 ^ _11924;
  wire _18570 = _18568 ^ _18569;
  wire _18571 = _18566 ^ _18570;
  wire _18572 = _18564 ^ _18571;
  wire _18573 = _18557 ^ _18572;
  wire _18574 = _11383 ^ _71;
  wire _18575 = uncoded_block[158] ^ uncoded_block[162];
  wire _18576 = _1748 ^ _18575;
  wire _18577 = _18574 ^ _18576;
  wire _18578 = _8589 ^ _11390;
  wire _18579 = _4060 ^ _86;
  wire _18580 = _18578 ^ _18579;
  wire _18581 = _18577 ^ _18580;
  wire _18582 = _9196 ^ _6798;
  wire _18583 = uncoded_block[195] ^ uncoded_block[197];
  wire _18584 = _89 ^ _18583;
  wire _18585 = _18582 ^ _18584;
  wire _18586 = _14622 ^ _4070;
  wire _18587 = _18586 ^ _16613;
  wire _18588 = _18585 ^ _18587;
  wire _18589 = _18581 ^ _18588;
  wire _18590 = _8606 ^ _15644;
  wire _18591 = _18590 ^ _14629;
  wire _18592 = _1775 ^ _2550;
  wire _18593 = _9208 ^ _2552;
  wire _18594 = _18592 ^ _18593;
  wire _18595 = _18591 ^ _18594;
  wire _18596 = _1780 ^ _116;
  wire _18597 = _7434 ^ _3311;
  wire _18598 = _18596 ^ _18597;
  wire _18599 = _8041 ^ _7438;
  wire _18600 = uncoded_block[265] ^ uncoded_block[271];
  wire _18601 = _6831 ^ _18600;
  wire _18602 = _18599 ^ _18601;
  wire _18603 = _18598 ^ _18602;
  wire _18604 = _18595 ^ _18603;
  wire _18605 = _18589 ^ _18604;
  wire _18606 = _18573 ^ _18605;
  wire _18607 = _10872 ^ _5513;
  wire _18608 = uncoded_block[281] ^ uncoded_block[288];
  wire _18609 = _18608 ^ _10876;
  wire _18610 = _18607 ^ _18609;
  wire _18611 = uncoded_block[293] ^ uncoded_block[301];
  wire _18612 = _18611 ^ _6845;
  wire _18613 = _4115 ^ _3338;
  wire _18614 = _18612 ^ _18613;
  wire _18615 = _18610 ^ _18614;
  wire _18616 = _3340 ^ _4832;
  wire _18617 = uncoded_block[325] ^ uncoded_block[332];
  wire _18618 = _3347 ^ _18617;
  wire _18619 = _18616 ^ _18618;
  wire _18620 = _8646 ^ _6217;
  wire _18621 = uncoded_block[344] ^ uncoded_block[348];
  wire _18622 = _18621 ^ _4132;
  wire _18623 = _18620 ^ _18622;
  wire _18624 = _18619 ^ _18623;
  wire _18625 = _18615 ^ _18624;
  wire _18626 = _12530 ^ _7470;
  wire _18627 = _14666 ^ _18626;
  wire _18628 = _1835 ^ _10895;
  wire _18629 = _7474 ^ _7476;
  wire _18630 = _18628 ^ _18629;
  wire _18631 = _18627 ^ _18630;
  wire _18632 = uncoded_block[381] ^ uncoded_block[387];
  wire _18633 = uncoded_block[389] ^ uncoded_block[391];
  wire _18634 = _18632 ^ _18633;
  wire _18635 = _1046 ^ _1048;
  wire _18636 = _18634 ^ _18635;
  wire _18637 = _181 ^ _1051;
  wire _18638 = _1052 ^ _5564;
  wire _18639 = _18637 ^ _18638;
  wire _18640 = _18636 ^ _18639;
  wire _18641 = _18631 ^ _18640;
  wire _18642 = _18625 ^ _18641;
  wire _18643 = uncoded_block[420] ^ uncoded_block[425];
  wire _18644 = _5565 ^ _18643;
  wire _18645 = _16184 ^ _1857;
  wire _18646 = _18644 ^ _18645;
  wire _18647 = _4169 ^ _3408;
  wire _18648 = _1864 ^ _3411;
  wire _18649 = _18647 ^ _18648;
  wire _18650 = _18646 ^ _18649;
  wire _18651 = _1870 ^ _2653;
  wire _18652 = uncoded_block[465] ^ uncoded_block[469];
  wire _18653 = _18652 ^ _8686;
  wire _18654 = _18651 ^ _18653;
  wire _18655 = _9286 ^ _3422;
  wire _18656 = _18654 ^ _18655;
  wire _18657 = _18650 ^ _18656;
  wire _18658 = _1086 ^ _4897;
  wire _18659 = _9832 ^ _2664;
  wire _18660 = _18658 ^ _18659;
  wire _18661 = _8117 ^ _5604;
  wire _18662 = _18661 ^ _1098;
  wire _18663 = _18660 ^ _18662;
  wire _18664 = _1893 ^ _13676;
  wire _18665 = uncoded_block[517] ^ uncoded_block[521];
  wire _18666 = _8706 ^ _18665;
  wire _18667 = _18664 ^ _18666;
  wire _18668 = _6289 ^ _11513;
  wire _18669 = uncoded_block[530] ^ uncoded_block[537];
  wire _18670 = uncoded_block[541] ^ uncoded_block[547];
  wire _18671 = _18669 ^ _18670;
  wire _18672 = _18668 ^ _18671;
  wire _18673 = _18667 ^ _18672;
  wire _18674 = _18663 ^ _18673;
  wire _18675 = _18657 ^ _18674;
  wire _18676 = _18642 ^ _18675;
  wire _18677 = _18606 ^ _18676;
  wire _18678 = _8720 ^ _1122;
  wire _18679 = uncoded_block[558] ^ uncoded_block[562];
  wire _18680 = _18679 ^ _3465;
  wire _18681 = _18678 ^ _18680;
  wire _18682 = uncoded_block[566] ^ uncoded_block[568];
  wire _18683 = _18682 ^ _3468;
  wire _18684 = uncoded_block[576] ^ uncoded_block[578];
  wire _18685 = _4941 ^ _18684;
  wire _18686 = _18683 ^ _18685;
  wire _18687 = _18681 ^ _18686;
  wire _18688 = _3475 ^ _3478;
  wire _18689 = uncoded_block[589] ^ uncoded_block[592];
  wire _18690 = _18689 ^ _6316;
  wire _18691 = _18688 ^ _18690;
  wire _18692 = _4952 ^ _1145;
  wire _18693 = uncoded_block[605] ^ uncoded_block[611];
  wire _18694 = _18693 ^ _7563;
  wire _18695 = _18692 ^ _18694;
  wire _18696 = _18691 ^ _18695;
  wire _18697 = _18687 ^ _18696;
  wire _18698 = _5653 ^ _6328;
  wire _18699 = _18698 ^ _12619;
  wire _18700 = _12620 ^ _290;
  wire _18701 = _4249 ^ _8751;
  wire _18702 = _18700 ^ _18701;
  wire _18703 = _18699 ^ _18702;
  wire _18704 = uncoded_block[651] ^ uncoded_block[657];
  wire _18705 = uncoded_block[658] ^ uncoded_block[660];
  wire _18706 = _18704 ^ _18705;
  wire _18707 = _15266 ^ _18706;
  wire _18708 = _12630 ^ _309;
  wire _18709 = uncoded_block[668] ^ uncoded_block[670];
  wire _18710 = uncoded_block[671] ^ uncoded_block[680];
  wire _18711 = _18709 ^ _18710;
  wire _18712 = _18708 ^ _18711;
  wire _18713 = _18707 ^ _18712;
  wire _18714 = _18703 ^ _18713;
  wire _18715 = _18697 ^ _18714;
  wire _18716 = uncoded_block[685] ^ uncoded_block[687];
  wire _18717 = _3522 ^ _18716;
  wire _18718 = _18717 ^ _15283;
  wire _18719 = uncoded_block[696] ^ uncoded_block[698];
  wire _18720 = _328 ^ _18719;
  wire _18721 = uncoded_block[702] ^ uncoded_block[704];
  wire _18722 = _3532 ^ _18721;
  wire _18723 = _18720 ^ _18722;
  wire _18724 = _18718 ^ _18723;
  wire _18725 = uncoded_block[707] ^ uncoded_block[714];
  wire _18726 = uncoded_block[715] ^ uncoded_block[719];
  wire _18727 = _18725 ^ _18726;
  wire _18728 = _12648 ^ _3544;
  wire _18729 = _18727 ^ _18728;
  wire _18730 = uncoded_block[730] ^ uncoded_block[736];
  wire _18731 = _5693 ^ _18730;
  wire _18732 = _1996 ^ _7006;
  wire _18733 = _18731 ^ _18732;
  wire _18734 = _18729 ^ _18733;
  wire _18735 = _18724 ^ _18734;
  wire _18736 = _353 ^ _356;
  wire _18737 = _2002 ^ _12663;
  wire _18738 = _18736 ^ _18737;
  wire _18739 = _15305 ^ _359;
  wire _18740 = uncoded_block[762] ^ uncoded_block[764];
  wire _18741 = _9914 ^ _18740;
  wire _18742 = _18739 ^ _18741;
  wire _18743 = _18738 ^ _18742;
  wire _18744 = _4301 ^ _5027;
  wire _18745 = _11019 ^ _15799;
  wire _18746 = _18744 ^ _18745;
  wire _18747 = _4309 ^ _371;
  wire _18748 = _14279 ^ _18747;
  wire _18749 = _18746 ^ _18748;
  wire _18750 = _18743 ^ _18749;
  wire _18751 = _18735 ^ _18750;
  wire _18752 = _18715 ^ _18751;
  wire _18753 = _4314 ^ _375;
  wire _18754 = _5034 ^ _18753;
  wire _18755 = _3581 ^ _5041;
  wire _18756 = _8225 ^ _18755;
  wire _18757 = _18754 ^ _18756;
  wire _18758 = _2809 ^ _1246;
  wire _18759 = _14801 ^ _18758;
  wire _18760 = _1249 ^ _401;
  wire _18761 = _18760 ^ _7044;
  wire _18762 = _18759 ^ _18761;
  wire _18763 = _18757 ^ _18762;
  wire _18764 = _3600 ^ _14300;
  wire _18765 = _11049 ^ _18764;
  wire _18766 = _5747 ^ _14302;
  wire _18767 = _5752 ^ _2835;
  wire _18768 = _18766 ^ _18767;
  wire _18769 = _18765 ^ _18768;
  wire _18770 = uncoded_block[882] ^ uncoded_block[887];
  wire _18771 = _18770 ^ _12704;
  wire _18772 = _2843 ^ _18311;
  wire _18773 = _18771 ^ _18772;
  wire _18774 = _3623 ^ _6428;
  wire _18775 = uncoded_block[918] ^ uncoded_block[921];
  wire _18776 = _6430 ^ _18775;
  wire _18777 = _18774 ^ _18776;
  wire _18778 = _18773 ^ _18777;
  wire _18779 = _18769 ^ _18778;
  wire _18780 = _18763 ^ _18779;
  wire _18781 = _7075 ^ _15848;
  wire _18782 = _2856 ^ _18781;
  wire _18783 = _3641 ^ _9975;
  wire _18784 = _13266 ^ _14329;
  wire _18785 = _18783 ^ _18784;
  wire _18786 = _18782 ^ _18785;
  wire _18787 = uncoded_block[956] ^ uncoded_block[964];
  wire _18788 = _18787 ^ _2092;
  wire _18789 = _11648 ^ _8847;
  wire _18790 = _18788 ^ _18789;
  wire _18791 = _11092 ^ _2882;
  wire _18792 = _18326 ^ _18791;
  wire _18793 = _18790 ^ _18792;
  wire _18794 = _18786 ^ _18793;
  wire _18795 = _7691 ^ _1326;
  wire _18796 = _15856 ^ _18795;
  wire _18797 = _1327 ^ _18344;
  wire _18798 = _14855 ^ _8301;
  wire _18799 = _18797 ^ _18798;
  wire _18800 = _18796 ^ _18799;
  wire _18801 = uncoded_block[1026] ^ uncoded_block[1028];
  wire _18802 = _18801 ^ _4418;
  wire _18803 = _18802 ^ _10555;
  wire _18804 = _5812 ^ _515;
  wire _18805 = _13844 ^ _1359;
  wire _18806 = _18804 ^ _18805;
  wire _18807 = _18803 ^ _18806;
  wire _18808 = _18800 ^ _18807;
  wire _18809 = _18794 ^ _18808;
  wire _18810 = _18780 ^ _18809;
  wire _18811 = _18752 ^ _18810;
  wire _18812 = _18677 ^ _18811;
  wire _18813 = uncoded_block[1055] ^ uncoded_block[1061];
  wire _18814 = _18813 ^ _522;
  wire _18815 = _8888 ^ _11122;
  wire _18816 = _18814 ^ _18815;
  wire _18817 = _527 ^ _3692;
  wire _18818 = _8895 ^ _530;
  wire _18819 = _18817 ^ _18818;
  wire _18820 = _18816 ^ _18819;
  wire _18821 = _4438 ^ _13311;
  wire _18822 = _10021 ^ _11137;
  wire _18823 = _18821 ^ _18822;
  wire _18824 = _542 ^ _5846;
  wire _18825 = _8910 ^ _8914;
  wire _18826 = _18824 ^ _18825;
  wire _18827 = _18823 ^ _18826;
  wire _18828 = _18820 ^ _18827;
  wire _18829 = _2164 ^ _552;
  wire _18830 = _13322 ^ _8339;
  wire _18831 = _18829 ^ _18830;
  wire _18832 = uncoded_block[1126] ^ uncoded_block[1128];
  wire _18833 = _5176 ^ _18832;
  wire _18834 = uncoded_block[1131] ^ uncoded_block[1137];
  wire _18835 = _18834 ^ _5182;
  wire _18836 = _18833 ^ _18835;
  wire _18837 = _18831 ^ _18836;
  wire _18838 = _5184 ^ _2185;
  wire _18839 = _10037 ^ _18838;
  wire _18840 = _12244 ^ _14896;
  wire _18841 = _18839 ^ _18840;
  wire _18842 = _18837 ^ _18841;
  wire _18843 = _18828 ^ _18842;
  wire _18844 = _10046 ^ _7154;
  wire _18845 = _14901 ^ _589;
  wire _18846 = _18844 ^ _18845;
  wire _18847 = _3742 ^ _2195;
  wire _18848 = uncoded_block[1185] ^ uncoded_block[1192];
  wire _18849 = _18848 ^ _11719;
  wire _18850 = _18847 ^ _18849;
  wire _18851 = _18846 ^ _18850;
  wire _18852 = _15431 ^ _2979;
  wire _18853 = _5889 ^ _3763;
  wire _18854 = _18852 ^ _18853;
  wire _18855 = _10059 ^ _11177;
  wire _18856 = _11732 ^ _15441;
  wire _18857 = _18855 ^ _18856;
  wire _18858 = _18854 ^ _18857;
  wire _18859 = _18851 ^ _18858;
  wire _18860 = uncoded_block[1242] ^ uncoded_block[1245];
  wire _18861 = _18860 ^ _1449;
  wire _18862 = _8385 ^ _6546;
  wire _18863 = _18861 ^ _18862;
  wire _18864 = _18863 ^ _3788;
  wire _18865 = _11746 ^ _3793;
  wire _18866 = uncoded_block[1287] ^ uncoded_block[1289];
  wire _18867 = _2248 ^ _18866;
  wire _18868 = _18865 ^ _18867;
  wire _18869 = _9545 ^ _10646;
  wire _18870 = uncoded_block[1299] ^ uncoded_block[1301];
  wire _18871 = _645 ^ _18870;
  wire _18872 = _18869 ^ _18871;
  wire _18873 = _18868 ^ _18872;
  wire _18874 = _18864 ^ _18873;
  wire _18875 = _18859 ^ _18874;
  wire _18876 = _18843 ^ _18875;
  wire _18877 = _3805 ^ _3807;
  wire _18878 = _8407 ^ _2261;
  wire _18879 = _18877 ^ _18878;
  wire _18880 = _5926 ^ _9555;
  wire _18881 = _8411 ^ _16435;
  wire _18882 = _18880 ^ _18881;
  wire _18883 = _18879 ^ _18882;
  wire _18884 = _3820 ^ _661;
  wire _18885 = _4553 ^ _12854;
  wire _18886 = _18884 ^ _18885;
  wire _18887 = _5268 ^ _670;
  wire _18888 = _18436 ^ _10097;
  wire _18889 = _18887 ^ _18888;
  wire _18890 = _18886 ^ _18889;
  wire _18891 = _18883 ^ _18890;
  wire _18892 = uncoded_block[1358] ^ uncoded_block[1361];
  wire _18893 = _18892 ^ _1504;
  wire _18894 = _2284 ^ _10669;
  wire _18895 = _18893 ^ _18894;
  wire _18896 = uncoded_block[1382] ^ uncoded_block[1386];
  wire _18897 = _4564 ^ _18896;
  wire _18898 = _3838 ^ _13412;
  wire _18899 = _18897 ^ _18898;
  wire _18900 = _18895 ^ _18899;
  wire _18901 = uncoded_block[1392] ^ uncoded_block[1397];
  wire _18902 = _18901 ^ _1517;
  wire _18903 = uncoded_block[1402] ^ uncoded_block[1408];
  wire _18904 = _18903 ^ _4580;
  wire _18905 = _18902 ^ _18904;
  wire _18906 = _12322 ^ _10120;
  wire _18907 = _9022 ^ _2308;
  wire _18908 = _18906 ^ _18907;
  wire _18909 = _18905 ^ _18908;
  wire _18910 = _18900 ^ _18909;
  wire _18911 = _18891 ^ _18910;
  wire _18912 = _14977 ^ _1533;
  wire _18913 = _2318 ^ _4590;
  wire _18914 = _18912 ^ _18913;
  wire _18915 = _3865 ^ _720;
  wire _18916 = _11244 ^ _18915;
  wire _18917 = _18914 ^ _18916;
  wire _18918 = _12335 ^ _7243;
  wire _18919 = uncoded_block[1469] ^ uncoded_block[1470];
  wire _18920 = _5314 ^ _18919;
  wire _18921 = _18918 ^ _18920;
  wire _18922 = _3097 ^ _733;
  wire _18923 = _735 ^ _11807;
  wire _18924 = _18922 ^ _18923;
  wire _18925 = _18921 ^ _18924;
  wire _18926 = _18917 ^ _18925;
  wire _18927 = _16981 ^ _1565;
  wire _18928 = uncoded_block[1497] ^ uncoded_block[1502];
  wire _18929 = _3890 ^ _18928;
  wire _18930 = _18927 ^ _18929;
  wire _18931 = uncoded_block[1505] ^ uncoded_block[1510];
  wire _18932 = _1572 ^ _18931;
  wire _18933 = _6642 ^ _14488;
  wire _18934 = _18932 ^ _18933;
  wire _18935 = _18930 ^ _18934;
  wire _18936 = _11270 ^ _11272;
  wire _18937 = _9631 ^ _12914;
  wire _18938 = _18936 ^ _18937;
  wire _18939 = _15009 ^ _6651;
  wire _18940 = uncoded_block[1542] ^ uncoded_block[1555];
  wire _18941 = uncoded_block[1556] ^ uncoded_block[1561];
  wire _18942 = _18940 ^ _18941;
  wire _18943 = _18939 ^ _18942;
  wire _18944 = _18938 ^ _18943;
  wire _18945 = _18935 ^ _18944;
  wire _18946 = _18926 ^ _18945;
  wire _18947 = _18911 ^ _18946;
  wire _18948 = _18876 ^ _18947;
  wire _18949 = uncoded_block[1572] ^ uncoded_block[1575];
  wire _18950 = _18949 ^ _6663;
  wire _18951 = _7286 ^ _18950;
  wire _18952 = uncoded_block[1580] ^ uncoded_block[1582];
  wire _18953 = _18952 ^ _15537;
  wire _18954 = _10172 ^ _2394;
  wire _18955 = _18953 ^ _18954;
  wire _18956 = _18951 ^ _18955;
  wire _18957 = uncoded_block[1600] ^ uncoded_block[1603];
  wire _18958 = _8499 ^ _18957;
  wire _18959 = uncoded_block[1605] ^ uncoded_block[1609];
  wire _18960 = _18959 ^ _3937;
  wire _18961 = _18958 ^ _18960;
  wire _18962 = _18961 ^ _10184;
  wire _18963 = _18956 ^ _18962;
  wire _18964 = _6046 ^ _14525;
  wire _18965 = uncoded_block[1633] ^ uncoded_block[1636];
  wire _18966 = _15551 ^ _18965;
  wire _18967 = _18964 ^ _18966;
  wire _18968 = _5392 ^ _815;
  wire _18969 = uncoded_block[1645] ^ uncoded_block[1648];
  wire _18970 = _18969 ^ _10757;
  wire _18971 = _18968 ^ _18970;
  wire _18972 = _18967 ^ _18971;
  wire _18973 = _18030 ^ _11862;
  wire _18974 = _3175 ^ _3179;
  wire _18975 = _18973 ^ _18974;
  wire _18976 = _5399 ^ _7928;
  wire _18977 = _17537 ^ _9113;
  wire _18978 = _18976 ^ _18977;
  wire _18979 = _18975 ^ _18978;
  wire _18980 = _18972 ^ _18979;
  wire _18981 = _18963 ^ _18980;
  wire _18982 = uncoded_block[1683] ^ uncoded_block[1685];
  wire _18983 = _18982 ^ _1665;
  wire _18984 = _6707 ^ _18041;
  wire _18985 = _18983 ^ _18984;
  wire _18986 = _9677 ^ _11327;
  wire _18987 = _14028 ^ _2437;
  wire _18988 = _18986 ^ _18987;
  wire _18989 = _18985 ^ _18988;
  wire _18990 = uncoded_block[1713] ^ uncoded_block[1717];
  wire _18991 = _2438 ^ _18990;
  wire _18992 = _3988 ^ _12976;
  wire _18993 = _18991 ^ _18992;
  wire _18994 = _18993 ^ uncoded_block[1722];
  wire _18995 = _18989 ^ _18994;
  wire _18996 = _18981 ^ _18995;
  wire _18997 = _18948 ^ _18996;
  wire _18998 = _18812 ^ _18997;
  wire _18999 = uncoded_block[3] ^ uncoded_block[9];
  wire _19000 = _4710 ^ _18999;
  wire _19001 = uncoded_block[10] ^ uncoded_block[13];
  wire _19002 = _19001 ^ _868;
  wire _19003 = _19000 ^ _19002;
  wire _19004 = _12419 ^ _7354;
  wire _19005 = _19003 ^ _19004;
  wire _19006 = uncoded_block[36] ^ uncoded_block[41];
  wire _19007 = _3225 ^ _19006;
  wire _19008 = _14048 ^ _9150;
  wire _19009 = _19007 ^ _19008;
  wire _19010 = _14575 ^ _2471;
  wire _19011 = uncoded_block[61] ^ uncoded_block[65];
  wire _19012 = _7364 ^ _19011;
  wire _19013 = _19010 ^ _19012;
  wire _19014 = _19009 ^ _19013;
  wire _19015 = _19005 ^ _19014;
  wire _19016 = _11357 ^ _6745;
  wire _19017 = _4020 ^ _39;
  wire _19018 = _19016 ^ _19017;
  wire _19019 = uncoded_block[80] ^ uncoded_block[82];
  wire _19020 = _19019 ^ _14586;
  wire _19021 = _2484 ^ _2487;
  wire _19022 = _19020 ^ _19021;
  wire _19023 = _19018 ^ _19022;
  wire _19024 = _1718 ^ _4026;
  wire _19025 = uncoded_block[102] ^ uncoded_block[104];
  wire _19026 = _10251 ^ _19025;
  wire _19027 = _19024 ^ _19026;
  wire _19028 = _8572 ^ _5453;
  wire _19029 = uncoded_block[115] ^ uncoded_block[124];
  wire _19030 = _6763 ^ _19029;
  wire _19031 = _19028 ^ _19030;
  wire _19032 = _19027 ^ _19031;
  wire _19033 = _19023 ^ _19032;
  wire _19034 = _19015 ^ _19033;
  wire _19035 = uncoded_block[128] ^ uncoded_block[132];
  wire _19036 = uncoded_block[136] ^ uncoded_block[141];
  wire _19037 = _19035 ^ _19036;
  wire _19038 = _4046 ^ _15623;
  wire _19039 = _19037 ^ _19038;
  wire _19040 = uncoded_block[159] ^ uncoded_block[161];
  wire _19041 = _6784 ^ _19040;
  wire _19042 = uncoded_block[162] ^ uncoded_block[167];
  wire _19043 = _19042 ^ _8591;
  wire _19044 = _19041 ^ _19043;
  wire _19045 = _19039 ^ _19044;
  wire _19046 = _82 ^ _9195;
  wire _19047 = _7402 ^ _19046;
  wire _19048 = uncoded_block[185] ^ uncoded_block[193];
  wire _19049 = _19048 ^ _3284;
  wire _19050 = uncoded_block[200] ^ uncoded_block[209];
  wire _19051 = _2532 ^ _19050;
  wire _19052 = _19049 ^ _19051;
  wire _19053 = _19047 ^ _19052;
  wire _19054 = _19045 ^ _19053;
  wire _19055 = _4787 ^ _5497;
  wire _19056 = _14625 ^ _19055;
  wire _19057 = _2545 ^ _6168;
  wire _19058 = _6821 ^ _968;
  wire _19059 = _19057 ^ _19058;
  wire _19060 = _19056 ^ _19059;
  wire _19061 = uncoded_block[253] ^ uncoded_block[258];
  wire _19062 = _1781 ^ _19061;
  wire _19063 = _3306 ^ _19062;
  wire _19064 = _7438 ^ _6187;
  wire _19065 = _14122 ^ _6192;
  wire _19066 = _19064 ^ _19065;
  wire _19067 = _19063 ^ _19066;
  wire _19068 = _19060 ^ _19067;
  wire _19069 = _19054 ^ _19068;
  wire _19070 = _19034 ^ _19069;
  wire _19071 = uncoded_block[276] ^ uncoded_block[281];
  wire _19072 = uncoded_block[283] ^ uncoded_block[285];
  wire _19073 = _19071 ^ _19072;
  wire _19074 = _992 ^ _995;
  wire _19075 = _19073 ^ _19074;
  wire _19076 = _13615 ^ _8636;
  wire _19077 = uncoded_block[304] ^ uncoded_block[309];
  wire _19078 = _142 ^ _19077;
  wire _19079 = _19076 ^ _19078;
  wire _19080 = _19075 ^ _19079;
  wire _19081 = _14654 ^ _11439;
  wire _19082 = _6208 ^ _11441;
  wire _19083 = _19081 ^ _19082;
  wire _19084 = _4123 ^ _12521;
  wire _19085 = _4838 ^ _2592;
  wire _19086 = _19084 ^ _19085;
  wire _19087 = _19083 ^ _19086;
  wire _19088 = _19080 ^ _19087;
  wire _19089 = _1825 ^ _6859;
  wire _19090 = _161 ^ _4132;
  wire _19091 = _19089 ^ _19090;
  wire _19092 = uncoded_block[352] ^ uncoded_block[354];
  wire _19093 = _19092 ^ _5548;
  wire _19094 = _7470 ^ _13093;
  wire _19095 = _19093 ^ _19094;
  wire _19096 = _19091 ^ _19095;
  wire _19097 = _6873 ^ _10895;
  wire _19098 = _8079 ^ _2609;
  wire _19099 = _19097 ^ _19098;
  wire _19100 = _1038 ^ _3377;
  wire _19101 = _3380 ^ _7483;
  wire _19102 = _19100 ^ _19101;
  wire _19103 = _19099 ^ _19102;
  wire _19104 = _19096 ^ _19103;
  wire _19105 = _19088 ^ _19104;
  wire _19106 = uncoded_block[400] ^ uncoded_block[408];
  wire _19107 = _19106 ^ _14682;
  wire _19108 = _18635 ^ _19107;
  wire _19109 = _13112 ^ _4163;
  wire _19110 = _4164 ^ _11479;
  wire _19111 = _19109 ^ _19110;
  wire _19112 = _19108 ^ _19111;
  wire _19113 = uncoded_block[434] ^ uncoded_block[438];
  wire _19114 = _12553 ^ _19113;
  wire _19115 = uncoded_block[439] ^ uncoded_block[442];
  wire _19116 = _19115 ^ _12559;
  wire _19117 = _19114 ^ _19116;
  wire _19118 = uncoded_block[448] ^ uncoded_block[450];
  wire _19119 = _19118 ^ _4177;
  wire _19120 = _1075 ^ _1870;
  wire _19121 = _19119 ^ _19120;
  wire _19122 = _19117 ^ _19121;
  wire _19123 = _19112 ^ _19122;
  wire _19124 = _3415 ^ _5586;
  wire _19125 = _4185 ^ _13665;
  wire _19126 = _19124 ^ _19125;
  wire _19127 = _4188 ^ _11494;
  wire _19128 = uncoded_block[478] ^ uncoded_block[481];
  wire _19129 = _5590 ^ _19128;
  wire _19130 = _19127 ^ _19129;
  wire _19131 = _19126 ^ _19130;
  wire _19132 = _1086 ^ _12577;
  wire _19133 = _12578 ^ _9837;
  wire _19134 = _19132 ^ _19133;
  wire _19135 = uncoded_block[501] ^ uncoded_block[502];
  wire _19136 = _19135 ^ _6921;
  wire _19137 = _10376 ^ _4908;
  wire _19138 = _19136 ^ _19137;
  wire _19139 = _19134 ^ _19138;
  wire _19140 = _19131 ^ _19139;
  wire _19141 = _19123 ^ _19140;
  wire _19142 = _19105 ^ _19141;
  wire _19143 = _19070 ^ _19142;
  wire _19144 = _13676 ^ _17205;
  wire _19145 = _19144 ^ _3446;
  wire _19146 = _14716 ^ _1111;
  wire _19147 = _9309 ^ _6292;
  wire _19148 = _19146 ^ _19147;
  wire _19149 = _19145 ^ _19148;
  wire _19150 = _8718 ^ _1909;
  wire _19151 = _19150 ^ _1914;
  wire _19152 = _1123 ^ _4937;
  wire _19153 = uncoded_block[565] ^ uncoded_block[568];
  wire _19154 = _9319 ^ _19153;
  wire _19155 = _19152 ^ _19154;
  wire _19156 = _19151 ^ _19155;
  wire _19157 = _19149 ^ _19156;
  wire _19158 = _3468 ^ _3472;
  wire _19159 = _6312 ^ _8733;
  wire _19160 = _19158 ^ _19159;
  wire _19161 = _3479 ^ _2702;
  wire _19162 = _19160 ^ _19161;
  wire _19163 = uncoded_block[599] ^ uncoded_block[605];
  wire _19164 = _2706 ^ _19163;
  wire _19165 = _1942 ^ _8154;
  wire _19166 = _19164 ^ _19165;
  wire _19167 = _4960 ^ _14224;
  wire _19168 = _7565 ^ _19167;
  wire _19169 = _19166 ^ _19168;
  wire _19170 = _19162 ^ _19169;
  wire _19171 = _19157 ^ _19170;
  wire _19172 = uncoded_block[626] ^ uncoded_block[630];
  wire _19173 = _19172 ^ _14228;
  wire _19174 = _3501 ^ _1160;
  wire _19175 = _19173 ^ _19174;
  wire _19176 = _1163 ^ _296;
  wire _19177 = uncoded_block[648] ^ uncoded_block[650];
  wire _19178 = _19177 ^ _1960;
  wire _19179 = _19176 ^ _19178;
  wire _19180 = _19175 ^ _19179;
  wire _19181 = uncoded_block[653] ^ uncoded_block[655];
  wire _19182 = _19181 ^ _1962;
  wire _19183 = _15768 ^ _308;
  wire _19184 = _19182 ^ _19183;
  wire _19185 = uncoded_block[673] ^ uncoded_block[675];
  wire _19186 = _311 ^ _19185;
  wire _19187 = _10991 ^ _19186;
  wire _19188 = _19184 ^ _19187;
  wire _19189 = _19180 ^ _19188;
  wire _19190 = _8177 ^ _1968;
  wire _19191 = uncoded_block[681] ^ uncoded_block[684];
  wire _19192 = _19191 ^ _15281;
  wire _19193 = _19190 ^ _19192;
  wire _19194 = uncoded_block[689] ^ uncoded_block[693];
  wire _19195 = uncoded_block[697] ^ uncoded_block[698];
  wire _19196 = _19194 ^ _19195;
  wire _19197 = uncoded_block[699] ^ uncoded_block[705];
  wire _19198 = _19197 ^ _4995;
  wire _19199 = _19196 ^ _19198;
  wire _19200 = _19193 ^ _19199;
  wire _19201 = uncoded_block[713] ^ uncoded_block[715];
  wire _19202 = _19201 ^ _12648;
  wire _19203 = _3544 ^ _10457;
  wire _19204 = _19202 ^ _19203;
  wire _19205 = _1991 ^ _5006;
  wire _19206 = _2770 ^ _5699;
  wire _19207 = _19205 ^ _19206;
  wire _19208 = _19204 ^ _19207;
  wire _19209 = _19200 ^ _19208;
  wire _19210 = _19189 ^ _19209;
  wire _19211 = _19171 ^ _19210;
  wire _19212 = uncoded_block[746] ^ uncoded_block[754];
  wire _19213 = _19212 ^ _7015;
  wire _19214 = _19213 ^ _361;
  wire _19215 = uncoded_block[764] ^ uncoded_block[769];
  wire _19216 = _19215 ^ _15310;
  wire _19217 = uncoded_block[777] ^ uncoded_block[780];
  wire _19218 = uncoded_block[785] ^ uncoded_block[788];
  wire _19219 = _19217 ^ _19218;
  wire _19220 = _19216 ^ _19219;
  wire _19221 = _19214 ^ _19220;
  wire _19222 = uncoded_block[790] ^ uncoded_block[794];
  wire _19223 = uncoded_block[796] ^ uncoded_block[799];
  wire _19224 = _19222 ^ _19223;
  wire _19225 = _12126 ^ _389;
  wire _19226 = _19224 ^ _19225;
  wire _19227 = _16791 ^ _5041;
  wire _19228 = _2806 ^ _5046;
  wire _19229 = _19227 ^ _19228;
  wire _19230 = _19226 ^ _19229;
  wire _19231 = _19221 ^ _19230;
  wire _19232 = _3587 ^ _2032;
  wire _19233 = _4331 ^ _16801;
  wire _19234 = _19232 ^ _19233;
  wire _19235 = _9938 ^ _5058;
  wire _19236 = uncoded_block[852] ^ uncoded_block[859];
  wire _19237 = _5060 ^ _19236;
  wire _19238 = _19235 ^ _19237;
  wire _19239 = _19234 ^ _19238;
  wire _19240 = _5071 ^ _2828;
  wire _19241 = _5070 ^ _19240;
  wire _19242 = _6415 ^ _7654;
  wire _19243 = _2836 ^ _1272;
  wire _19244 = _19242 ^ _19243;
  wire _19245 = _19241 ^ _19244;
  wire _19246 = _19239 ^ _19245;
  wire _19247 = _19231 ^ _19246;
  wire _19248 = _18307 ^ _8826;
  wire _19249 = _429 ^ _9960;
  wire _19250 = _19248 ^ _19249;
  wire _19251 = uncoded_block[906] ^ uncoded_block[909];
  wire _19252 = uncoded_block[910] ^ uncoded_block[912];
  wire _19253 = _19251 ^ _19252;
  wire _19254 = _6434 ^ _5766;
  wire _19255 = _19253 ^ _19254;
  wire _19256 = _19250 ^ _19255;
  wire _19257 = _4370 ^ _1296;
  wire _19258 = _2078 ^ _2862;
  wire _19259 = _19257 ^ _19258;
  wire _19260 = _7080 ^ _6439;
  wire _19261 = uncoded_block[945] ^ uncoded_block[949];
  wire _19262 = _2865 ^ _19261;
  wire _19263 = _19260 ^ _19262;
  wire _19264 = _19259 ^ _19263;
  wire _19265 = _19256 ^ _19264;
  wire _19266 = _8276 ^ _9980;
  wire _19267 = _2872 ^ _2092;
  wire _19268 = uncoded_block[971] ^ uncoded_block[973];
  wire _19269 = _11648 ^ _19268;
  wire _19270 = _19267 ^ _19269;
  wire _19271 = _19266 ^ _19270;
  wire _19272 = uncoded_block[983] ^ uncoded_block[989];
  wire _19273 = _19272 ^ _2882;
  wire _19274 = _14847 ^ _19273;
  wire _19275 = uncoded_block[992] ^ uncoded_block[994];
  wire _19276 = _19275 ^ _6453;
  wire _19277 = uncoded_block[998] ^ uncoded_block[1002];
  wire _19278 = _19277 ^ _2886;
  wire _19279 = _19276 ^ _19278;
  wire _19280 = _19274 ^ _19279;
  wire _19281 = _19271 ^ _19280;
  wire _19282 = _19265 ^ _19281;
  wire _19283 = _19247 ^ _19282;
  wire _19284 = _19211 ^ _19283;
  wire _19285 = _19143 ^ _19284;
  wire _19286 = uncoded_block[1016] ^ uncoded_block[1020];
  wire _19287 = _19286 ^ _1334;
  wire _19288 = _7695 ^ _19287;
  wire _19289 = uncoded_block[1023] ^ uncoded_block[1027];
  wire _19290 = uncoded_block[1028] ^ uncoded_block[1033];
  wire _19291 = _19289 ^ _19290;
  wire _19292 = _7707 ^ _12199;
  wire _19293 = _19291 ^ _19292;
  wire _19294 = _19288 ^ _19293;
  wire _19295 = uncoded_block[1048] ^ uncoded_block[1050];
  wire _19296 = _19295 ^ _2136;
  wire _19297 = _19296 ^ _1361;
  wire _19298 = uncoded_block[1060] ^ uncoded_block[1063];
  wire _19299 = _19298 ^ _2142;
  wire _19300 = uncoded_block[1068] ^ uncoded_block[1078];
  wire _19301 = uncoded_block[1079] ^ uncoded_block[1082];
  wire _19302 = _19300 ^ _19301;
  wire _19303 = _19299 ^ _19302;
  wire _19304 = _19297 ^ _19303;
  wire _19305 = _19294 ^ _19304;
  wire _19306 = uncoded_block[1087] ^ uncoded_block[1091];
  wire _19307 = _2928 ^ _19306;
  wire _19308 = _19307 ^ _4443;
  wire _19309 = _5843 ^ _5169;
  wire _19310 = _19309 ^ _7732;
  wire _19311 = _19308 ^ _19310;
  wire _19312 = _549 ^ _4450;
  wire _19313 = uncoded_block[1115] ^ uncoded_block[1117];
  wire _19314 = _4451 ^ _19313;
  wire _19315 = _19312 ^ _19314;
  wire _19316 = _8920 ^ _5176;
  wire _19317 = _2944 ^ _18832;
  wire _19318 = _19316 ^ _19317;
  wire _19319 = _19315 ^ _19318;
  wire _19320 = _19311 ^ _19319;
  wire _19321 = _19305 ^ _19320;
  wire _19322 = uncoded_block[1129] ^ uncoded_block[1133];
  wire _19323 = _19322 ^ _5856;
  wire _19324 = _10593 ^ _5182;
  wire _19325 = _19323 ^ _19324;
  wire _19326 = _1400 ^ _5862;
  wire _19327 = _8933 ^ _5188;
  wire _19328 = _19326 ^ _19327;
  wire _19329 = _19325 ^ _19328;
  wire _19330 = uncoded_block[1157] ^ uncoded_block[1161];
  wire _19331 = _19330 ^ _3734;
  wire _19332 = _11160 ^ _10602;
  wire _19333 = _19331 ^ _19332;
  wire _19334 = _17396 ^ _5873;
  wire _19335 = _5200 ^ _3746;
  wire _19336 = _19334 ^ _19335;
  wire _19337 = _19333 ^ _19336;
  wire _19338 = _19329 ^ _19337;
  wire _19339 = uncoded_block[1187] ^ uncoded_block[1190];
  wire _19340 = _19339 ^ _3749;
  wire _19341 = _14398 ^ _2206;
  wire _19342 = _19340 ^ _19341;
  wire _19343 = _2207 ^ _5885;
  wire _19344 = _7765 ^ _16403;
  wire _19345 = _19343 ^ _19344;
  wire _19346 = _19342 ^ _19345;
  wire _19347 = uncoded_block[1220] ^ uncoded_block[1224];
  wire _19348 = _14914 ^ _19347;
  wire _19349 = _11177 ^ _1439;
  wire _19350 = _19348 ^ _19349;
  wire _19351 = _2225 ^ _14921;
  wire _19352 = _19351 ^ _5222;
  wire _19353 = _19350 ^ _19352;
  wire _19354 = _19346 ^ _19353;
  wire _19355 = _19338 ^ _19354;
  wire _19356 = _19321 ^ _19355;
  wire _19357 = _6536 ^ _6538;
  wire _19358 = uncoded_block[1251] ^ uncoded_block[1254];
  wire _19359 = _19358 ^ _3783;
  wire _19360 = _19357 ^ _19359;
  wire _19361 = _3784 ^ _16919;
  wire _19362 = _19361 ^ _14929;
  wire _19363 = _19360 ^ _19362;
  wire _19364 = _7792 ^ _3793;
  wire _19365 = uncoded_block[1283] ^ uncoded_block[1286];
  wire _19366 = _3794 ^ _19365;
  wire _19367 = _19364 ^ _19366;
  wire _19368 = _18866 ^ _9545;
  wire _19369 = uncoded_block[1295] ^ uncoded_block[1298];
  wire _19370 = _19369 ^ _18870;
  wire _19371 = _19368 ^ _19370;
  wire _19372 = _19367 ^ _19371;
  wire _19373 = _19363 ^ _19372;
  wire _19374 = _1481 ^ _17931;
  wire _19375 = uncoded_block[1323] ^ uncoded_block[1325];
  wire _19376 = _5254 ^ _19375;
  wire _19377 = uncoded_block[1326] ^ uncoded_block[1329];
  wire _19378 = _19377 ^ _5256;
  wire _19379 = _19376 ^ _19378;
  wire _19380 = _19374 ^ _19379;
  wire _19381 = _661 ^ _3038;
  wire _19382 = uncoded_block[1353] ^ uncoded_block[1358];
  wire _19383 = _12855 ^ _19382;
  wire _19384 = _19381 ^ _19383;
  wire _19385 = _6588 ^ _677;
  wire _19386 = _19385 ^ _9011;
  wire _19387 = _19384 ^ _19386;
  wire _19388 = _19380 ^ _19387;
  wire _19389 = _19373 ^ _19388;
  wire _19390 = _684 ^ _12305;
  wire _19391 = uncoded_block[1377] ^ uncoded_block[1384];
  wire _19392 = _19391 ^ _12867;
  wire _19393 = _19390 ^ _19392;
  wire _19394 = uncoded_block[1392] ^ uncoded_block[1398];
  wire _19395 = _19394 ^ _3841;
  wire _19396 = _3068 ^ _13947;
  wire _19397 = _19395 ^ _19396;
  wire _19398 = _19393 ^ _19397;
  wire _19399 = _15972 ^ _2306;
  wire _19400 = _11792 ^ _1527;
  wire _19401 = _19399 ^ _19400;
  wire _19402 = _10684 ^ _3081;
  wire _19403 = _1534 ^ _712;
  wire _19404 = _19402 ^ _19403;
  wire _19405 = _19401 ^ _19404;
  wire _19406 = _19398 ^ _19405;
  wire _19407 = _2319 ^ _5305;
  wire _19408 = uncoded_block[1452] ^ uncoded_block[1456];
  wire _19409 = _1543 ^ _19408;
  wire _19410 = _19407 ^ _19409;
  wire _19411 = uncoded_block[1461] ^ uncoded_block[1468];
  wire _19412 = _13437 ^ _19411;
  wire _19413 = _5983 ^ _3097;
  wire _19414 = _19412 ^ _19413;
  wire _19415 = _19410 ^ _19414;
  wire _19416 = uncoded_block[1476] ^ uncoded_block[1483];
  wire _19417 = _19416 ^ _739;
  wire _19418 = _1563 ^ _2352;
  wire _19419 = _19417 ^ _19418;
  wire _19420 = _747 ^ _7866;
  wire _19421 = uncoded_block[1505] ^ uncoded_block[1511];
  wire _19422 = _1572 ^ _19421;
  wire _19423 = _19420 ^ _19422;
  wire _19424 = _19419 ^ _19423;
  wire _19425 = _19415 ^ _19424;
  wire _19426 = _19406 ^ _19425;
  wire _19427 = _19389 ^ _19426;
  wire _19428 = _19356 ^ _19427;
  wire _19429 = uncoded_block[1512] ^ uncoded_block[1514];
  wire _19430 = _19429 ^ _9621;
  wire _19431 = uncoded_block[1517] ^ uncoded_block[1523];
  wire _19432 = _19431 ^ _1581;
  wire _19433 = _19430 ^ _19432;
  wire _19434 = _11272 ^ _9631;
  wire _19435 = _9064 ^ _3906;
  wire _19436 = _19434 ^ _19435;
  wire _19437 = _19433 ^ _19436;
  wire _19438 = _8482 ^ _14496;
  wire _19439 = _16500 ^ _19438;
  wire _19440 = _4638 ^ _4644;
  wire _19441 = _6658 ^ _19440;
  wire _19442 = _19439 ^ _19441;
  wire _19443 = _19437 ^ _19442;
  wire _19444 = _4645 ^ _4647;
  wire _19445 = _15535 ^ _6031;
  wire _19446 = _19444 ^ _19445;
  wire _19447 = _2386 ^ _3927;
  wire _19448 = uncoded_block[1591] ^ uncoded_block[1595];
  wire _19449 = _19448 ^ _8499;
  wire _19450 = _19447 ^ _19449;
  wire _19451 = _19446 ^ _19450;
  wire _19452 = _14517 ^ _10743;
  wire _19453 = _7297 ^ _6684;
  wire _19454 = _19452 ^ _19453;
  wire _19455 = uncoded_block[1624] ^ uncoded_block[1630];
  wire _19456 = _19455 ^ _5388;
  wire _19457 = _9099 ^ _7309;
  wire _19458 = _19456 ^ _19457;
  wire _19459 = _19454 ^ _19458;
  wire _19460 = _19451 ^ _19459;
  wire _19461 = _19443 ^ _19460;
  wire _19462 = _3169 ^ _2412;
  wire _19463 = _3172 ^ _18030;
  wire _19464 = _19462 ^ _19463;
  wire _19465 = _13508 ^ _4680;
  wire _19466 = uncoded_block[1664] ^ uncoded_block[1666];
  wire _19467 = _3175 ^ _19466;
  wire _19468 = _19465 ^ _19467;
  wire _19469 = _19464 ^ _19468;
  wire _19470 = uncoded_block[1667] ^ uncoded_block[1669];
  wire _19471 = uncoded_block[1670] ^ uncoded_block[1672];
  wire _19472 = _19470 ^ _19471;
  wire _19473 = _7323 ^ _5401;
  wire _19474 = _19472 ^ _19473;
  wire _19475 = uncoded_block[1684] ^ uncoded_block[1687];
  wire _19476 = _19475 ^ _837;
  wire _19477 = _17039 ^ _19476;
  wire _19478 = _19474 ^ _19477;
  wire _19479 = _19469 ^ _19478;
  wire _19480 = _6707 ^ _840;
  wire _19481 = _18045 ^ _4700;
  wire _19482 = _19480 ^ _19481;
  wire _19483 = uncoded_block[1706] ^ uncoded_block[1714];
  wire _19484 = _3976 ^ _19483;
  wire _19485 = _2441 ^ _2443;
  wire _19486 = _19484 ^ _19485;
  wire _19487 = _19482 ^ _19486;
  wire _19488 = _19487 ^ uncoded_block[1719];
  wire _19489 = _19479 ^ _19488;
  wire _19490 = _19461 ^ _19489;
  wire _19491 = _19428 ^ _19490;
  wire _19492 = _19285 ^ _19491;
  wire _19493 = _4710 ^ _3993;
  wire _19494 = _4 ^ _1686;
  wire _19495 = _19493 ^ _19494;
  wire _19496 = uncoded_block[20] ^ uncoded_block[22];
  wire _19497 = _9692 ^ _19496;
  wire _19498 = _3220 ^ _15;
  wire _19499 = _19497 ^ _19498;
  wire _19500 = _19495 ^ _19499;
  wire _19501 = uncoded_block[35] ^ uncoded_block[37];
  wire _19502 = _19501 ^ _19;
  wire _19503 = _6736 ^ _6099;
  wire _19504 = _19502 ^ _19503;
  wire _19505 = _6101 ^ _1700;
  wire _19506 = uncoded_block[57] ^ uncoded_block[61];
  wire _19507 = _888 ^ _19506;
  wire _19508 = _19505 ^ _19507;
  wire _19509 = _19504 ^ _19508;
  wire _19510 = _19500 ^ _19509;
  wire _19511 = uncoded_block[72] ^ uncoded_block[75];
  wire _19512 = _34 ^ _19511;
  wire _19513 = _19512 ^ _17076;
  wire _19514 = _14586 ^ _14065;
  wire _19515 = uncoded_block[90] ^ uncoded_block[93];
  wire _19516 = _19515 ^ _6758;
  wire _19517 = _19514 ^ _19516;
  wire _19518 = _19513 ^ _19517;
  wire _19519 = _9718 ^ _7986;
  wire _19520 = uncoded_block[109] ^ uncoded_block[111];
  wire _19521 = _6122 ^ _19520;
  wire _19522 = _19519 ^ _19521;
  wire _19523 = _6763 ^ _6769;
  wire _19524 = _19523 ^ _2499;
  wire _19525 = _19522 ^ _19524;
  wire _19526 = _19518 ^ _19525;
  wire _19527 = _19510 ^ _19526;
  wire _19528 = _9727 ^ _8579;
  wire _19529 = _2510 ^ _3265;
  wire _19530 = _19528 ^ _19529;
  wire _19531 = uncoded_block[149] ^ uncoded_block[154];
  wire _19532 = _19531 ^ _3271;
  wire _19533 = _17096 ^ _19532;
  wire _19534 = _19530 ^ _19533;
  wire _19535 = _73 ^ _19040;
  wire _19536 = uncoded_block[163] ^ uncoded_block[166];
  wire _19537 = _19536 ^ _6788;
  wire _19538 = _19535 ^ _19537;
  wire _19539 = uncoded_block[173] ^ uncoded_block[174];
  wire _19540 = _81 ^ _19539;
  wire _19541 = _19540 ^ _12471;
  wire _19542 = _19538 ^ _19541;
  wire _19543 = _19534 ^ _19542;
  wire _19544 = uncoded_block[189] ^ uncoded_block[193];
  wire _19545 = _4772 ^ _19544;
  wire _19546 = uncoded_block[201] ^ uncoded_block[205];
  wire _19547 = _2532 ^ _19546;
  wire _19548 = _19545 ^ _19547;
  wire _19549 = uncoded_block[211] ^ uncoded_block[213];
  wire _19550 = _19549 ^ _8606;
  wire _19551 = _16613 ^ _19550;
  wire _19552 = _19548 ^ _19551;
  wire _19553 = _102 ^ _4788;
  wire _19554 = _4076 ^ _3299;
  wire _19555 = _19553 ^ _19554;
  wire _19556 = _3303 ^ _3305;
  wire _19557 = _8612 ^ _11952;
  wire _19558 = _19556 ^ _19557;
  wire _19559 = _19555 ^ _19558;
  wire _19560 = _19552 ^ _19559;
  wire _19561 = _19543 ^ _19560;
  wire _19562 = _19527 ^ _19561;
  wire _19563 = _974 ^ _3311;
  wire _19564 = _14639 ^ _119;
  wire _19565 = _19563 ^ _19564;
  wire _19566 = uncoded_block[271] ^ uncoded_block[274];
  wire _19567 = _984 ^ _19566;
  wire _19568 = _4805 ^ _19567;
  wire _19569 = _19565 ^ _19568;
  wire _19570 = uncoded_block[275] ^ uncoded_block[277];
  wire _19571 = _19570 ^ _7445;
  wire _19572 = _10304 ^ _991;
  wire _19573 = _19571 ^ _19572;
  wire _19574 = uncoded_block[288] ^ uncoded_block[292];
  wire _19575 = _19574 ^ _2573;
  wire _19576 = _17142 ^ _143;
  wire _19577 = _19575 ^ _19576;
  wire _19578 = _19573 ^ _19577;
  wire _19579 = _19569 ^ _19578;
  wire _19580 = _149 ^ _6852;
  wire _19581 = _10316 ^ _19580;
  wire _19582 = _2584 ^ _4125;
  wire _19583 = uncoded_block[333] ^ uncoded_block[339];
  wire _19584 = _19583 ^ _4129;
  wire _19585 = _19582 ^ _19584;
  wire _19586 = _19581 ^ _19585;
  wire _19587 = _7465 ^ _5541;
  wire _19588 = _162 ^ _6221;
  wire _19589 = _19587 ^ _19588;
  wire _19590 = uncoded_block[368] ^ uncoded_block[371];
  wire _19591 = _17163 ^ _19590;
  wire _19592 = _16660 ^ _19591;
  wire _19593 = _19589 ^ _19592;
  wire _19594 = _19586 ^ _19593;
  wire _19595 = _19579 ^ _19594;
  wire _19596 = _13094 ^ _10898;
  wire _19597 = _10899 ^ _4857;
  wire _19598 = _19596 ^ _19597;
  wire _19599 = uncoded_block[385] ^ uncoded_block[387];
  wire _19600 = _3377 ^ _19599;
  wire _19601 = _3381 ^ _2615;
  wire _19602 = _19600 ^ _19601;
  wire _19603 = _19598 ^ _19602;
  wire _19604 = uncoded_block[392] ^ uncoded_block[394];
  wire _19605 = _19604 ^ _3384;
  wire _19606 = _1849 ^ _2625;
  wire _19607 = _19605 ^ _19606;
  wire _19608 = _6244 ^ _13106;
  wire _19609 = _19608 ^ _8664;
  wire _19610 = _19607 ^ _19609;
  wire _19611 = _19603 ^ _19610;
  wire _19612 = uncoded_block[413] ^ uncoded_block[415];
  wire _19613 = uncoded_block[417] ^ uncoded_block[420];
  wire _19614 = _19612 ^ _19613;
  wire _19615 = _19614 ^ _8673;
  wire _19616 = _13115 ^ _10352;
  wire _19617 = uncoded_block[436] ^ uncoded_block[442];
  wire _19618 = _19617 ^ _10356;
  wire _19619 = _19616 ^ _19618;
  wire _19620 = _19615 ^ _19619;
  wire _19621 = uncoded_block[451] ^ uncoded_block[454];
  wire _19622 = _3411 ^ _19621;
  wire _19623 = _1870 ^ _13127;
  wire _19624 = _19622 ^ _19623;
  wire _19625 = uncoded_block[472] ^ uncoded_block[476];
  wire _19626 = _1874 ^ _19625;
  wire _19627 = _5598 ^ _1090;
  wire _19628 = _19626 ^ _19627;
  wire _19629 = _19624 ^ _19628;
  wire _19630 = _19620 ^ _19629;
  wire _19631 = _19611 ^ _19630;
  wire _19632 = _19595 ^ _19631;
  wire _19633 = _19562 ^ _19632;
  wire _19634 = _1091 ^ _3432;
  wire _19635 = _6919 ^ _12033;
  wire _19636 = _19634 ^ _19635;
  wire _19637 = _2671 ^ _8701;
  wire _19638 = uncoded_block[518] ^ uncoded_block[519];
  wire _19639 = _9840 ^ _19638;
  wire _19640 = _19637 ^ _19639;
  wire _19641 = _19636 ^ _19640;
  wire _19642 = uncoded_block[522] ^ uncoded_block[531];
  wire _19643 = _1107 ^ _19642;
  wire _19644 = _5617 ^ _8718;
  wire _19645 = _19643 ^ _19644;
  wire _19646 = _16715 ^ _8720;
  wire _19647 = _8724 ^ _6940;
  wire _19648 = _19646 ^ _19647;
  wire _19649 = _19645 ^ _19648;
  wire _19650 = _19641 ^ _19649;
  wire _19651 = _9319 ^ _18682;
  wire _19652 = uncoded_block[576] ^ uncoded_block[579];
  wire _19653 = _4224 ^ _19652;
  wire _19654 = _19651 ^ _19653;
  wire _19655 = _1138 ^ _8733;
  wire _19656 = uncoded_block[587] ^ uncoded_block[591];
  wire _19657 = _19656 ^ _8148;
  wire _19658 = _19655 ^ _19657;
  wire _19659 = _19654 ^ _19658;
  wire _19660 = _8149 ^ _2707;
  wire _19661 = _2710 ^ _12609;
  wire _19662 = _19660 ^ _19661;
  wire _19663 = _8744 ^ _6959;
  wire _19664 = _6960 ^ _4246;
  wire _19665 = _19663 ^ _19664;
  wire _19666 = _19662 ^ _19665;
  wire _19667 = _19659 ^ _19666;
  wire _19668 = _19650 ^ _19667;
  wire _19669 = uncoded_block[628] ^ uncoded_block[635];
  wire _19670 = _2720 ^ _19669;
  wire _19671 = _293 ^ _8751;
  wire _19672 = _19670 ^ _19671;
  wire _19673 = _296 ^ _15766;
  wire _19674 = uncoded_block[655] ^ uncoded_block[661];
  wire _19675 = _4975 ^ _19674;
  wire _19676 = _19673 ^ _19675;
  wire _19677 = _19672 ^ _19676;
  wire _19678 = _12630 ^ _1177;
  wire _19679 = _19678 ^ _8178;
  wire _19680 = _1971 ^ _6353;
  wire _19681 = _4271 ^ _326;
  wire _19682 = _19680 ^ _19681;
  wire _19683 = _19679 ^ _19682;
  wire _19684 = _19677 ^ _19683;
  wire _19685 = _6985 ^ _8186;
  wire _19686 = _4275 ^ _18721;
  wire _19687 = _19685 ^ _19686;
  wire _19688 = uncoded_block[708] ^ uncoded_block[711];
  wire _19689 = _19688 ^ _3536;
  wire _19690 = _12647 ^ _5002;
  wire _19691 = _19689 ^ _19690;
  wire _19692 = _19687 ^ _19691;
  wire _19693 = _5690 ^ _6374;
  wire _19694 = _1990 ^ _7605;
  wire _19695 = _19693 ^ _19694;
  wire _19696 = _4293 ^ _1214;
  wire _19697 = _12105 ^ _19696;
  wire _19698 = _19695 ^ _19697;
  wire _19699 = _19692 ^ _19698;
  wire _19700 = _19684 ^ _19699;
  wire _19701 = _19668 ^ _19700;
  wire _19702 = _5017 ^ _4299;
  wire _19703 = _19702 ^ _14782;
  wire _19704 = _2784 ^ _11019;
  wire _19705 = uncoded_block[778] ^ uncoded_block[781];
  wire _19706 = _7620 ^ _19705;
  wire _19707 = _19704 ^ _19706;
  wire _19708 = _19703 ^ _19707;
  wire _19709 = uncoded_block[787] ^ uncoded_block[792];
  wire _19710 = _2015 ^ _19709;
  wire _19711 = _11024 ^ _11591;
  wire _19712 = _19710 ^ _19711;
  wire _19713 = _2801 ^ _5726;
  wire _19714 = _19713 ^ _8229;
  wire _19715 = _19712 ^ _19714;
  wire _19716 = _19708 ^ _19715;
  wire _19717 = uncoded_block[815] ^ uncoded_block[821];
  wire _19718 = _19717 ^ _1246;
  wire _19719 = _2032 ^ _2812;
  wire _19720 = _19718 ^ _19719;
  wire _19721 = _12137 ^ _1253;
  wire _19722 = _11043 ^ _2036;
  wire _19723 = _19721 ^ _19722;
  wire _19724 = _19720 ^ _19723;
  wire _19725 = uncoded_block[847] ^ uncoded_block[849];
  wire _19726 = _19725 ^ _408;
  wire _19727 = _9948 ^ _14302;
  wire _19728 = _19726 ^ _19727;
  wire _19729 = _2828 ^ _1269;
  wire _19730 = _2831 ^ _2835;
  wire _19731 = _19729 ^ _19730;
  wire _19732 = _19728 ^ _19731;
  wire _19733 = _19724 ^ _19732;
  wire _19734 = _19716 ^ _19733;
  wire _19735 = uncoded_block[894] ^ uncoded_block[896];
  wire _19736 = _421 ^ _19735;
  wire _19737 = _428 ^ _15345;
  wire _19738 = _19736 ^ _19737;
  wire _19739 = uncoded_block[912] ^ uncoded_block[919];
  wire _19740 = _1285 ^ _19739;
  wire _19741 = _3632 ^ _2855;
  wire _19742 = _19740 ^ _19741;
  wire _19743 = _19738 ^ _19742;
  wire _19744 = _7075 ^ _2079;
  wire _19745 = _5101 ^ _16832;
  wire _19746 = _19744 ^ _19745;
  wire _19747 = uncoded_block[944] ^ uncoded_block[946];
  wire _19748 = uncoded_block[951] ^ uncoded_block[954];
  wire _19749 = _19747 ^ _19748;
  wire _19750 = uncoded_block[956] ^ uncoded_block[961];
  wire _19751 = _19750 ^ _2092;
  wire _19752 = _19749 ^ _19751;
  wire _19753 = _19746 ^ _19752;
  wire _19754 = _19743 ^ _19753;
  wire _19755 = _2093 ^ _1314;
  wire _19756 = _13821 ^ _8855;
  wire _19757 = _19755 ^ _19756;
  wire _19758 = _5118 ^ _4401;
  wire _19759 = _2883 ^ _6457;
  wire _19760 = _19758 ^ _19759;
  wire _19761 = _19757 ^ _19760;
  wire _19762 = _7691 ^ _8866;
  wire _19763 = uncoded_block[1012] ^ uncoded_block[1015];
  wire _19764 = _5129 ^ _19763;
  wire _19765 = _19762 ^ _19764;
  wire _19766 = uncoded_block[1023] ^ uncoded_block[1025];
  wire _19767 = _5135 ^ _19766;
  wire _19768 = uncoded_block[1033] ^ uncoded_block[1035];
  wire _19769 = _18801 ^ _19768;
  wire _19770 = _19767 ^ _19769;
  wire _19771 = _19765 ^ _19770;
  wire _19772 = _19761 ^ _19771;
  wire _19773 = _19754 ^ _19772;
  wire _19774 = _19734 ^ _19773;
  wire _19775 = _19701 ^ _19774;
  wire _19776 = _19633 ^ _19775;
  wire _19777 = uncoded_block[1041] ^ uncoded_block[1044];
  wire _19778 = _502 ^ _19777;
  wire _19779 = _1356 ^ _10564;
  wire _19780 = _19778 ^ _19779;
  wire _19781 = _7117 ^ _13849;
  wire _19782 = uncoded_block[1063] ^ uncoded_block[1067];
  wire _19783 = _19782 ^ _8892;
  wire _19784 = _19781 ^ _19783;
  wire _19785 = _19780 ^ _19784;
  wire _19786 = _5158 ^ _2147;
  wire _19787 = _8904 ^ _7725;
  wire _19788 = _19786 ^ _19787;
  wire _19789 = _5840 ^ _537;
  wire _19790 = _10026 ^ _545;
  wire _19791 = _19789 ^ _19790;
  wire _19792 = _19788 ^ _19791;
  wire _19793 = _19785 ^ _19792;
  wire _19794 = uncoded_block[1102] ^ uncoded_block[1104];
  wire _19795 = uncoded_block[1106] ^ uncoded_block[1111];
  wire _19796 = _19794 ^ _19795;
  wire _19797 = _7133 ^ _13322;
  wire _19798 = _19796 ^ _19797;
  wire _19799 = _3714 ^ _5176;
  wire _19800 = _19799 ^ _15895;
  wire _19801 = _19798 ^ _19800;
  wire _19802 = _13866 ^ _5856;
  wire _19803 = _2177 ^ _5861;
  wire _19804 = _19802 ^ _19803;
  wire _19805 = uncoded_block[1151] ^ uncoded_block[1156];
  wire _19806 = _2956 ^ _19805;
  wire _19807 = _578 ^ _13335;
  wire _19808 = _19806 ^ _19807;
  wire _19809 = _19804 ^ _19808;
  wire _19810 = _19801 ^ _19809;
  wire _19811 = _19793 ^ _19810;
  wire _19812 = _10602 ^ _5872;
  wire _19813 = _590 ^ _1418;
  wire _19814 = _19812 ^ _19813;
  wire _19815 = uncoded_block[1192] ^ uncoded_block[1195];
  wire _19816 = _2971 ^ _19815;
  wire _19817 = _7160 ^ _2209;
  wire _19818 = _19816 ^ _19817;
  wire _19819 = _19814 ^ _19818;
  wire _19820 = _2979 ^ _10617;
  wire _19821 = _19820 ^ _18853;
  wire _19822 = _10059 ^ _609;
  wire _19823 = _14919 ^ _14921;
  wire _19824 = _19822 ^ _19823;
  wire _19825 = _19821 ^ _19824;
  wire _19826 = _19819 ^ _19825;
  wire _19827 = uncoded_block[1237] ^ uncoded_block[1239];
  wire _19828 = _19827 ^ _6536;
  wire _19829 = uncoded_block[1243] ^ uncoded_block[1245];
  wire _19830 = _19829 ^ _1451;
  wire _19831 = _19828 ^ _19830;
  wire _19832 = _12824 ^ _7782;
  wire _19833 = _19831 ^ _19832;
  wire _19834 = uncoded_block[1268] ^ uncoded_block[1272];
  wire _19835 = _3786 ^ _19834;
  wire _19836 = _3005 ^ _19835;
  wire _19837 = _7792 ^ _7183;
  wire _19838 = _4525 ^ _15456;
  wire _19839 = _19837 ^ _19838;
  wire _19840 = _19836 ^ _19839;
  wire _19841 = _19833 ^ _19840;
  wire _19842 = _19826 ^ _19841;
  wire _19843 = _19811 ^ _19842;
  wire _19844 = uncoded_block[1297] ^ uncoded_block[1306];
  wire _19845 = _9547 ^ _19844;
  wire _19846 = _1480 ^ _14432;
  wire _19847 = _19845 ^ _19846;
  wire _19848 = _9555 ^ _7201;
  wire _19849 = _1494 ^ _4551;
  wire _19850 = _19848 ^ _19849;
  wire _19851 = _19847 ^ _19850;
  wire _19852 = _3822 ^ _5262;
  wire _19853 = _11771 ^ _12857;
  wire _19854 = _19852 ^ _19853;
  wire _19855 = _6588 ^ _5275;
  wire _19856 = _3047 ^ _3052;
  wire _19857 = _19855 ^ _19856;
  wire _19858 = _19854 ^ _19857;
  wire _19859 = _19851 ^ _19858;
  wire _19860 = _8423 ^ _9573;
  wire _19861 = uncoded_block[1383] ^ uncoded_block[1386];
  wire _19862 = _3834 ^ _19861;
  wire _19863 = _19860 ^ _19862;
  wire _19864 = uncoded_block[1390] ^ uncoded_block[1395];
  wire _19865 = _691 ^ _19864;
  wire _19866 = uncoded_block[1398] ^ uncoded_block[1405];
  wire _19867 = _13938 ^ _19866;
  wire _19868 = _19865 ^ _19867;
  wire _19869 = _19863 ^ _19868;
  wire _19870 = _2300 ^ _6606;
  wire _19871 = _13422 ^ _1526;
  wire _19872 = _19870 ^ _19871;
  wire _19873 = _709 ^ _3081;
  wire _19874 = _19873 ^ _16968;
  wire _19875 = _19872 ^ _19874;
  wire _19876 = _19869 ^ _19875;
  wire _19877 = _19859 ^ _19876;
  wire _19878 = _3084 ^ _11246;
  wire _19879 = _719 ^ _6622;
  wire _19880 = _19878 ^ _19879;
  wire _19881 = _723 ^ _8455;
  wire _19882 = uncoded_block[1465] ^ uncoded_block[1469];
  wire _19883 = _19882 ^ _16977;
  wire _19884 = _19881 ^ _19883;
  wire _19885 = _19880 ^ _19884;
  wire _19886 = _1555 ^ _13963;
  wire _19887 = uncoded_block[1483] ^ uncoded_block[1486];
  wire _19888 = _19887 ^ _7251;
  wire _19889 = _19886 ^ _19888;
  wire _19890 = uncoded_block[1496] ^ uncoded_block[1501];
  wire _19891 = _17489 ^ _19890;
  wire _19892 = uncoded_block[1506] ^ uncoded_block[1510];
  wire _19893 = _19892 ^ _19429;
  wire _19894 = _19891 ^ _19893;
  wire _19895 = _19889 ^ _19894;
  wire _19896 = _19885 ^ _19895;
  wire _19897 = uncoded_block[1518] ^ uncoded_block[1522];
  wire _19898 = _9621 ^ _19897;
  wire _19899 = uncoded_block[1523] ^ uncoded_block[1527];
  wire _19900 = uncoded_block[1528] ^ uncoded_block[1533];
  wire _19901 = _19899 ^ _19900;
  wire _19902 = _19898 ^ _19901;
  wire _19903 = uncoded_block[1536] ^ uncoded_block[1540];
  wire _19904 = _19903 ^ _6008;
  wire _19905 = _5355 ^ _8482;
  wire _19906 = _19904 ^ _19905;
  wire _19907 = _19902 ^ _19906;
  wire _19908 = _14496 ^ _15528;
  wire _19909 = _15022 ^ _5361;
  wire _19910 = _19908 ^ _19909;
  wire _19911 = _14506 ^ _3921;
  wire _19912 = _18006 ^ _19911;
  wire _19913 = _19910 ^ _19912;
  wire _19914 = _19907 ^ _19913;
  wire _19915 = _19896 ^ _19914;
  wire _19916 = _19877 ^ _19915;
  wire _19917 = _19843 ^ _19916;
  wire _19918 = uncoded_block[1582] ^ uncoded_block[1587];
  wire _19919 = _19918 ^ _5371;
  wire _19920 = _19919 ^ _14516;
  wire _19921 = uncoded_block[1601] ^ uncoded_block[1608];
  wire _19922 = _19921 ^ _3937;
  wire _19923 = _16032 ^ _12376;
  wire _19924 = _19922 ^ _19923;
  wire _19925 = _19920 ^ _19924;
  wire _19926 = _7912 ^ _3941;
  wire _19927 = _807 ^ _14525;
  wire _19928 = _19926 ^ _19927;
  wire _19929 = uncoded_block[1631] ^ uncoded_block[1633];
  wire _19930 = _19929 ^ _2405;
  wire _19931 = uncoded_block[1637] ^ uncoded_block[1642];
  wire _19932 = _19931 ^ _3169;
  wire _19933 = _19930 ^ _19932;
  wire _19934 = _19928 ^ _19933;
  wire _19935 = _19925 ^ _19934;
  wire _19936 = _18030 ^ _820;
  wire _19937 = _3174 ^ _823;
  wire _19938 = _19936 ^ _19937;
  wire _19939 = uncoded_block[1669] ^ uncoded_block[1671];
  wire _19940 = _17032 ^ _19939;
  wire _19941 = _6700 ^ _1662;
  wire _19942 = _19940 ^ _19941;
  wire _19943 = _19938 ^ _19942;
  wire _19944 = _4691 ^ _6705;
  wire _19945 = _2429 ^ _11325;
  wire _19946 = _19944 ^ _19945;
  wire _19947 = _840 ^ _5409;
  wire _19948 = _845 ^ _8536;
  wire _19949 = _19947 ^ _19948;
  wire _19950 = _19946 ^ _19949;
  wire _19951 = _19943 ^ _19950;
  wire _19952 = _19935 ^ _19951;
  wire _19953 = uncoded_block[1709] ^ uncoded_block[1713];
  wire _19954 = _19953 ^ _7944;
  wire _19955 = _19954 ^ _10217;
  wire _19956 = _19952 ^ _19955;
  wire _19957 = _19917 ^ _19956;
  wire _19958 = _19776 ^ _19957;
  wire _19959 = uncoded_block[7] ^ uncoded_block[9];
  wire _19960 = _4712 ^ _19959;
  wire _19961 = _6086 ^ _871;
  wire _19962 = _19960 ^ _19961;
  wire _19963 = uncoded_block[20] ^ uncoded_block[23];
  wire _19964 = _10226 ^ _19963;
  wire _19965 = uncoded_block[27] ^ uncoded_block[32];
  wire _19966 = _4001 ^ _19965;
  wire _19967 = _19964 ^ _19966;
  wire _19968 = _19962 ^ _19967;
  wire _19969 = _16 ^ _18;
  wire _19970 = _19 ^ _8554;
  wire _19971 = _19969 ^ _19970;
  wire _19972 = uncoded_block[48] ^ uncoded_block[51];
  wire _19973 = _19972 ^ _4014;
  wire _19974 = uncoded_block[58] ^ uncoded_block[61];
  wire _19975 = _19974 ^ _2474;
  wire _19976 = _19973 ^ _19975;
  wire _19977 = _19971 ^ _19976;
  wire _19978 = _19968 ^ _19977;
  wire _19979 = _1706 ^ _3241;
  wire _19980 = uncoded_block[83] ^ uncoded_block[88];
  wire _19981 = _4733 ^ _19980;
  wire _19982 = _19979 ^ _19981;
  wire _19983 = _47 ^ _910;
  wire _19984 = _18081 ^ _19983;
  wire _19985 = _19982 ^ _19984;
  wire _19986 = _7986 ^ _2491;
  wire _19987 = _19986 ^ _17089;
  wire _19988 = _6128 ^ _10256;
  wire _19989 = uncoded_block[127] ^ uncoded_block[133];
  wire _19990 = _19989 ^ _926;
  wire _19991 = _19988 ^ _19990;
  wire _19992 = _19987 ^ _19991;
  wire _19993 = _19985 ^ _19992;
  wire _19994 = _19978 ^ _19993;
  wire _19995 = _4760 ^ _4043;
  wire _19996 = _7392 ^ _3269;
  wire _19997 = _19995 ^ _19996;
  wire _19998 = uncoded_block[159] ^ uncoded_block[162];
  wire _19999 = _5470 ^ _19998;
  wire _20000 = _19999 ^ _8590;
  wire _20001 = _19997 ^ _20000;
  wire _20002 = _10841 ^ _1757;
  wire _20003 = _10839 ^ _20002;
  wire _20004 = uncoded_block[185] ^ uncoded_block[187];
  wire _20005 = _86 ^ _20004;
  wire _20006 = _4773 ^ _6798;
  wire _20007 = _20005 ^ _20006;
  wire _20008 = _20003 ^ _20007;
  wire _20009 = _20001 ^ _20008;
  wire _20010 = _7411 ^ _4068;
  wire _20011 = _20010 ^ _11406;
  wire _20012 = _19549 ^ _3296;
  wire _20013 = uncoded_block[218] ^ uncoded_block[221];
  wire _20014 = _20013 ^ _7419;
  wire _20015 = _20012 ^ _20014;
  wire _20016 = _20011 ^ _20015;
  wire _20017 = _8028 ^ _968;
  wire _20018 = _2552 ^ _1780;
  wire _20019 = _20017 ^ _20018;
  wire _20020 = uncoded_block[243] ^ uncoded_block[247];
  wire _20021 = uncoded_block[248] ^ uncoded_block[252];
  wire _20022 = _20020 ^ _20021;
  wire _20023 = uncoded_block[255] ^ uncoded_block[259];
  wire _20024 = _20023 ^ _7438;
  wire _20025 = _20022 ^ _20024;
  wire _20026 = _20019 ^ _20025;
  wire _20027 = _20016 ^ _20026;
  wire _20028 = _20009 ^ _20027;
  wire _20029 = _19994 ^ _20028;
  wire _20030 = uncoded_block[270] ^ uncoded_block[276];
  wire _20031 = _985 ^ _20030;
  wire _20032 = _5509 ^ _20031;
  wire _20033 = _4814 ^ _5515;
  wire _20034 = _11424 ^ _991;
  wire _20035 = _20033 ^ _20034;
  wire _20036 = _20032 ^ _20035;
  wire _20037 = _992 ^ _2571;
  wire _20038 = uncoded_block[294] ^ uncoded_block[296];
  wire _20039 = _20038 ^ _8636;
  wire _20040 = _20037 ^ _20039;
  wire _20041 = _7453 ^ _8055;
  wire _20042 = _4115 ^ _145;
  wire _20043 = _20041 ^ _20042;
  wire _20044 = _20040 ^ _20043;
  wire _20045 = _20036 ^ _20044;
  wire _20046 = uncoded_block[324] ^ uncoded_block[329];
  wire _20047 = _20046 ^ _4125;
  wire _20048 = _3352 ^ _13629;
  wire _20049 = _20047 ^ _20048;
  wire _20050 = uncoded_block[346] ^ uncoded_block[350];
  wire _20051 = _20050 ^ _1024;
  wire _20052 = _13631 ^ _20051;
  wire _20053 = _20049 ^ _20052;
  wire _20054 = _6864 ^ _18158;
  wire _20055 = _20054 ^ _19094;
  wire _20056 = uncoded_block[377] ^ uncoded_block[379];
  wire _20057 = _4141 ^ _20056;
  wire _20058 = _1841 ^ _6876;
  wire _20059 = _20057 ^ _20058;
  wire _20060 = _20055 ^ _20059;
  wire _20061 = _20053 ^ _20060;
  wire _20062 = _20045 ^ _20061;
  wire _20063 = _9255 ^ _6239;
  wire _20064 = _10908 ^ _2622;
  wire _20065 = _20063 ^ _20064;
  wire _20066 = _17668 ^ _6244;
  wire _20067 = _184 ^ _1052;
  wire _20068 = _20066 ^ _20067;
  wire _20069 = _20065 ^ _20068;
  wire _20070 = _18172 ^ _13113;
  wire _20071 = uncoded_block[431] ^ uncoded_block[434];
  wire _20072 = _9816 ^ _20071;
  wire _20073 = _201 ^ _5577;
  wire _20074 = _20072 ^ _20073;
  wire _20075 = _20070 ^ _20074;
  wire _20076 = _20069 ^ _20075;
  wire _20077 = _206 ^ _16191;
  wire _20078 = uncoded_block[456] ^ uncoded_block[460];
  wire _20079 = _2650 ^ _20078;
  wire _20080 = _20077 ^ _20079;
  wire _20081 = _13662 ^ _4186;
  wire _20082 = _20081 ^ _1084;
  wire _20083 = _20080 ^ _20082;
  wire _20084 = uncoded_block[481] ^ uncoded_block[486];
  wire _20085 = _15719 ^ _20084;
  wire _20086 = _12578 ^ _2667;
  wire _20087 = _20085 ^ _20086;
  wire _20088 = uncoded_block[504] ^ uncoded_block[508];
  wire _20089 = _2668 ^ _20088;
  wire _20090 = _9295 ^ _13676;
  wire _20091 = _20089 ^ _20090;
  wire _20092 = _20087 ^ _20091;
  wire _20093 = _20083 ^ _20092;
  wire _20094 = _20076 ^ _20093;
  wire _20095 = _20062 ^ _20094;
  wire _20096 = _20029 ^ _20095;
  wire _20097 = uncoded_block[520] ^ uncoded_block[523];
  wire _20098 = _1895 ^ _20097;
  wire _20099 = uncoded_block[524] ^ uncoded_block[526];
  wire _20100 = _20099 ^ _3447;
  wire _20101 = _20098 ^ _20100;
  wire _20102 = _16215 ^ _14197;
  wire _20103 = _9854 ^ _1117;
  wire _20104 = _20102 ^ _20103;
  wire _20105 = _20101 ^ _20104;
  wire _20106 = _6300 ^ _247;
  wire _20107 = uncoded_block[552] ^ uncoded_block[556];
  wire _20108 = _20107 ^ _3461;
  wire _20109 = _20106 ^ _20108;
  wire _20110 = uncoded_block[564] ^ uncoded_block[567];
  wire _20111 = _20110 ^ _14208;
  wire _20112 = _4941 ^ _17718;
  wire _20113 = _20111 ^ _20112;
  wire _20114 = _20109 ^ _20113;
  wire _20115 = _20105 ^ _20114;
  wire _20116 = uncoded_block[586] ^ uncoded_block[588];
  wire _20117 = _1933 ^ _20116;
  wire _20118 = _1141 ^ _2701;
  wire _20119 = _20117 ^ _20118;
  wire _20120 = _14737 ^ _6954;
  wire _20121 = _6323 ^ _8154;
  wire _20122 = _20120 ^ _20121;
  wire _20123 = _20119 ^ _20122;
  wire _20124 = _7563 ^ _7567;
  wire _20125 = uncoded_block[619] ^ uncoded_block[621];
  wire _20126 = uncoded_block[623] ^ uncoded_block[626];
  wire _20127 = _20125 ^ _20126;
  wire _20128 = _20124 ^ _20127;
  wire _20129 = _7576 ^ _16740;
  wire _20130 = _20129 ^ _19673;
  wire _20131 = _20128 ^ _20130;
  wire _20132 = _20123 ^ _20131;
  wire _20133 = _20115 ^ _20132;
  wire _20134 = uncoded_block[651] ^ uncoded_block[656];
  wire _20135 = _20134 ^ _4261;
  wire _20136 = _6344 ^ _1174;
  wire _20137 = _20135 ^ _20136;
  wire _20138 = _8176 ^ _1968;
  wire _20139 = _6353 ^ _13194;
  wire _20140 = _20138 ^ _20139;
  wire _20141 = _20137 ^ _20140;
  wire _20142 = _6357 ^ _328;
  wire _20143 = uncoded_block[699] ^ uncoded_block[703];
  wire _20144 = _19195 ^ _20143;
  wire _20145 = _20142 ^ _20144;
  wire _20146 = _1191 ^ _11004;
  wire _20147 = _340 ^ _9369;
  wire _20148 = _20146 ^ _20147;
  wire _20149 = _20145 ^ _20148;
  wire _20150 = _20141 ^ _20149;
  wire _20151 = uncoded_block[723] ^ uncoded_block[726];
  wire _20152 = _20151 ^ _13749;
  wire _20153 = uncoded_block[734] ^ uncoded_block[737];
  wire _20154 = _1991 ^ _20153;
  wire _20155 = _20152 ^ _20154;
  wire _20156 = uncoded_block[739] ^ uncoded_block[742];
  wire _20157 = _20156 ^ _11576;
  wire _20158 = _2775 ^ _5704;
  wire _20159 = _20157 ^ _20158;
  wire _20160 = _20155 ^ _20159;
  wire _20161 = _2002 ^ _2778;
  wire _20162 = _359 ^ _8781;
  wire _20163 = _20161 ^ _20162;
  wire _20164 = _364 ^ _2784;
  wire _20165 = uncoded_block[775] ^ uncoded_block[777];
  wire _20166 = _20165 ^ _7021;
  wire _20167 = _20164 ^ _20166;
  wire _20168 = _20163 ^ _20167;
  wire _20169 = _20160 ^ _20168;
  wire _20170 = _20150 ^ _20169;
  wire _20171 = _20133 ^ _20170;
  wire _20172 = _2794 ^ _371;
  wire _20173 = _12675 ^ _8791;
  wire _20174 = _20172 ^ _20173;
  wire _20175 = _4317 ^ _3577;
  wire _20176 = _15807 ^ _20175;
  wire _20177 = _20174 ^ _20176;
  wire _20178 = _12127 ^ _5041;
  wire _20179 = _5729 ^ _6398;
  wire _20180 = _20178 ^ _20179;
  wire _20181 = _7037 ^ _11034;
  wire _20182 = _12135 ^ _12686;
  wire _20183 = _20181 ^ _20182;
  wire _20184 = _20180 ^ _20183;
  wire _20185 = _20177 ^ _20184;
  wire _20186 = uncoded_block[839] ^ uncoded_block[842];
  wire _20187 = _2814 ^ _20186;
  wire _20188 = uncoded_block[844] ^ uncoded_block[848];
  wire _20189 = _20188 ^ _7643;
  wire _20190 = _20187 ^ _20189;
  wire _20191 = _8237 ^ _14300;
  wire _20192 = _3603 ^ _413;
  wire _20193 = _20191 ^ _20192;
  wire _20194 = _20190 ^ _20193;
  wire _20195 = _414 ^ _2828;
  wire _20196 = _20195 ^ _7061;
  wire _20197 = _8820 ^ _11059;
  wire _20198 = _13799 ^ _1277;
  wire _20199 = _20197 ^ _20198;
  wire _20200 = _20196 ^ _20199;
  wire _20201 = _20194 ^ _20200;
  wire _20202 = _20185 ^ _20201;
  wire _20203 = _5758 ^ _7066;
  wire _20204 = _8254 ^ _7070;
  wire _20205 = _20203 ^ _20204;
  wire _20206 = uncoded_block[912] ^ uncoded_block[916];
  wire _20207 = _6428 ^ _20206;
  wire _20208 = _17820 ^ _6435;
  wire _20209 = _20207 ^ _20208;
  wire _20210 = _20205 ^ _20209;
  wire _20211 = uncoded_block[933] ^ uncoded_block[939];
  wire _20212 = _448 ^ _20211;
  wire _20213 = _20212 ^ _457;
  wire _20214 = _14326 ^ _16326;
  wire _20215 = _9438 ^ _2093;
  wire _20216 = _20214 ^ _20215;
  wire _20217 = _20213 ^ _20216;
  wire _20218 = _20210 ^ _20217;
  wire _20219 = uncoded_block[972] ^ uncoded_block[976];
  wire _20220 = _1314 ^ _20219;
  wire _20221 = uncoded_block[982] ^ uncoded_block[988];
  wire _20222 = _471 ^ _20221;
  wire _20223 = _20220 ^ _20222;
  wire _20224 = _16338 ^ _479;
  wire _20225 = _480 ^ _3666;
  wire _20226 = _20224 ^ _20225;
  wire _20227 = _20223 ^ _20226;
  wire _20228 = _13283 ^ _2117;
  wire _20229 = _11663 ^ _1334;
  wire _20230 = _20228 ^ _20229;
  wire _20231 = _8301 ^ _18801;
  wire _20232 = _2898 ^ _499;
  wire _20233 = _20231 ^ _20232;
  wire _20234 = _20230 ^ _20233;
  wire _20235 = _20227 ^ _20234;
  wire _20236 = _20218 ^ _20235;
  wire _20237 = _20202 ^ _20236;
  wire _20238 = _20171 ^ _20237;
  wire _20239 = _20096 ^ _20238;
  wire _20240 = _7707 ^ _5810;
  wire _20241 = _6478 ^ _2133;
  wire _20242 = _20240 ^ _20241;
  wire _20243 = _515 ^ _13844;
  wire _20244 = _13846 ^ _1363;
  wire _20245 = _20243 ^ _20244;
  wire _20246 = _20242 ^ _20245;
  wire _20247 = uncoded_block[1062] ^ uncoded_block[1065];
  wire _20248 = _20247 ^ _3689;
  wire _20249 = _15396 ^ _529;
  wire _20250 = _20248 ^ _20249;
  wire _20251 = uncoded_block[1078] ^ uncoded_block[1080];
  wire _20252 = _20251 ^ _7724;
  wire _20253 = uncoded_block[1087] ^ uncoded_block[1090];
  wire _20254 = _2928 ^ _20253;
  wire _20255 = _20252 ^ _20254;
  wire _20256 = _20250 ^ _20255;
  wire _20257 = _20246 ^ _20256;
  wire _20258 = _11689 ^ _8910;
  wire _20259 = _20258 ^ _2162;
  wire _20260 = _8915 ^ _7132;
  wire _20261 = _8917 ^ _19313;
  wire _20262 = _20260 ^ _20261;
  wire _20263 = _20259 ^ _20262;
  wire _20264 = _9489 ^ _4459;
  wire _20265 = uncoded_block[1128] ^ uncoded_block[1131];
  wire _20266 = uncoded_block[1136] ^ uncoded_block[1138];
  wire _20267 = _20265 ^ _20266;
  wire _20268 = _20264 ^ _20267;
  wire _20269 = uncoded_block[1139] ^ uncoded_block[1143];
  wire _20270 = _20269 ^ _2953;
  wire _20271 = _1401 ^ _4466;
  wire _20272 = _20270 ^ _20271;
  wire _20273 = _20268 ^ _20272;
  wire _20274 = _20263 ^ _20273;
  wire _20275 = _20257 ^ _20274;
  wire _20276 = _4468 ^ _8354;
  wire _20277 = _20276 ^ _16892;
  wire _20278 = _1407 ^ _2189;
  wire _20279 = _11161 ^ _2192;
  wire _20280 = _20278 ^ _20279;
  wire _20281 = _20277 ^ _20280;
  wire _20282 = _1411 ^ _6520;
  wire _20283 = _12808 ^ _7756;
  wire _20284 = _20282 ^ _20283;
  wire _20285 = _6525 ^ _11721;
  wire _20286 = uncoded_block[1202] ^ uncoded_block[1206];
  wire _20287 = _7162 ^ _20286;
  wire _20288 = _20285 ^ _20287;
  wire _20289 = _20284 ^ _20288;
  wire _20290 = _20281 ^ _20289;
  wire _20291 = _1427 ^ _10059;
  wire _20292 = uncoded_block[1222] ^ uncoded_block[1228];
  wire _20293 = _20292 ^ _1439;
  wire _20294 = _20291 ^ _20293;
  wire _20295 = _2225 ^ _2989;
  wire _20296 = _15441 ^ _4509;
  wire _20297 = _20295 ^ _20296;
  wire _20298 = _20294 ^ _20297;
  wire _20299 = uncoded_block[1246] ^ uncoded_block[1251];
  wire _20300 = _11734 ^ _20299;
  wire _20301 = _5231 ^ _15934;
  wire _20302 = _20300 ^ _20301;
  wire _20303 = uncoded_block[1269] ^ uncoded_block[1274];
  wire _20304 = _3008 ^ _20303;
  wire _20305 = _3005 ^ _20304;
  wire _20306 = _20302 ^ _20305;
  wire _20307 = _20298 ^ _20306;
  wire _20308 = _20290 ^ _20307;
  wire _20309 = _20275 ^ _20308;
  wire _20310 = uncoded_block[1280] ^ uncoded_block[1287];
  wire _20311 = _5908 ^ _20310;
  wire _20312 = _20311 ^ _7187;
  wire _20313 = _7193 ^ _16424;
  wire _20314 = uncoded_block[1311] ^ uncoded_block[1313];
  wire _20315 = _3025 ^ _20314;
  wire _20316 = _20313 ^ _20315;
  wire _20317 = _20312 ^ _20316;
  wire _20318 = _3811 ^ _4540;
  wire _20319 = _5254 ^ _4543;
  wire _20320 = _20318 ^ _20319;
  wire _20321 = uncoded_block[1325] ^ uncoded_block[1330];
  wire _20322 = _20321 ^ _8998;
  wire _20323 = _4551 ^ _3822;
  wire _20324 = _20322 ^ _20323;
  wire _20325 = _20320 ^ _20324;
  wire _20326 = _20317 ^ _20325;
  wire _20327 = uncoded_block[1346] ^ uncoded_block[1351];
  wire _20328 = _10092 ^ _20327;
  wire _20329 = uncoded_block[1356] ^ uncoded_block[1362];
  wire _20330 = _5272 ^ _20329;
  wire _20331 = _20328 ^ _20330;
  wire _20332 = uncoded_block[1363] ^ uncoded_block[1370];
  wire _20333 = _20332 ^ _8423;
  wire _20334 = uncoded_block[1377] ^ uncoded_block[1379];
  wire _20335 = _3054 ^ _20334;
  wire _20336 = _20333 ^ _20335;
  wire _20337 = _20331 ^ _20336;
  wire _20338 = _7222 ^ _691;
  wire _20339 = _3836 ^ _20338;
  wire _20340 = uncoded_block[1393] ^ uncoded_block[1396];
  wire _20341 = _20340 ^ _5955;
  wire _20342 = _2297 ^ _10678;
  wire _20343 = _20341 ^ _20342;
  wire _20344 = _20339 ^ _20343;
  wire _20345 = _20337 ^ _20344;
  wire _20346 = _20326 ^ _20345;
  wire _20347 = uncoded_block[1413] ^ uncoded_block[1414];
  wire _20348 = _8436 ^ _20347;
  wire _20349 = _2306 ^ _10120;
  wire _20350 = _20348 ^ _20349;
  wire _20351 = _9588 ^ _13429;
  wire _20352 = _1530 ^ _9591;
  wire _20353 = _20351 ^ _20352;
  wire _20354 = _20350 ^ _20353;
  wire _20355 = uncoded_block[1439] ^ uncoded_block[1443];
  wire _20356 = _2314 ^ _20355;
  wire _20357 = uncoded_block[1444] ^ uncoded_block[1446];
  wire _20358 = _20357 ^ _3864;
  wire _20359 = _20356 ^ _20358;
  wire _20360 = _1544 ^ _9037;
  wire _20361 = uncoded_block[1461] ^ uncoded_block[1463];
  wire _20362 = uncoded_block[1464] ^ uncoded_block[1468];
  wire _20363 = _20361 ^ _20362;
  wire _20364 = _20360 ^ _20363;
  wire _20365 = _20359 ^ _20364;
  wire _20366 = _20354 ^ _20365;
  wire _20367 = uncoded_block[1469] ^ uncoded_block[1473];
  wire _20368 = _20367 ^ _4604;
  wire _20369 = uncoded_block[1481] ^ uncoded_block[1485];
  wire _20370 = _3884 ^ _20369;
  wire _20371 = _20368 ^ _20370;
  wire _20372 = _8462 ^ _5993;
  wire _20373 = _741 ^ _20372;
  wire _20374 = _20371 ^ _20373;
  wire _20375 = _1572 ^ _4616;
  wire _20376 = _15002 ^ _7264;
  wire _20377 = _20375 ^ _20376;
  wire _20378 = _7265 ^ _12352;
  wire _20379 = _20378 ^ _16492;
  wire _20380 = _20377 ^ _20379;
  wire _20381 = _20374 ^ _20380;
  wire _20382 = _20366 ^ _20381;
  wire _20383 = _20346 ^ _20382;
  wire _20384 = _20309 ^ _20383;
  wire _20385 = _4624 ^ _6648;
  wire _20386 = uncoded_block[1537] ^ uncoded_block[1541];
  wire _20387 = uncoded_block[1542] ^ uncoded_block[1544];
  wire _20388 = _20386 ^ _20387;
  wire _20389 = _20385 ^ _20388;
  wire _20390 = uncoded_block[1552] ^ uncoded_block[1558];
  wire _20391 = _2367 ^ _20390;
  wire _20392 = uncoded_block[1565] ^ uncoded_block[1566];
  wire _20393 = _2372 ^ _20392;
  wire _20394 = _20391 ^ _20393;
  wire _20395 = _20389 ^ _20394;
  wire _20396 = _16020 ^ _1608;
  wire _20397 = uncoded_block[1579] ^ uncoded_block[1582];
  wire _20398 = _6663 ^ _20397;
  wire _20399 = _20396 ^ _20398;
  wire _20400 = _3925 ^ _3927;
  wire _20401 = uncoded_block[1590] ^ uncoded_block[1592];
  wire _20402 = _20401 ^ _6673;
  wire _20403 = _20400 ^ _20402;
  wire _20404 = _20399 ^ _20403;
  wire _20405 = _20395 ^ _20404;
  wire _20406 = uncoded_block[1603] ^ uncoded_block[1605];
  wire _20407 = _20406 ^ _4662;
  wire _20408 = _12938 ^ _20407;
  wire _20409 = uncoded_block[1612] ^ uncoded_block[1616];
  wire _20410 = _20409 ^ _804;
  wire _20411 = _9095 ^ _3941;
  wire _20412 = _20410 ^ _20411;
  wire _20413 = _20408 ^ _20412;
  wire _20414 = _4665 ^ _4668;
  wire _20415 = _18516 ^ _3172;
  wire _20416 = _20414 ^ _20415;
  wire _20417 = uncoded_block[1652] ^ uncoded_block[1655];
  wire _20418 = _20417 ^ _12390;
  wire _20419 = _12394 ^ _3179;
  wire _20420 = _20418 ^ _20419;
  wire _20421 = _20416 ^ _20420;
  wire _20422 = _20413 ^ _20421;
  wire _20423 = _20405 ^ _20422;
  wire _20424 = _2422 ^ _8521;
  wire _20425 = _7323 ^ _3962;
  wire _20426 = _20424 ^ _20425;
  wire _20427 = uncoded_block[1679] ^ uncoded_block[1680];
  wire _20428 = _20427 ^ _4691;
  wire _20429 = uncoded_block[1686] ^ uncoded_block[1689];
  wire _20430 = _4693 ^ _20429;
  wire _20431 = _20428 ^ _20430;
  wire _20432 = _20426 ^ _20431;
  wire _20433 = _7331 ^ _9675;
  wire _20434 = _10771 ^ _11327;
  wire _20435 = _20433 ^ _20434;
  wire _20436 = uncoded_block[1700] ^ uncoded_block[1702];
  wire _20437 = uncoded_block[1704] ^ uncoded_block[1707];
  wire _20438 = _20436 ^ _20437;
  wire _20439 = _11879 ^ _854;
  wire _20440 = _20438 ^ _20439;
  wire _20441 = _20435 ^ _20440;
  wire _20442 = _20432 ^ _20441;
  wire _20443 = _20442 ^ _3989;
  wire _20444 = _20423 ^ _20443;
  wire _20445 = _20384 ^ _20444;
  wire _20446 = _20239 ^ _20445;
  wire _20447 = _3209 ^ _2453;
  wire _20448 = _20447 ^ _7349;
  wire _20449 = _3216 ^ _871;
  wire _20450 = _10226 ^ _1690;
  wire _20451 = _20449 ^ _20450;
  wire _20452 = _20448 ^ _20451;
  wire _20453 = uncoded_block[22] ^ uncoded_block[25];
  wire _20454 = _20453 ^ _11344;
  wire _20455 = _11890 ^ _879;
  wire _20456 = _20454 ^ _20455;
  wire _20457 = uncoded_block[41] ^ uncoded_block[43];
  wire _20458 = _2466 ^ _20457;
  wire _20459 = uncoded_block[44] ^ uncoded_block[46];
  wire _20460 = _20459 ^ _3232;
  wire _20461 = _20458 ^ _20460;
  wire _20462 = _20456 ^ _20461;
  wire _20463 = _20452 ^ _20462;
  wire _20464 = _3233 ^ _12429;
  wire _20465 = uncoded_block[59] ^ uncoded_block[61];
  wire _20466 = _1703 ^ _20465;
  wire _20467 = _20464 ^ _20466;
  wire _20468 = _9156 ^ _4017;
  wire _20469 = _900 ^ _6749;
  wire _20470 = _20468 ^ _20469;
  wire _20471 = _20467 ^ _20470;
  wire _20472 = uncoded_block[83] ^ uncoded_block[87];
  wire _20473 = _20472 ^ _15603;
  wire _20474 = uncoded_block[91] ^ uncoded_block[98];
  wire _20475 = _20474 ^ _15097;
  wire _20476 = _20473 ^ _20475;
  wire _20477 = _7986 ^ _50;
  wire _20478 = _6126 ^ _1727;
  wire _20479 = _20477 ^ _20478;
  wire _20480 = _20476 ^ _20479;
  wire _20481 = _20471 ^ _20480;
  wire _20482 = _20463 ^ _20481;
  wire _20483 = _2501 ^ _1730;
  wire _20484 = uncoded_block[133] ^ uncoded_block[140];
  wire _20485 = _4754 ^ _20484;
  wire _20486 = _20483 ^ _20485;
  wire _20487 = _16600 ^ _67;
  wire _20488 = uncoded_block[153] ^ uncoded_block[156];
  wire _20489 = _1745 ^ _20488;
  wire _20490 = _20487 ^ _20489;
  wire _20491 = _20486 ^ _20490;
  wire _20492 = _9188 ^ _8589;
  wire _20493 = _6788 ^ _8591;
  wire _20494 = _20492 ^ _20493;
  wire _20495 = _6149 ^ _940;
  wire _20496 = _11935 ^ _7409;
  wire _20497 = _20495 ^ _20496;
  wire _20498 = _20494 ^ _20497;
  wire _20499 = _20491 ^ _20498;
  wire _20500 = uncoded_block[192] ^ uncoded_block[195];
  wire _20501 = _20500 ^ _16116;
  wire _20502 = uncoded_block[203] ^ uncoded_block[207];
  wire _20503 = _8018 ^ _20502;
  wire _20504 = _20501 ^ _20503;
  wire _20505 = _5489 ^ _4787;
  wire _20506 = _5492 ^ _4076;
  wire _20507 = _20505 ^ _20506;
  wire _20508 = _20504 ^ _20507;
  wire _20509 = _3299 ^ _4791;
  wire _20510 = _968 ^ _3305;
  wire _20511 = _20509 ^ _20510;
  wire _20512 = _10292 ^ _6179;
  wire _20513 = _9212 ^ _4800;
  wire _20514 = _20512 ^ _20513;
  wire _20515 = _20511 ^ _20514;
  wire _20516 = _20508 ^ _20515;
  wire _20517 = _20499 ^ _20516;
  wire _20518 = _20482 ^ _20517;
  wire _20519 = _15656 ^ _14639;
  wire _20520 = uncoded_block[260] ^ uncoded_block[262];
  wire _20521 = _20520 ^ _6187;
  wire _20522 = _20519 ^ _20521;
  wire _20523 = uncoded_block[265] ^ uncoded_block[267];
  wire _20524 = _20523 ^ _985;
  wire _20525 = _20524 ^ _3322;
  wire _20526 = _20522 ^ _20525;
  wire _20527 = uncoded_block[278] ^ uncoded_block[280];
  wire _20528 = _1795 ^ _20527;
  wire _20529 = _11967 ^ _4105;
  wire _20530 = _20528 ^ _20529;
  wire _20531 = _5522 ^ _2571;
  wire _20532 = _20531 ^ _8050;
  wire _20533 = _20530 ^ _20532;
  wire _20534 = _20526 ^ _20533;
  wire _20535 = _8636 ^ _142;
  wire _20536 = uncoded_block[306] ^ uncoded_block[310];
  wire _20537 = _8052 ^ _20536;
  wire _20538 = _20535 ^ _20537;
  wire _20539 = uncoded_block[315] ^ uncoded_block[318];
  wire _20540 = _16648 ^ _20539;
  wire _20541 = _4832 ^ _6852;
  wire _20542 = _20540 ^ _20541;
  wire _20543 = _20538 ^ _20542;
  wire _20544 = _4126 ^ _2592;
  wire _20545 = _16153 ^ _20544;
  wire _20546 = uncoded_block[338] ^ uncoded_block[342];
  wire _20547 = uncoded_block[343] ^ uncoded_block[346];
  wire _20548 = _20546 ^ _20547;
  wire _20549 = _20548 ^ _18155;
  wire _20550 = _20545 ^ _20549;
  wire _20551 = _20543 ^ _20550;
  wire _20552 = _20534 ^ _20551;
  wire _20553 = _162 ^ _2601;
  wire _20554 = uncoded_block[356] ^ uncoded_block[358];
  wire _20555 = uncoded_block[359] ^ uncoded_block[366];
  wire _20556 = _20554 ^ _20555;
  wire _20557 = _20553 ^ _20556;
  wire _20558 = _3369 ^ _6873;
  wire _20559 = _4141 ^ _4854;
  wire _20560 = _20558 ^ _20559;
  wire _20561 = _20557 ^ _20560;
  wire _20562 = _1842 ^ _1045;
  wire _20563 = _4152 ^ _10910;
  wire _20564 = _20562 ^ _20563;
  wire _20565 = _2625 ^ _6244;
  wire _20566 = _1049 ^ _20565;
  wire _20567 = _20564 ^ _20566;
  wire _20568 = _20561 ^ _20567;
  wire _20569 = uncoded_block[407] ^ uncoded_block[413];
  wire _20570 = _20569 ^ _4871;
  wire _20571 = _20570 ^ _16678;
  wire _20572 = uncoded_block[428] ^ uncoded_block[434];
  wire _20573 = _20572 ^ _5574;
  wire _20574 = uncoded_block[447] ^ uncoded_block[454];
  wire _20575 = _12559 ^ _20574;
  wire _20576 = _20573 ^ _20575;
  wire _20577 = _20571 ^ _20576;
  wire _20578 = _212 ^ _8681;
  wire _20579 = _13662 ^ _7507;
  wire _20580 = _20578 ^ _20579;
  wire _20581 = _13665 ^ _19625;
  wire _20582 = _20581 ^ _17195;
  wire _20583 = _20580 ^ _20582;
  wire _20584 = _20577 ^ _20583;
  wire _20585 = _20568 ^ _20584;
  wire _20586 = _20552 ^ _20585;
  wire _20587 = _20518 ^ _20586;
  wire _20588 = uncoded_block[484] ^ uncoded_block[487];
  wire _20589 = _20588 ^ _9832;
  wire _20590 = _2664 ^ _5604;
  wire _20591 = _20589 ^ _20590;
  wire _20592 = uncoded_block[499] ^ uncoded_block[502];
  wire _20593 = _20592 ^ _1887;
  wire _20594 = uncoded_block[509] ^ uncoded_block[514];
  wire _20595 = _5611 ^ _20594;
  wire _20596 = _20593 ^ _20595;
  wire _20597 = _20591 ^ _20596;
  wire _20598 = uncoded_block[517] ^ uncoded_block[518];
  wire _20599 = _8706 ^ _20598;
  wire _20600 = _9841 ^ _13684;
  wire _20601 = _20599 ^ _20600;
  wire _20602 = uncoded_block[526] ^ uncoded_block[528];
  wire _20603 = uncoded_block[530] ^ uncoded_block[532];
  wire _20604 = _20602 ^ _20603;
  wire _20605 = _16215 ^ _6932;
  wire _20606 = _20604 ^ _20605;
  wire _20607 = _20601 ^ _20606;
  wire _20608 = _20597 ^ _20607;
  wire _20609 = _5620 ^ _1117;
  wire _20610 = _2688 ^ _8721;
  wire _20611 = _20609 ^ _20610;
  wire _20612 = _1916 ^ _1924;
  wire _20613 = _20612 ^ _14729;
  wire _20614 = _20611 ^ _20613;
  wire _20615 = uncoded_block[569] ^ uncoded_block[573];
  wire _20616 = _20615 ^ _263;
  wire _20617 = _20616 ^ _267;
  wire _20618 = uncoded_block[591] ^ uncoded_block[593];
  wire _20619 = _9864 ^ _20618;
  wire _20620 = _15247 ^ _4952;
  wire _20621 = _20619 ^ _20620;
  wire _20622 = _20617 ^ _20621;
  wire _20623 = _20614 ^ _20622;
  wire _20624 = _20608 ^ _20623;
  wire _20625 = _3487 ^ _2710;
  wire _20626 = uncoded_block[608] ^ uncoded_block[611];
  wire _20627 = uncoded_block[612] ^ uncoded_block[616];
  wire _20628 = _20626 ^ _20627;
  wire _20629 = _20625 ^ _20628;
  wire _20630 = uncoded_block[619] ^ uncoded_block[622];
  wire _20631 = _6959 ^ _20630;
  wire _20632 = _12618 ^ _4247;
  wire _20633 = _20631 ^ _20632;
  wire _20634 = _20629 ^ _20633;
  wire _20635 = _14745 ^ _4249;
  wire _20636 = _20635 ^ _13723;
  wire _20637 = _15766 ^ _301;
  wire _20638 = uncoded_block[659] ^ uncoded_block[662];
  wire _20639 = _3508 ^ _20638;
  wire _20640 = _20637 ^ _20639;
  wire _20641 = _20636 ^ _20640;
  wire _20642 = _20634 ^ _20641;
  wire _20643 = uncoded_block[666] ^ uncoded_block[671];
  wire _20644 = _308 ^ _20643;
  wire _20645 = _1178 ^ _10434;
  wire _20646 = _20644 ^ _20645;
  wire _20647 = _6352 ^ _3522;
  wire _20648 = uncoded_block[685] ^ uncoded_block[690];
  wire _20649 = _3526 ^ _20648;
  wire _20650 = _20647 ^ _20649;
  wire _20651 = _20646 ^ _20650;
  wire _20652 = _6360 ^ _17258;
  wire _20653 = _7591 ^ _20652;
  wire _20654 = uncoded_block[703] ^ uncoded_block[706];
  wire _20655 = _20654 ^ _8190;
  wire _20656 = _1192 ^ _337;
  wire _20657 = _20655 ^ _20656;
  wire _20658 = _20653 ^ _20657;
  wire _20659 = _20651 ^ _20658;
  wire _20660 = _20642 ^ _20659;
  wire _20661 = _20624 ^ _20660;
  wire _20662 = _4999 ^ _340;
  wire _20663 = _8198 ^ _14774;
  wire _20664 = _20662 ^ _20663;
  wire _20665 = _7002 ^ _1203;
  wire _20666 = _5702 ^ _5013;
  wire _20667 = _20665 ^ _20666;
  wire _20668 = _20664 ^ _20667;
  wire _20669 = uncoded_block[752] ^ uncoded_block[757];
  wire _20670 = _1210 ^ _20669;
  wire _20671 = _5019 ^ _14271;
  wire _20672 = _20670 ^ _20671;
  wire _20673 = _5711 ^ _14278;
  wire _20674 = _17284 ^ _2019;
  wire _20675 = _20673 ^ _20674;
  wire _20676 = _20672 ^ _20675;
  wire _20677 = _20668 ^ _20676;
  wire _20678 = _11591 ^ _8224;
  wire _20679 = _3575 ^ _20678;
  wire _20680 = _1235 ^ _5041;
  wire _20681 = _5042 ^ _1241;
  wire _20682 = _20680 ^ _20681;
  wire _20683 = _20679 ^ _20682;
  wire _20684 = _12135 ^ _14807;
  wire _20685 = _4329 ^ _20684;
  wire _20686 = _5054 ^ _20186;
  wire _20687 = _2043 ^ _14814;
  wire _20688 = _20686 ^ _20687;
  wire _20689 = _20685 ^ _20688;
  wire _20690 = _20683 ^ _20689;
  wire _20691 = _20677 ^ _20690;
  wire _20692 = uncoded_block[857] ^ uncoded_block[859];
  wire _20693 = _7049 ^ _20692;
  wire _20694 = _20693 ^ _415;
  wire _20695 = _2828 ^ _6416;
  wire _20696 = uncoded_block[879] ^ uncoded_block[881];
  wire _20697 = _11620 ^ _20696;
  wire _20698 = _20695 ^ _20697;
  wire _20699 = _20694 ^ _20698;
  wire _20700 = _423 ^ _7660;
  wire _20701 = uncoded_block[891] ^ uncoded_block[893];
  wire _20702 = _20701 ^ _5085;
  wire _20703 = _20700 ^ _20702;
  wire _20704 = uncoded_block[897] ^ uncoded_block[900];
  wire _20705 = _20704 ^ _7070;
  wire _20706 = _1287 ^ _438;
  wire _20707 = _20705 ^ _20706;
  wire _20708 = _20703 ^ _20707;
  wire _20709 = _20699 ^ _20708;
  wire _20710 = _439 ^ _446;
  wire _20711 = _1296 ^ _15848;
  wire _20712 = _20710 ^ _20711;
  wire _20713 = _2084 ^ _8271;
  wire _20714 = _456 ^ _3643;
  wire _20715 = _20713 ^ _20714;
  wire _20716 = _20712 ^ _20715;
  wire _20717 = _461 ^ _7680;
  wire _20718 = _20717 ^ _8281;
  wire _20719 = _12180 ^ _1314;
  wire _20720 = _20719 ^ _18326;
  wire _20721 = _20718 ^ _20720;
  wire _20722 = _20716 ^ _20721;
  wire _20723 = _20709 ^ _20722;
  wire _20724 = _20691 ^ _20723;
  wire _20725 = _20661 ^ _20724;
  wire _20726 = _20587 ^ _20725;
  wire _20727 = _10535 ^ _8857;
  wire _20728 = uncoded_block[993] ^ uncoded_block[998];
  wire _20729 = _8859 ^ _20728;
  wire _20730 = uncoded_block[1003] ^ uncoded_block[1005];
  wire _20731 = _2111 ^ _20730;
  wire _20732 = _20729 ^ _20731;
  wire _20733 = _20727 ^ _20732;
  wire _20734 = _487 ^ _2117;
  wire _20735 = _7703 ^ _8871;
  wire _20736 = _20734 ^ _20735;
  wire _20737 = _2120 ^ _9454;
  wire _20738 = _495 ^ _2898;
  wire _20739 = _20737 ^ _20738;
  wire _20740 = _20736 ^ _20739;
  wire _20741 = _20733 ^ _20740;
  wire _20742 = _499 ^ _6474;
  wire _20743 = _20742 ^ _513;
  wire _20744 = uncoded_block[1044] ^ uncoded_block[1047];
  wire _20745 = _20744 ^ _518;
  wire _20746 = _12762 ^ _6483;
  wire _20747 = _20745 ^ _20746;
  wire _20748 = _20743 ^ _20747;
  wire _20749 = _2140 ^ _2921;
  wire _20750 = _1366 ^ _5158;
  wire _20751 = _20749 ^ _20750;
  wire _20752 = _2146 ^ _8895;
  wire _20753 = uncoded_block[1083] ^ uncoded_block[1085];
  wire _20754 = _20753 ^ _19306;
  wire _20755 = _20752 ^ _20754;
  wire _20756 = _20751 ^ _20755;
  wire _20757 = _20748 ^ _20756;
  wire _20758 = _20741 ^ _20757;
  wire _20759 = _11137 ^ _11139;
  wire _20760 = uncoded_block[1100] ^ uncoded_block[1103];
  wire _20761 = uncoded_block[1104] ^ uncoded_block[1109];
  wire _20762 = _20760 ^ _20761;
  wire _20763 = _20759 ^ _20762;
  wire _20764 = _15407 ^ _19313;
  wire _20765 = _2941 ^ _12789;
  wire _20766 = _20764 ^ _20765;
  wire _20767 = _20763 ^ _20766;
  wire _20768 = _14887 ^ _14380;
  wire _20769 = _15895 ^ _20768;
  wire _20770 = _4462 ^ _18377;
  wire _20771 = _10597 ^ _6505;
  wire _20772 = _20770 ^ _20771;
  wire _20773 = _20769 ^ _20772;
  wire _20774 = _20767 ^ _20773;
  wire _20775 = _8354 ^ _3733;
  wire _20776 = uncoded_block[1164] ^ uncoded_block[1169];
  wire _20777 = _20776 ^ _1410;
  wire _20778 = _20775 ^ _20777;
  wire _20779 = _17890 ^ _3742;
  wire _20780 = _1417 ^ _19339;
  wire _20781 = _20779 ^ _20780;
  wire _20782 = _20778 ^ _20781;
  wire _20783 = _7159 ^ _8951;
  wire _20784 = _2206 ^ _7763;
  wire _20785 = _20783 ^ _20784;
  wire _20786 = _2978 ^ _2217;
  wire _20787 = _18395 ^ _2982;
  wire _20788 = _20786 ^ _20787;
  wire _20789 = _20785 ^ _20788;
  wire _20790 = _20782 ^ _20789;
  wire _20791 = _20774 ^ _20790;
  wire _20792 = _20758 ^ _20791;
  wire _20793 = _10620 ^ _5215;
  wire _20794 = _5891 ^ _5218;
  wire _20795 = _20793 ^ _20794;
  wire _20796 = _8962 ^ _18860;
  wire _20797 = _18405 ^ _20796;
  wire _20798 = _20795 ^ _20797;
  wire _20799 = _2235 ^ _3001;
  wire _20800 = _10070 ^ _20799;
  wire _20801 = uncoded_block[1257] ^ uncoded_block[1259];
  wire _20802 = _20801 ^ _1458;
  wire _20803 = _1459 ^ _628;
  wire _20804 = _20802 ^ _20803;
  wire _20805 = _20800 ^ _20804;
  wire _20806 = _20798 ^ _20805;
  wire _20807 = _7791 ^ _631;
  wire _20808 = uncoded_block[1284] ^ uncoded_block[1288];
  wire _20809 = _9541 ^ _20808;
  wire _20810 = _20807 ^ _20809;
  wire _20811 = _4529 ^ _642;
  wire _20812 = uncoded_block[1302] ^ uncoded_block[1305];
  wire _20813 = _645 ^ _20812;
  wire _20814 = _20811 ^ _20813;
  wire _20815 = _20810 ^ _20814;
  wire _20816 = uncoded_block[1312] ^ uncoded_block[1315];
  wire _20817 = _3808 ^ _20816;
  wire _20818 = _5926 ^ _654;
  wire _20819 = _20817 ^ _20818;
  wire _20820 = _3814 ^ _8411;
  wire _20821 = _20820 ^ _6579;
  wire _20822 = _20819 ^ _20821;
  wire _20823 = _20815 ^ _20822;
  wire _20824 = _20806 ^ _20823;
  wire _20825 = _1495 ^ _17938;
  wire _20826 = _11771 ^ _4558;
  wire _20827 = _20825 ^ _20826;
  wire _20828 = _5940 ^ _3045;
  wire _20829 = uncoded_block[1370] ^ uncoded_block[1373];
  wire _20830 = _5281 ^ _20829;
  wire _20831 = _20828 ^ _20830;
  wire _20832 = _20827 ^ _20831;
  wire _20833 = _12305 ^ _20334;
  wire _20834 = uncoded_block[1386] ^ uncoded_block[1393];
  wire _20835 = uncoded_block[1394] ^ uncoded_block[1398];
  wire _20836 = _20834 ^ _20835;
  wire _20837 = _20833 ^ _20836;
  wire _20838 = _1517 ^ _3847;
  wire _20839 = _5294 ^ _17461;
  wire _20840 = _20838 ^ _20839;
  wire _20841 = _20837 ^ _20840;
  wire _20842 = _20832 ^ _20841;
  wire _20843 = _13422 ^ _705;
  wire _20844 = _9021 ^ _3074;
  wire _20845 = _20843 ^ _20844;
  wire _20846 = uncoded_block[1429] ^ uncoded_block[1433];
  wire _20847 = _2308 ^ _20846;
  wire _20848 = _14978 ^ _6613;
  wire _20849 = _20847 ^ _20848;
  wire _20850 = _20845 ^ _20849;
  wire _20851 = _20357 ^ _2325;
  wire _20852 = uncoded_block[1453] ^ uncoded_block[1456];
  wire _20853 = _2326 ^ _20852;
  wire _20854 = _20851 ^ _20853;
  wire _20855 = uncoded_block[1463] ^ uncoded_block[1467];
  wire _20856 = _7241 ^ _20855;
  wire _20857 = _7247 ^ _18470;
  wire _20858 = _20856 ^ _20857;
  wire _20859 = _20854 ^ _20858;
  wire _20860 = _20850 ^ _20859;
  wire _20861 = _20842 ^ _20860;
  wire _20862 = _20824 ^ _20861;
  wire _20863 = _20792 ^ _20862;
  wire _20864 = _2342 ^ _1558;
  wire _20865 = _1559 ^ _16981;
  wire _20866 = _20864 ^ _20865;
  wire _20867 = _4610 ^ _6631;
  wire _20868 = _6634 ^ _3111;
  wire _20869 = _20867 ^ _20868;
  wire _20870 = _20866 ^ _20869;
  wire _20871 = _5334 ^ _3117;
  wire _20872 = _12347 ^ _20871;
  wire _20873 = _2357 ^ _3118;
  wire _20874 = uncoded_block[1526] ^ uncoded_block[1531];
  wire _20875 = _20874 ^ _12914;
  wire _20876 = _20873 ^ _20875;
  wire _20877 = _20872 ^ _20876;
  wire _20878 = _20870 ^ _20877;
  wire _20879 = _12917 ^ _1589;
  wire _20880 = uncoded_block[1545] ^ uncoded_block[1556];
  wire _20881 = _20880 ^ _11281;
  wire _20882 = _20879 ^ _20881;
  wire _20883 = _774 ^ _11284;
  wire _20884 = _7891 ^ _4648;
  wire _20885 = _20883 ^ _20884;
  wire _20886 = _20882 ^ _20885;
  wire _20887 = _4651 ^ _784;
  wire _20888 = _15538 ^ _14512;
  wire _20889 = _20887 ^ _20888;
  wire _20890 = _13996 ^ _1621;
  wire _20891 = _20406 ^ _800;
  wire _20892 = _20890 ^ _20891;
  wire _20893 = _20889 ^ _20892;
  wire _20894 = _20886 ^ _20893;
  wire _20895 = _20878 ^ _20894;
  wire _20896 = _6040 ^ _801;
  wire _20897 = _16032 ^ _9095;
  wire _20898 = _20896 ^ _20897;
  wire _20899 = _7300 ^ _9656;
  wire _20900 = uncoded_block[1632] ^ uncoded_block[1636];
  wire _20901 = uncoded_block[1638] ^ uncoded_block[1641];
  wire _20902 = _20900 ^ _20901;
  wire _20903 = _20899 ^ _20902;
  wire _20904 = _20898 ^ _20903;
  wire _20905 = uncoded_block[1645] ^ uncoded_block[1649];
  wire _20906 = _13500 ^ _20905;
  wire _20907 = _3172 ^ _20417;
  wire _20908 = _20906 ^ _20907;
  wire _20909 = uncoded_block[1658] ^ uncoded_block[1660];
  wire _20910 = _12390 ^ _20909;
  wire _20911 = _2419 ^ _5399;
  wire _20912 = _20910 ^ _20911;
  wire _20913 = _20908 ^ _20912;
  wire _20914 = _20904 ^ _20913;
  wire _20915 = _14537 ^ _17037;
  wire _20916 = _11321 ^ _9669;
  wire _20917 = _20916 ^ _18042;
  wire _20918 = _20915 ^ _20917;
  wire _20919 = _11327 ^ _6068;
  wire _20920 = uncoded_block[1702] ^ uncoded_block[1704];
  wire _20921 = _20920 ^ _848;
  wire _20922 = _20919 ^ _20921;
  wire _20923 = uncoded_block[1717] ^ uncoded_block[1719];
  wire _20924 = _11879 ^ _20923;
  wire _20925 = _20924 ^ uncoded_block[1722];
  wire _20926 = _20922 ^ _20925;
  wire _20927 = _20918 ^ _20926;
  wire _20928 = _20914 ^ _20927;
  wire _20929 = _20895 ^ _20928;
  wire _20930 = _20863 ^ _20929;
  wire _20931 = _20726 ^ _20930;
  wire _20932 = uncoded_block[4] ^ uncoded_block[9];
  wire _20933 = _0 ^ _20932;
  wire _20934 = _15075 ^ _871;
  wire _20935 = _20933 ^ _20934;
  wire _20936 = _13537 ^ _3219;
  wire _20937 = uncoded_block[27] ^ uncoded_block[31];
  wire _20938 = _6089 ^ _20937;
  wire _20939 = _20936 ^ _20938;
  wire _20940 = _20935 ^ _20939;
  wire _20941 = uncoded_block[40] ^ uncoded_block[43];
  wire _20942 = _2462 ^ _20941;
  wire _20943 = _12425 ^ _5435;
  wire _20944 = _20942 ^ _20943;
  wire _20945 = _888 ^ _19974;
  wire _20946 = _2474 ^ _12435;
  wire _20947 = _20945 ^ _20946;
  wire _20948 = _20944 ^ _20947;
  wire _20949 = _20940 ^ _20948;
  wire _20950 = _34 ^ _4020;
  wire _20951 = _20950 ^ _10247;
  wire _20952 = uncoded_block[94] ^ uncoded_block[96];
  wire _20953 = _19515 ^ _20952;
  wire _20954 = _10251 ^ _15101;
  wire _20955 = _20953 ^ _20954;
  wire _20956 = _20951 ^ _20955;
  wire _20957 = uncoded_block[108] ^ uncoded_block[110];
  wire _20958 = _20957 ^ _10816;
  wire _20959 = _16592 ^ _2501;
  wire _20960 = _20958 ^ _20959;
  wire _20961 = uncoded_block[123] ^ uncoded_block[125];
  wire _20962 = _20961 ^ _917;
  wire _20963 = uncoded_block[132] ^ uncoded_block[134];
  wire _20964 = _923 ^ _20963;
  wire _20965 = _20962 ^ _20964;
  wire _20966 = _20960 ^ _20965;
  wire _20967 = _20956 ^ _20966;
  wire _20968 = _20949 ^ _20967;
  wire _20969 = uncoded_block[135] ^ uncoded_block[137];
  wire _20970 = _20969 ^ _4043;
  wire _20971 = _7392 ^ _1744;
  wire _20972 = _20970 ^ _20971;
  wire _20973 = uncoded_block[154] ^ uncoded_block[158];
  wire _20974 = _15623 ^ _20973;
  wire _20975 = uncoded_block[159] ^ uncoded_block[163];
  wire _20976 = _20975 ^ _4054;
  wire _20977 = _20974 ^ _20976;
  wire _20978 = _20972 ^ _20977;
  wire _20979 = uncoded_block[174] ^ uncoded_block[177];
  wire _20980 = _79 ^ _20979;
  wire _20981 = _5477 ^ _86;
  wire _20982 = _20980 ^ _20981;
  wire _20983 = _945 ^ _947;
  wire _20984 = _4776 ^ _7411;
  wire _20985 = _20983 ^ _20984;
  wire _20986 = _20982 ^ _20985;
  wire _20987 = _20978 ^ _20986;
  wire _20988 = _15135 ^ _14099;
  wire _20989 = _20988 ^ _13043;
  wire _20990 = uncoded_block[225] ^ uncoded_block[230];
  wire _20991 = _15644 ^ _20990;
  wire _20992 = _3297 ^ _20991;
  wire _20993 = _20989 ^ _20992;
  wire _20994 = uncoded_block[235] ^ uncoded_block[239];
  wire _20995 = _1775 ^ _20994;
  wire _20996 = _10860 ^ _6179;
  wire _20997 = _20995 ^ _20996;
  wire _20998 = _16626 ^ _11954;
  wire _20999 = uncoded_block[254] ^ uncoded_block[256];
  wire _21000 = _13053 ^ _20999;
  wire _21001 = _20998 ^ _21000;
  wire _21002 = _20997 ^ _21001;
  wire _21003 = _20993 ^ _21002;
  wire _21004 = _20987 ^ _21003;
  wire _21005 = _20968 ^ _21004;
  wire _21006 = _14639 ^ _6185;
  wire _21007 = uncoded_block[266] ^ uncoded_block[270];
  wire _21008 = _6187 ^ _21007;
  wire _21009 = _21006 ^ _21008;
  wire _21010 = _3320 ^ _130;
  wire _21011 = _4103 ^ _11967;
  wire _21012 = _21010 ^ _21011;
  wire _21013 = _21009 ^ _21012;
  wire _21014 = uncoded_block[294] ^ uncoded_block[297];
  wire _21015 = _134 ^ _21014;
  wire _21016 = uncoded_block[298] ^ uncoded_block[304];
  wire _21017 = uncoded_block[308] ^ uncoded_block[309];
  wire _21018 = _21016 ^ _21017;
  wire _21019 = _21015 ^ _21018;
  wire _21020 = _1006 ^ _4832;
  wire _21021 = _2583 ^ _12521;
  wire _21022 = _21020 ^ _21021;
  wire _21023 = _21019 ^ _21022;
  wire _21024 = _21013 ^ _21023;
  wire _21025 = _15172 ^ _5536;
  wire _21026 = _10323 ^ _3355;
  wire _21027 = _21025 ^ _21026;
  wire _21028 = uncoded_block[349] ^ uncoded_block[355];
  wire _21029 = _21028 ^ _2602;
  wire _21030 = uncoded_block[362] ^ uncoded_block[363];
  wire _21031 = _6864 ^ _21030;
  wire _21032 = _21029 ^ _21031;
  wire _21033 = _21027 ^ _21032;
  wire _21034 = _13094 ^ _1038;
  wire _21035 = _8077 ^ _21034;
  wire _21036 = _3380 ^ _18633;
  wire _21037 = _21036 ^ _2624;
  wire _21038 = _21035 ^ _21037;
  wire _21039 = _21033 ^ _21038;
  wire _21040 = _21024 ^ _21039;
  wire _21041 = _12545 ^ _2629;
  wire _21042 = _3394 ^ _9266;
  wire _21043 = _21041 ^ _21042;
  wire _21044 = _4871 ^ _15197;
  wire _21045 = _14160 ^ _1060;
  wire _21046 = _21044 ^ _21045;
  wire _21047 = _21043 ^ _21046;
  wire _21048 = _14163 ^ _9271;
  wire _21049 = uncoded_block[440] ^ uncoded_block[442];
  wire _21050 = _6255 ^ _21049;
  wire _21051 = _21048 ^ _21050;
  wire _21052 = uncoded_block[443] ^ uncoded_block[445];
  wire _21053 = _21052 ^ _4177;
  wire _21054 = _21053 ^ _17684;
  wire _21055 = _21051 ^ _21054;
  wire _21056 = _21047 ^ _21055;
  wire _21057 = uncoded_block[460] ^ uncoded_block[463];
  wire _21058 = _21057 ^ _4890;
  wire _21059 = uncoded_block[466] ^ uncoded_block[470];
  wire _21060 = _21059 ^ _11494;
  wire _21061 = _21058 ^ _21060;
  wire _21062 = _5592 ^ _8110;
  wire _21063 = _15212 ^ _8115;
  wire _21064 = _21062 ^ _21063;
  wire _21065 = _21061 ^ _21064;
  wire _21066 = _10937 ^ _5603;
  wire _21067 = uncoded_block[498] ^ uncoded_block[500];
  wire _21068 = _21067 ^ _6921;
  wire _21069 = _21066 ^ _21068;
  wire _21070 = _19137 ^ _16702;
  wire _21071 = _21069 ^ _21070;
  wire _21072 = _21065 ^ _21071;
  wire _21073 = _21056 ^ _21072;
  wire _21074 = _21040 ^ _21073;
  wire _21075 = _21005 ^ _21074;
  wire _21076 = _20598 ^ _3445;
  wire _21077 = _13684 ^ _12586;
  wire _21078 = _21076 ^ _21077;
  wire _21079 = uncoded_block[538] ^ uncoded_block[540];
  wire _21080 = _21079 ^ _8132;
  wire _21081 = _19147 ^ _21080;
  wire _21082 = _21078 ^ _21081;
  wire _21083 = _244 ^ _246;
  wire _21084 = _247 ^ _8724;
  wire _21085 = _21083 ^ _21084;
  wire _21086 = _6305 ^ _9319;
  wire _21087 = uncoded_block[568] ^ uncoded_block[573];
  wire _21088 = _9320 ^ _21087;
  wire _21089 = _21086 ^ _21088;
  wire _21090 = _21085 ^ _21089;
  wire _21091 = _21082 ^ _21090;
  wire _21092 = _1138 ^ _266;
  wire _21093 = _12058 ^ _21092;
  wire _21094 = uncoded_block[598] ^ uncoded_block[603];
  wire _21095 = _18222 ^ _21094;
  wire _21096 = _21095 ^ _20121;
  wire _21097 = _21093 ^ _21096;
  wire _21098 = uncoded_block[614] ^ uncoded_block[616];
  wire _21099 = _7563 ^ _21098;
  wire _21100 = _6959 ^ _4963;
  wire _21101 = _21099 ^ _21100;
  wire _21102 = _10418 ^ _1154;
  wire _21103 = _1156 ^ _10420;
  wire _21104 = _21102 ^ _21103;
  wire _21105 = _21101 ^ _21104;
  wire _21106 = _21097 ^ _21105;
  wire _21107 = _21091 ^ _21106;
  wire _21108 = _4255 ^ _294;
  wire _21109 = _296 ^ _14234;
  wire _21110 = _21108 ^ _21109;
  wire _21111 = uncoded_block[654] ^ uncoded_block[658];
  wire _21112 = _21111 ^ _4261;
  wire _21113 = uncoded_block[663] ^ uncoded_block[666];
  wire _21114 = _15768 ^ _21113;
  wire _21115 = _21112 ^ _21114;
  wire _21116 = _21110 ^ _21115;
  wire _21117 = _9886 ^ _1178;
  wire _21118 = _8760 ^ _13731;
  wire _21119 = _21117 ^ _21118;
  wire _21120 = _6352 ^ _1972;
  wire _21121 = _325 ^ _11556;
  wire _21122 = _21120 ^ _21121;
  wire _21123 = _21119 ^ _21122;
  wire _21124 = _21116 ^ _21123;
  wire _21125 = _6990 ^ _20143;
  wire _21126 = uncoded_block[714] ^ uncoded_block[720];
  wire _21127 = _11565 ^ _21126;
  wire _21128 = _21125 ^ _21127;
  wire _21129 = uncoded_block[724] ^ uncoded_block[727];
  wire _21130 = _9369 ^ _21129;
  wire _21131 = uncoded_block[730] ^ uncoded_block[735];
  wire _21132 = _7001 ^ _21131;
  wire _21133 = _21130 ^ _21132;
  wire _21134 = _21128 ^ _21133;
  wire _21135 = _350 ^ _1207;
  wire _21136 = uncoded_block[743] ^ uncoded_block[746];
  wire _21137 = _21136 ^ _5013;
  wire _21138 = _21135 ^ _21137;
  wire _21139 = uncoded_block[749] ^ uncoded_block[753];
  wire _21140 = _21139 ^ _11012;
  wire _21141 = _2781 ^ _2784;
  wire _21142 = _21140 ^ _21141;
  wire _21143 = _21138 ^ _21142;
  wire _21144 = _21134 ^ _21143;
  wire _21145 = _21124 ^ _21144;
  wire _21146 = _21107 ^ _21145;
  wire _21147 = _2791 ^ _5711;
  wire _21148 = _21147 ^ _13220;
  wire _21149 = uncoded_block[792] ^ uncoded_block[797];
  wire _21150 = _6388 ^ _21149;
  wire _21151 = _16791 ^ _11596;
  wire _21152 = _21150 ^ _21151;
  wire _21153 = _21148 ^ _21152;
  wire _21154 = _1239 ^ _7634;
  wire _21155 = uncoded_block[821] ^ uncoded_block[824];
  wire _21156 = _21155 ^ _12135;
  wire _21157 = _21154 ^ _21156;
  wire _21158 = _10490 ^ _1250;
  wire _21159 = uncoded_block[838] ^ uncoded_block[842];
  wire _21160 = _12138 ^ _21159;
  wire _21161 = _21158 ^ _21160;
  wire _21162 = _21157 ^ _21161;
  wire _21163 = _21153 ^ _21162;
  wire _21164 = _1256 ^ _405;
  wire _21165 = uncoded_block[851] ^ uncoded_block[855];
  wire _21166 = _21165 ^ _17803;
  wire _21167 = _21164 ^ _21166;
  wire _21168 = _17304 ^ _12696;
  wire _21169 = _417 ^ _16304;
  wire _21170 = _21168 ^ _21169;
  wire _21171 = _21167 ^ _21170;
  wire _21172 = uncoded_block[882] ^ uncoded_block[888];
  wire _21173 = _21172 ^ _4354;
  wire _21174 = _14827 ^ _5758;
  wire _21175 = _21173 ^ _21174;
  wire _21176 = _3617 ^ _2844;
  wire _21177 = _19251 ^ _12708;
  wire _21178 = _21176 ^ _21177;
  wire _21179 = _21175 ^ _21178;
  wire _21180 = _21171 ^ _21179;
  wire _21181 = _21163 ^ _21180;
  wire _21182 = uncoded_block[913] ^ uncoded_block[919];
  wire _21183 = _21182 ^ _15840;
  wire _21184 = _16827 ^ _4371;
  wire _21185 = _21183 ^ _21184;
  wire _21186 = _9431 ^ _7080;
  wire _21187 = uncoded_block[942] ^ uncoded_block[946];
  wire _21188 = _453 ^ _21187;
  wire _21189 = _21186 ^ _21188;
  wire _21190 = _21185 ^ _21189;
  wire _21191 = uncoded_block[949] ^ uncoded_block[951];
  wire _21192 = _9975 ^ _21191;
  wire _21193 = _461 ^ _8277;
  wire _21194 = _21192 ^ _21193;
  wire _21195 = _467 ^ _1315;
  wire _21196 = _8281 ^ _21195;
  wire _21197 = _21194 ^ _21196;
  wire _21198 = _21190 ^ _21197;
  wire _21199 = _5789 ^ _8853;
  wire _21200 = _7689 ^ _11098;
  wire _21201 = _21199 ^ _21200;
  wire _21202 = _12737 ^ _479;
  wire _21203 = _11101 ^ _483;
  wire _21204 = _21202 ^ _21203;
  wire _21205 = _21201 ^ _21204;
  wire _21206 = uncoded_block[1008] ^ uncoded_block[1013];
  wire _21207 = _21206 ^ _2893;
  wire _21208 = _1334 ^ _1338;
  wire _21209 = _21207 ^ _21208;
  wire _21210 = _5806 ^ _501;
  wire _21211 = _8876 ^ _21210;
  wire _21212 = _21209 ^ _21211;
  wire _21213 = _21205 ^ _21212;
  wire _21214 = _21198 ^ _21213;
  wire _21215 = _21181 ^ _21214;
  wire _21216 = _21146 ^ _21215;
  wire _21217 = _21075 ^ _21216;
  wire _21218 = uncoded_block[1036] ^ uncoded_block[1039];
  wire _21219 = _21218 ^ _1346;
  wire _21220 = _2130 ^ _9464;
  wire _21221 = _21219 ^ _21220;
  wire _21222 = _9465 ^ _7117;
  wire _21223 = uncoded_block[1069] ^ uncoded_block[1073];
  wire _21224 = _7717 ^ _21223;
  wire _21225 = _21222 ^ _21224;
  wire _21226 = _21221 ^ _21225;
  wire _21227 = _6486 ^ _5162;
  wire _21228 = uncoded_block[1080] ^ uncoded_block[1084];
  wire _21229 = _21228 ^ _2149;
  wire _21230 = _21227 ^ _21229;
  wire _21231 = _11137 ^ _543;
  wire _21232 = _20760 ^ _8914;
  wire _21233 = _21231 ^ _21232;
  wire _21234 = _21230 ^ _21233;
  wire _21235 = _21226 ^ _21234;
  wire _21236 = _2164 ^ _7132;
  wire _21237 = _12782 ^ _3714;
  wire _21238 = _21236 ^ _21237;
  wire _21239 = _14376 ^ _4459;
  wire _21240 = _20265 ^ _8929;
  wire _21241 = _21239 ^ _21240;
  wire _21242 = _21238 ^ _21241;
  wire _21243 = _4462 ^ _2952;
  wire _21244 = uncoded_block[1146] ^ uncoded_block[1150];
  wire _21245 = _21244 ^ _2185;
  wire _21246 = _21243 ^ _21245;
  wire _21247 = _6510 ^ _2958;
  wire _21248 = uncoded_block[1167] ^ uncoded_block[1170];
  wire _21249 = _21248 ^ _1410;
  wire _21250 = _21247 ^ _21249;
  wire _21251 = _21246 ^ _21250;
  wire _21252 = _21242 ^ _21251;
  wire _21253 = _21235 ^ _21252;
  wire _21254 = _2967 ^ _1411;
  wire _21255 = _4482 ^ _4486;
  wire _21256 = _21254 ^ _21255;
  wire _21257 = uncoded_block[1189] ^ uncoded_block[1193];
  wire _21258 = _5201 ^ _21257;
  wire _21259 = uncoded_block[1195] ^ uncoded_block[1198];
  wire _21260 = _21259 ^ _599;
  wire _21261 = _21258 ^ _21260;
  wire _21262 = _21256 ^ _21261;
  wire _21263 = uncoded_block[1206] ^ uncoded_block[1213];
  wire _21264 = _7163 ^ _21263;
  wire _21265 = _2219 ^ _3763;
  wire _21266 = _21264 ^ _21265;
  wire _21267 = _3765 ^ _13355;
  wire _21268 = _612 ^ _7169;
  wire _21269 = _21267 ^ _21268;
  wire _21270 = _21266 ^ _21269;
  wire _21271 = _21262 ^ _21270;
  wire _21272 = _3771 ^ _616;
  wire _21273 = uncoded_block[1247] ^ uncoded_block[1253];
  wire _21274 = _21273 ^ _2238;
  wire _21275 = _21272 ^ _21274;
  wire _21276 = _3004 ^ _2239;
  wire _21277 = _12832 ^ _4523;
  wire _21278 = _21276 ^ _21277;
  wire _21279 = _21275 ^ _21278;
  wire _21280 = uncoded_block[1277] ^ uncoded_block[1279];
  wire _21281 = _1463 ^ _21280;
  wire _21282 = uncoded_block[1281] ^ uncoded_block[1285];
  wire _21283 = _21282 ^ _18417;
  wire _21284 = _21281 ^ _21283;
  wire _21285 = uncoded_block[1290] ^ uncoded_block[1298];
  wire _21286 = _21285 ^ _1472;
  wire _21287 = _21286 ^ _3809;
  wire _21288 = _21284 ^ _21287;
  wire _21289 = _21279 ^ _21288;
  wire _21290 = _21271 ^ _21289;
  wire _21291 = _21253 ^ _21290;
  wire _21292 = uncoded_block[1312] ^ uncoded_block[1316];
  wire _21293 = uncoded_block[1317] ^ uncoded_block[1318];
  wire _21294 = _21292 ^ _21293;
  wire _21295 = _2265 ^ _19375;
  wire _21296 = _21294 ^ _21295;
  wire _21297 = _16435 ^ _3820;
  wire _21298 = uncoded_block[1339] ^ uncoded_block[1345];
  wire _21299 = _661 ^ _21298;
  wire _21300 = _21297 ^ _21299;
  wire _21301 = _21296 ^ _21300;
  wire _21302 = _664 ^ _11218;
  wire _21303 = uncoded_block[1351] ^ uncoded_block[1355];
  wire _21304 = _21303 ^ _6588;
  wire _21305 = _21302 ^ _21304;
  wire _21306 = uncoded_block[1362] ^ uncoded_block[1365];
  wire _21307 = _21306 ^ _10668;
  wire _21308 = _11226 ^ _10103;
  wire _21309 = _21307 ^ _21308;
  wire _21310 = _21305 ^ _21309;
  wire _21311 = _21301 ^ _21310;
  wire _21312 = uncoded_block[1375] ^ uncoded_block[1382];
  wire _21313 = _21312 ^ _6596;
  wire _21314 = _9578 ^ _7828;
  wire _21315 = _21313 ^ _21314;
  wire _21316 = _5955 ^ _3066;
  wire _21317 = _1519 ^ _3847;
  wire _21318 = _21316 ^ _21317;
  wire _21319 = _21315 ^ _21318;
  wire _21320 = _5961 ^ _6607;
  wire _21321 = _3853 ^ _5967;
  wire _21322 = _21320 ^ _21321;
  wire _21323 = uncoded_block[1428] ^ uncoded_block[1433];
  wire _21324 = uncoded_block[1434] ^ uncoded_block[1441];
  wire _21325 = _21323 ^ _21324;
  wire _21326 = uncoded_block[1444] ^ uncoded_block[1451];
  wire _21327 = _6613 ^ _21326;
  wire _21328 = _21325 ^ _21327;
  wire _21329 = _21322 ^ _21328;
  wire _21330 = _21319 ^ _21329;
  wire _21331 = _21311 ^ _21330;
  wire _21332 = _2328 ^ _6623;
  wire _21333 = _21332 ^ _14988;
  wire _21334 = _3881 ^ _1556;
  wire _21335 = _17484 ^ _21334;
  wire _21336 = _21333 ^ _21335;
  wire _21337 = uncoded_block[1484] ^ uncoded_block[1488];
  wire _21338 = uncoded_block[1489] ^ uncoded_block[1498];
  wire _21339 = _21337 ^ _21338;
  wire _21340 = uncoded_block[1499] ^ uncoded_block[1507];
  wire _21341 = _21340 ^ _5333;
  wire _21342 = _21339 ^ _21341;
  wire _21343 = uncoded_block[1510] ^ uncoded_block[1514];
  wire _21344 = _21343 ^ _3117;
  wire _21345 = _9059 ^ _17499;
  wire _21346 = _21344 ^ _21345;
  wire _21347 = _21342 ^ _21346;
  wire _21348 = _21336 ^ _21347;
  wire _21349 = _6002 ^ _6005;
  wire _21350 = uncoded_block[1534] ^ uncoded_block[1537];
  wire _21351 = _21350 ^ _3908;
  wire _21352 = _21349 ^ _21351;
  wire _21353 = _3909 ^ _7274;
  wire _21354 = _5356 ^ _3131;
  wire _21355 = _21353 ^ _21354;
  wire _21356 = _21352 ^ _21355;
  wire _21357 = _773 ^ _13991;
  wire _21358 = _2376 ^ _11284;
  wire _21359 = _21357 ^ _21358;
  wire _21360 = _2377 ^ _5363;
  wire _21361 = uncoded_block[1572] ^ uncoded_block[1577];
  wire _21362 = _21361 ^ _3921;
  wire _21363 = _21360 ^ _21362;
  wire _21364 = _21359 ^ _21363;
  wire _21365 = _21356 ^ _21364;
  wire _21366 = _21348 ^ _21365;
  wire _21367 = _21331 ^ _21366;
  wire _21368 = _21291 ^ _21367;
  wire _21369 = uncoded_block[1583] ^ uncoded_block[1590];
  wire _21370 = _21369 ^ _792;
  wire _21371 = _3934 ^ _6039;
  wire _21372 = _21370 ^ _21371;
  wire _21373 = _10742 ^ _4662;
  wire _21374 = _7908 ^ _17020;
  wire _21375 = _21373 ^ _21374;
  wire _21376 = _21372 ^ _21375;
  wire _21377 = _9094 ^ _7300;
  wire _21378 = _6046 ^ _3942;
  wire _21379 = _21377 ^ _21378;
  wire _21380 = _18965 ^ _5392;
  wire _21381 = _1646 ^ _6691;
  wire _21382 = _21380 ^ _21381;
  wire _21383 = _21379 ^ _21382;
  wire _21384 = _21376 ^ _21383;
  wire _21385 = _12390 ^ _6055;
  wire _21386 = _4679 ^ _21385;
  wire _21387 = _7320 ^ _12962;
  wire _21388 = _21386 ^ _21387;
  wire _21389 = uncoded_block[1678] ^ uncoded_block[1686];
  wire _21390 = _11319 ^ _21389;
  wire _21391 = _3189 ^ _3967;
  wire _21392 = _21390 ^ _21391;
  wire _21393 = _6707 ^ _6066;
  wire _21394 = uncoded_block[1695] ^ uncoded_block[1697];
  wire _21395 = _21394 ^ _3973;
  wire _21396 = _21393 ^ _21395;
  wire _21397 = _21392 ^ _21396;
  wire _21398 = _21388 ^ _21397;
  wire _21399 = _21384 ^ _21398;
  wire _21400 = uncoded_block[1702] ^ uncoded_block[1710];
  wire _21401 = _21400 ^ _14552;
  wire _21402 = _3988 ^ uncoded_block[1721];
  wire _21403 = _21401 ^ _21402;
  wire _21404 = _21399 ^ _21403;
  wire _21405 = _21368 ^ _21404;
  wire _21406 = _21217 ^ _21405;
  wire _21407 = uncoded_block[0] ^ uncoded_block[3];
  wire _21408 = _21407 ^ _4712;
  wire _21409 = _3995 ^ _17058;
  wire _21410 = _21408 ^ _21409;
  wire _21411 = _2458 ^ _9694;
  wire _21412 = uncoded_block[27] ^ uncoded_block[30];
  wire _21413 = _21412 ^ _2466;
  wire _21414 = _21411 ^ _21413;
  wire _21415 = _21410 ^ _21414;
  wire _21416 = uncoded_block[41] ^ uncoded_block[46];
  wire _21417 = uncoded_block[49] ^ uncoded_block[54];
  wire _21418 = _21416 ^ _21417;
  wire _21419 = _888 ^ _7969;
  wire _21420 = _21418 ^ _21419;
  wire _21421 = _2474 ^ _11357;
  wire _21422 = _6745 ^ _12438;
  wire _21423 = _21421 ^ _21422;
  wire _21424 = _21420 ^ _21423;
  wire _21425 = _21415 ^ _21424;
  wire _21426 = _6749 ^ _2483;
  wire _21427 = _2484 ^ _6757;
  wire _21428 = _21426 ^ _21427;
  wire _21429 = uncoded_block[98] ^ uncoded_block[101];
  wire _21430 = _6758 ^ _21429;
  wire _21431 = _7986 ^ _1722;
  wire _21432 = _21430 ^ _21431;
  wire _21433 = _21428 ^ _21432;
  wire _21434 = _6123 ^ _10816;
  wire _21435 = _54 ^ _14602;
  wire _21436 = _21434 ^ _21435;
  wire _21437 = _15107 ^ _15113;
  wire _21438 = _21436 ^ _21437;
  wire _21439 = _21433 ^ _21438;
  wire _21440 = _21425 ^ _21439;
  wire _21441 = uncoded_block[140] ^ uncoded_block[149];
  wire _21442 = _21441 ^ _70;
  wire _21443 = uncoded_block[152] ^ uncoded_block[157];
  wire _21444 = _21443 ^ _4049;
  wire _21445 = _21442 ^ _21444;
  wire _21446 = _6145 ^ _18578;
  wire _21447 = _21445 ^ _21446;
  wire _21448 = uncoded_block[170] ^ uncoded_block[176];
  wire _21449 = _21448 ^ _17105;
  wire _21450 = uncoded_block[182] ^ uncoded_block[186];
  wire _21451 = _21450 ^ _18111;
  wire _21452 = _21449 ^ _21451;
  wire _21453 = _18113 ^ _89;
  wire _21454 = _10277 ^ _17112;
  wire _21455 = _21453 ^ _21454;
  wire _21456 = _21452 ^ _21455;
  wire _21457 = _21447 ^ _21456;
  wire _21458 = uncoded_block[203] ^ uncoded_block[208];
  wire _21459 = uncoded_block[209] ^ uncoded_block[213];
  wire _21460 = _21458 ^ _21459;
  wire _21461 = _3296 ^ _4787;
  wire _21462 = _21460 ^ _21461;
  wire _21463 = uncoded_block[229] ^ uncoded_block[236];
  wire _21464 = _109 ^ _21463;
  wire _21465 = uncoded_block[241] ^ uncoded_block[244];
  wire _21466 = _5500 ^ _21465;
  wire _21467 = _21464 ^ _21466;
  wire _21468 = _21462 ^ _21467;
  wire _21469 = _11954 ^ _11419;
  wire _21470 = _8618 ^ _21469;
  wire _21471 = _2559 ^ _7438;
  wire _21472 = uncoded_block[267] ^ uncoded_block[271];
  wire _21473 = _6831 ^ _21472;
  wire _21474 = _21471 ^ _21473;
  wire _21475 = _21470 ^ _21474;
  wire _21476 = _21468 ^ _21475;
  wire _21477 = _21457 ^ _21476;
  wire _21478 = _21440 ^ _21477;
  wire _21479 = uncoded_block[272] ^ uncoded_block[276];
  wire _21480 = _21479 ^ _20527;
  wire _21481 = _11967 ^ _991;
  wire _21482 = _21480 ^ _21481;
  wire _21483 = uncoded_block[295] ^ uncoded_block[299];
  wire _21484 = _12509 ^ _21483;
  wire _21485 = _21484 ^ _17640;
  wire _21486 = _21482 ^ _21485;
  wire _21487 = _21017 ^ _3340;
  wire _21488 = _21487 ^ _11440;
  wire _21489 = _9235 ^ _5536;
  wire _21490 = _11982 ^ _21489;
  wire _21491 = _21488 ^ _21490;
  wire _21492 = _21486 ^ _21491;
  wire _21493 = _3353 ^ _6859;
  wire _21494 = uncoded_block[347] ^ uncoded_block[351];
  wire _21495 = _21494 ^ _1028;
  wire _21496 = _21493 ^ _21495;
  wire _21497 = uncoded_block[356] ^ uncoded_block[359];
  wire _21498 = _21497 ^ _18160;
  wire _21499 = _13094 ^ _20056;
  wire _21500 = _21498 ^ _21499;
  wire _21501 = _21496 ^ _21500;
  wire _21502 = uncoded_block[380] ^ uncoded_block[384];
  wire _21503 = _21502 ^ _4149;
  wire _21504 = uncoded_block[389] ^ uncoded_block[393];
  wire _21505 = _21504 ^ _10910;
  wire _21506 = _21503 ^ _21505;
  wire _21507 = _10341 ^ _8088;
  wire _21508 = uncoded_block[414] ^ uncoded_block[416];
  wire _21509 = _12547 ^ _21508;
  wire _21510 = _21507 ^ _21509;
  wire _21511 = _21506 ^ _21510;
  wire _21512 = _21501 ^ _21511;
  wire _21513 = _21492 ^ _21512;
  wire _21514 = _3397 ^ _4874;
  wire _21515 = _21514 ^ _18177;
  wire _21516 = uncoded_block[440] ^ uncoded_block[443];
  wire _21517 = _14690 ^ _21516;
  wire _21518 = _9275 ^ _3411;
  wire _21519 = _21517 ^ _21518;
  wire _21520 = _21515 ^ _21519;
  wire _21521 = _12562 ^ _6261;
  wire _21522 = uncoded_block[459] ^ uncoded_block[462];
  wire _21523 = uncoded_block[468] ^ uncoded_block[471];
  wire _21524 = _21522 ^ _21523;
  wire _21525 = _21521 ^ _21524;
  wire _21526 = uncoded_block[477] ^ uncoded_block[479];
  wire _21527 = _4189 ^ _21526;
  wire _21528 = uncoded_block[483] ^ uncoded_block[485];
  wire _21529 = _4895 ^ _21528;
  wire _21530 = _21527 ^ _21529;
  wire _21531 = _21525 ^ _21530;
  wire _21532 = _21520 ^ _21531;
  wire _21533 = _224 ^ _10370;
  wire _21534 = _12578 ^ _1093;
  wire _21535 = _21533 ^ _21534;
  wire _21536 = uncoded_block[499] ^ uncoded_block[503];
  wire _21537 = _1094 ^ _21536;
  wire _21538 = _10375 ^ _231;
  wire _21539 = _21537 ^ _21538;
  wire _21540 = _21535 ^ _21539;
  wire _21541 = _3444 ^ _237;
  wire _21542 = _14709 ^ _21541;
  wire _21543 = _3447 ^ _10384;
  wire _21544 = _21543 ^ _20605;
  wire _21545 = _21542 ^ _21544;
  wire _21546 = _21540 ^ _21545;
  wire _21547 = _21532 ^ _21546;
  wire _21548 = _21513 ^ _21547;
  wire _21549 = _21478 ^ _21548;
  wire _21550 = uncoded_block[537] ^ uncoded_block[541];
  wire _21551 = _21550 ^ _9854;
  wire _21552 = uncoded_block[545] ^ uncoded_block[550];
  wire _21553 = _21552 ^ _8721;
  wire _21554 = _21551 ^ _21553;
  wire _21555 = uncoded_block[561] ^ uncoded_block[564];
  wire _21556 = _12051 ^ _21555;
  wire _21557 = _1126 ^ _13697;
  wire _21558 = _21556 ^ _21557;
  wire _21559 = _21554 ^ _21558;
  wire _21560 = uncoded_block[573] ^ uncoded_block[576];
  wire _21561 = _17221 ^ _21560;
  wire _21562 = _4946 ^ _1933;
  wire _21563 = _21561 ^ _21562;
  wire _21564 = _1934 ^ _4234;
  wire _21565 = uncoded_block[593] ^ uncoded_block[596];
  wire _21566 = _21565 ^ _12066;
  wire _21567 = _21564 ^ _21566;
  wire _21568 = _21563 ^ _21567;
  wire _21569 = _21559 ^ _21568;
  wire _21570 = _15252 ^ _1942;
  wire _21571 = _6957 ^ _7567;
  wire _21572 = _21570 ^ _21571;
  wire _21573 = _11538 ^ _5659;
  wire _21574 = _21572 ^ _21573;
  wire _21575 = uncoded_block[633] ^ uncoded_block[639];
  wire _21576 = _14745 ^ _21575;
  wire _21577 = _12624 ^ _6338;
  wire _21578 = _21576 ^ _21577;
  wire _21579 = _14234 ^ _6974;
  wire _21580 = _19674 ^ _12630;
  wire _21581 = _21579 ^ _21580;
  wire _21582 = _21578 ^ _21581;
  wire _21583 = _21574 ^ _21582;
  wire _21584 = _21569 ^ _21583;
  wire _21585 = _4978 ^ _16752;
  wire _21586 = uncoded_block[676] ^ uncoded_block[680];
  wire _21587 = _2748 ^ _21586;
  wire _21588 = _21585 ^ _21587;
  wire _21589 = _2750 ^ _11556;
  wire _21590 = _18719 ^ _11564;
  wire _21591 = _21589 ^ _21590;
  wire _21592 = _21588 ^ _21591;
  wire _21593 = uncoded_block[708] ^ uncoded_block[712];
  wire _21594 = _21593 ^ _6366;
  wire _21595 = uncoded_block[717] ^ uncoded_block[721];
  wire _21596 = uncoded_block[723] ^ uncoded_block[731];
  wire _21597 = _21595 ^ _21596;
  wire _21598 = _21594 ^ _21597;
  wire _21599 = _7002 ^ _7605;
  wire _21600 = uncoded_block[742] ^ uncoded_block[746];
  wire _21601 = _1996 ^ _21600;
  wire _21602 = _21599 ^ _21601;
  wire _21603 = _21598 ^ _21602;
  wire _21604 = _21592 ^ _21603;
  wire _21605 = uncoded_block[751] ^ uncoded_block[754];
  wire _21606 = _21605 ^ _3556;
  wire _21607 = _4299 ^ _18740;
  wire _21608 = _21606 ^ _21607;
  wire _21609 = _7616 ^ _7620;
  wire _21610 = uncoded_block[777] ^ uncoded_block[784];
  wire _21611 = _21610 ^ _371;
  wire _21612 = _21609 ^ _21611;
  wire _21613 = _21608 ^ _21612;
  wire _21614 = uncoded_block[793] ^ uncoded_block[797];
  wire _21615 = _372 ^ _21614;
  wire _21616 = _385 ^ _5726;
  wire _21617 = _21615 ^ _21616;
  wire _21618 = _4322 ^ _9397;
  wire _21619 = _21618 ^ _17292;
  wire _21620 = _21617 ^ _21619;
  wire _21621 = _21613 ^ _21620;
  wire _21622 = _21604 ^ _21621;
  wire _21623 = _21584 ^ _21622;
  wire _21624 = _1246 ^ _14807;
  wire _21625 = _401 ^ _7043;
  wire _21626 = _21624 ^ _21625;
  wire _21627 = _7640 ^ _3599;
  wire _21628 = _7643 ^ _6406;
  wire _21629 = _21627 ^ _21628;
  wire _21630 = _21626 ^ _21629;
  wire _21631 = uncoded_block[853] ^ uncoded_block[855];
  wire _21632 = _21631 ^ _20692;
  wire _21633 = _5069 ^ _8244;
  wire _21634 = _21632 ^ _21633;
  wire _21635 = _12151 ^ _20696;
  wire _21636 = uncoded_block[892] ^ uncoded_block[896];
  wire _21637 = _1272 ^ _21636;
  wire _21638 = _21635 ^ _21637;
  wire _21639 = _21634 ^ _21638;
  wire _21640 = _21630 ^ _21639;
  wire _21641 = _1278 ^ _10508;
  wire _21642 = _7070 ^ _1287;
  wire _21643 = _21641 ^ _21642;
  wire _21644 = uncoded_block[915] ^ uncoded_block[918];
  wire _21645 = _21644 ^ _17820;
  wire _21646 = _445 ^ _4370;
  wire _21647 = _21645 ^ _21646;
  wire _21648 = _21643 ^ _21647;
  wire _21649 = uncoded_block[932] ^ uncoded_block[936];
  wire _21650 = _7075 ^ _21649;
  wire _21651 = _10523 ^ _9975;
  wire _21652 = _21650 ^ _21651;
  wire _21653 = uncoded_block[950] ^ uncoded_block[954];
  wire _21654 = _21653 ^ _4384;
  wire _21655 = _7680 ^ _2872;
  wire _21656 = _21654 ^ _21655;
  wire _21657 = _21652 ^ _21656;
  wire _21658 = _21648 ^ _21657;
  wire _21659 = _21640 ^ _21658;
  wire _21660 = uncoded_block[977] ^ uncoded_block[981];
  wire _21661 = _11649 ^ _21660;
  wire _21662 = _2094 ^ _21661;
  wire _21663 = _20221 ^ _1323;
  wire _21664 = _10543 ^ _2107;
  wire _21665 = _21663 ^ _21664;
  wire _21666 = _21662 ^ _21665;
  wire _21667 = _483 ^ _4405;
  wire _21668 = uncoded_block[1009] ^ uncoded_block[1014];
  wire _21669 = _21668 ^ _9996;
  wire _21670 = _21667 ^ _21669;
  wire _21671 = _5135 ^ _8301;
  wire _21672 = _498 ^ _5806;
  wire _21673 = _21671 ^ _21672;
  wire _21674 = _21670 ^ _21673;
  wire _21675 = _21666 ^ _21674;
  wire _21676 = uncoded_block[1033] ^ uncoded_block[1037];
  wire _21677 = _21676 ^ _511;
  wire _21678 = uncoded_block[1042] ^ uncoded_block[1049];
  wire _21679 = _21678 ^ _3682;
  wire _21680 = _21677 ^ _21679;
  wire _21681 = _519 ^ _1363;
  wire _21682 = _10013 ^ _3689;
  wire _21683 = _21681 ^ _21682;
  wire _21684 = _21680 ^ _21683;
  wire _21685 = uncoded_block[1071] ^ uncoded_block[1075];
  wire _21686 = _1366 ^ _21685;
  wire _21687 = uncoded_block[1082] ^ uncoded_block[1085];
  wire _21688 = _21687 ^ _10021;
  wire _21689 = _21686 ^ _21688;
  wire _21690 = _19794 ^ _3708;
  wire _21691 = _1379 ^ _21690;
  wire _21692 = _21689 ^ _21691;
  wire _21693 = _21684 ^ _21692;
  wire _21694 = _21675 ^ _21693;
  wire _21695 = _21659 ^ _21694;
  wire _21696 = _21623 ^ _21695;
  wire _21697 = _21549 ^ _21696;
  wire _21698 = _4450 ^ _10585;
  wire _21699 = _1388 ^ _3714;
  wire _21700 = _21698 ^ _21699;
  wire _21701 = _2942 ^ _2944;
  wire _21702 = uncoded_block[1129] ^ uncoded_block[1137];
  wire _21703 = _15894 ^ _21702;
  wire _21704 = _21701 ^ _21703;
  wire _21705 = _21700 ^ _21704;
  wire _21706 = _2179 ^ _8932;
  wire _21707 = _21706 ^ _4467;
  wire _21708 = _8937 ^ _9500;
  wire _21709 = uncoded_block[1162] ^ uncoded_block[1171];
  wire _21710 = _10043 ^ _21709;
  wire _21711 = _21708 ^ _21710;
  wire _21712 = _21707 ^ _21711;
  wire _21713 = _21705 ^ _21712;
  wire _21714 = _3742 ^ _8944;
  wire _21715 = _16388 ^ _21714;
  wire _21716 = _2200 ^ _5203;
  wire _21717 = _21716 ^ _8950;
  wire _21718 = _21715 ^ _21717;
  wire _21719 = _2209 ^ _5209;
  wire _21720 = _1428 ^ _4498;
  wire _21721 = _21719 ^ _21720;
  wire _21722 = _3765 ^ _7168;
  wire _21723 = uncoded_block[1227] ^ uncoded_block[1231];
  wire _21724 = _11177 ^ _21723;
  wire _21725 = _21722 ^ _21724;
  wire _21726 = _21721 ^ _21725;
  wire _21727 = _21718 ^ _21726;
  wire _21728 = _21713 ^ _21727;
  wire _21729 = _2226 ^ _17416;
  wire _21730 = _8963 ^ _2232;
  wire _21731 = _21729 ^ _21730;
  wire _21732 = uncoded_block[1252] ^ uncoded_block[1257];
  wire _21733 = _6543 ^ _21732;
  wire _21734 = _7781 ^ _3004;
  wire _21735 = _21733 ^ _21734;
  wire _21736 = _21731 ^ _21735;
  wire _21737 = uncoded_block[1272] ^ uncoded_block[1276];
  wire _21738 = _9533 ^ _21737;
  wire _21739 = _21280 ^ _6560;
  wire _21740 = _21738 ^ _21739;
  wire _21741 = uncoded_block[1292] ^ uncoded_block[1296];
  wire _21742 = _11195 ^ _21741;
  wire _21743 = _17927 ^ _16424;
  wire _21744 = _21742 ^ _21743;
  wire _21745 = _21740 ^ _21744;
  wire _21746 = _21736 ^ _21745;
  wire _21747 = _3808 ^ _14430;
  wire _21748 = uncoded_block[1315] ^ uncoded_block[1316];
  wire _21749 = uncoded_block[1320] ^ uncoded_block[1324];
  wire _21750 = _21748 ^ _21749;
  wire _21751 = _21747 ^ _21750;
  wire _21752 = uncoded_block[1325] ^ uncoded_block[1329];
  wire _21753 = uncoded_block[1333] ^ uncoded_block[1335];
  wire _21754 = _21752 ^ _21753;
  wire _21755 = _1497 ^ _5266;
  wire _21756 = _21754 ^ _21755;
  wire _21757 = _21751 ^ _21756;
  wire _21758 = uncoded_block[1348] ^ uncoded_block[1352];
  wire _21759 = _4556 ^ _21758;
  wire _21760 = _673 ^ _12300;
  wire _21761 = _21759 ^ _21760;
  wire _21762 = uncoded_block[1365] ^ uncoded_block[1368];
  wire _21763 = _677 ^ _21762;
  wire _21764 = _680 ^ _10103;
  wire _21765 = _21763 ^ _21764;
  wire _21766 = _21761 ^ _21765;
  wire _21767 = _21757 ^ _21766;
  wire _21768 = _21746 ^ _21767;
  wire _21769 = _21728 ^ _21768;
  wire _21770 = _9573 ^ _2290;
  wire _21771 = uncoded_block[1386] ^ uncoded_block[1391];
  wire _21772 = _9575 ^ _21771;
  wire _21773 = _21770 ^ _21772;
  wire _21774 = uncoded_block[1393] ^ uncoded_block[1395];
  wire _21775 = _21774 ^ _13938;
  wire _21776 = _12315 ^ _3847;
  wire _21777 = _21775 ^ _21776;
  wire _21778 = _21773 ^ _21777;
  wire _21779 = _10113 ^ _13422;
  wire _21780 = uncoded_block[1421] ^ uncoded_block[1425];
  wire _21781 = _21780 ^ _7844;
  wire _21782 = _21779 ^ _21781;
  wire _21783 = uncoded_block[1431] ^ uncoded_block[1435];
  wire _21784 = _9590 ^ _21783;
  wire _21785 = _17470 ^ _3861;
  wire _21786 = _21784 ^ _21785;
  wire _21787 = _21782 ^ _21786;
  wire _21788 = _21778 ^ _21787;
  wire _21789 = _2319 ^ _2322;
  wire _21790 = _2325 ^ _6620;
  wire _21791 = _21789 ^ _21790;
  wire _21792 = _11247 ^ _3088;
  wire _21793 = uncoded_block[1460] ^ uncoded_block[1463];
  wire _21794 = _3089 ^ _21793;
  wire _21795 = _21792 ^ _21794;
  wire _21796 = _21791 ^ _21795;
  wire _21797 = uncoded_block[1470] ^ uncoded_block[1476];
  wire _21798 = _21797 ^ _1556;
  wire _21799 = uncoded_block[1481] ^ uncoded_block[1486];
  wire _21800 = uncoded_block[1487] ^ uncoded_block[1498];
  wire _21801 = _21799 ^ _21800;
  wire _21802 = _21798 ^ _21801;
  wire _21803 = uncoded_block[1499] ^ uncoded_block[1503];
  wire _21804 = _21803 ^ _11264;
  wire _21805 = _13973 ^ _9621;
  wire _21806 = _21804 ^ _21805;
  wire _21807 = _21802 ^ _21806;
  wire _21808 = _21796 ^ _21807;
  wire _21809 = _21788 ^ _21808;
  wire _21810 = _9058 ^ _1579;
  wire _21811 = _5343 ^ _4624;
  wire _21812 = _21810 ^ _21811;
  wire _21813 = _3906 ^ _1590;
  wire _21814 = _16995 ^ _14496;
  wire _21815 = _21813 ^ _21814;
  wire _21816 = _21812 ^ _21815;
  wire _21817 = _6657 ^ _17506;
  wire _21818 = uncoded_block[1559] ^ uncoded_block[1566];
  wire _21819 = _21818 ^ _7891;
  wire _21820 = _21817 ^ _21819;
  wire _21821 = uncoded_block[1579] ^ uncoded_block[1583];
  wire _21822 = _21821 ^ _2386;
  wire _21823 = _4649 ^ _21822;
  wire _21824 = _21820 ^ _21823;
  wire _21825 = _21816 ^ _21824;
  wire _21826 = uncoded_block[1587] ^ uncoded_block[1591];
  wire _21827 = uncoded_block[1592] ^ uncoded_block[1596];
  wire _21828 = _21826 ^ _21827;
  wire _21829 = _1620 ^ _6039;
  wire _21830 = _21828 ^ _21829;
  wire _21831 = uncoded_block[1609] ^ uncoded_block[1614];
  wire _21832 = _21831 ^ _10181;
  wire _21833 = _9095 ^ _13494;
  wire _21834 = _21832 ^ _21833;
  wire _21835 = _21830 ^ _21834;
  wire _21836 = uncoded_block[1634] ^ uncoded_block[1640];
  wire _21837 = _21836 ^ _13500;
  wire _21838 = _10187 ^ _21837;
  wire _21839 = _4674 ^ _15559;
  wire _21840 = _2414 ^ _16049;
  wire _21841 = _21839 ^ _21840;
  wire _21842 = _21838 ^ _21841;
  wire _21843 = _21835 ^ _21842;
  wire _21844 = _21825 ^ _21843;
  wire _21845 = _21809 ^ _21844;
  wire _21846 = _21769 ^ _21845;
  wire _21847 = _12395 ^ _7928;
  wire _21848 = _5401 ^ _10202;
  wire _21849 = _21847 ^ _21848;
  wire _21850 = _3965 ^ _837;
  wire _21851 = _7331 ^ _11874;
  wire _21852 = _21850 ^ _21851;
  wire _21853 = _21849 ^ _21852;
  wire _21854 = _3973 ^ _20437;
  wire _21855 = _21854 ^ _853;
  wire _21856 = _4703 ^ uncoded_block[1721];
  wire _21857 = _21855 ^ _21856;
  wire _21858 = _21853 ^ _21857;
  wire _21859 = _21846 ^ _21858;
  wire _21860 = _21697 ^ _21859;
  wire _21861 = uncoded_block[3] ^ uncoded_block[5];
  wire _21862 = _3209 ^ _21861;
  wire _21863 = _21862 ^ _6084;
  wire _21864 = _868 ^ _9692;
  wire _21865 = _3217 ^ _4000;
  wire _21866 = _21864 ^ _21865;
  wire _21867 = _21863 ^ _21866;
  wire _21868 = _9694 ^ _11344;
  wire _21869 = _2461 ^ _15;
  wire _21870 = _21868 ^ _21869;
  wire _21871 = uncoded_block[38] ^ uncoded_block[40];
  wire _21872 = _3227 ^ _21871;
  wire _21873 = _4008 ^ _22;
  wire _21874 = _21872 ^ _21873;
  wire _21875 = _21870 ^ _21874;
  wire _21876 = _21867 ^ _21875;
  wire _21877 = _23 ^ _6099;
  wire _21878 = _886 ^ _5436;
  wire _21879 = _21877 ^ _21878;
  wire _21880 = _7974 ^ _16085;
  wire _21881 = uncoded_block[75] ^ uncoded_block[78];
  wire _21882 = _3241 ^ _21881;
  wire _21883 = _21880 ^ _21882;
  wire _21884 = _21879 ^ _21883;
  wire _21885 = _6749 ^ _41;
  wire _21886 = _18077 ^ _14591;
  wire _21887 = _21885 ^ _21886;
  wire _21888 = uncoded_block[95] ^ uncoded_block[98];
  wire _21889 = uncoded_block[100] ^ uncoded_block[104];
  wire _21890 = _21888 ^ _21889;
  wire _21891 = uncoded_block[111] ^ uncoded_block[116];
  wire _21892 = _2491 ^ _21891;
  wire _21893 = _21890 ^ _21892;
  wire _21894 = _21887 ^ _21893;
  wire _21895 = _21884 ^ _21894;
  wire _21896 = _21876 ^ _21895;
  wire _21897 = _16592 ^ _3255;
  wire _21898 = uncoded_block[131] ^ uncoded_block[133];
  wire _21899 = _917 ^ _21898;
  wire _21900 = _21897 ^ _21899;
  wire _21901 = uncoded_block[146] ^ uncoded_block[149];
  wire _21902 = _4043 ^ _21901;
  wire _21903 = _21902 ^ _16107;
  wire _21904 = _21900 ^ _21903;
  wire _21905 = uncoded_block[157] ^ uncoded_block[159];
  wire _21906 = uncoded_block[160] ^ uncoded_block[161];
  wire _21907 = _21905 ^ _21906;
  wire _21908 = _4054 ^ _14614;
  wire _21909 = _21907 ^ _21908;
  wire _21910 = _8595 ^ _2525;
  wire _21911 = _2528 ^ _945;
  wire _21912 = _21910 ^ _21911;
  wire _21913 = _21909 ^ _21912;
  wire _21914 = _21904 ^ _21913;
  wire _21915 = _4773 ^ _89;
  wire _21916 = _10277 ^ _2537;
  wire _21917 = _21915 ^ _21916;
  wire _21918 = _4070 ^ _14101;
  wire _21919 = uncoded_block[208] ^ uncoded_block[213];
  wire _21920 = _21919 ^ _9750;
  wire _21921 = _21918 ^ _21920;
  wire _21922 = _21917 ^ _21921;
  wire _21923 = _5497 ^ _17118;
  wire _21924 = _14626 ^ _21923;
  wire _21925 = _21465 ^ _4799;
  wire _21926 = _10290 ^ _21925;
  wire _21927 = _21924 ^ _21926;
  wire _21928 = _21922 ^ _21927;
  wire _21929 = _21914 ^ _21928;
  wire _21930 = _21896 ^ _21929;
  wire _21931 = _2557 ^ _10864;
  wire _21932 = uncoded_block[262] ^ uncoded_block[267];
  wire _21933 = _21932 ^ _4102;
  wire _21934 = _21931 ^ _21933;
  wire _21935 = _6833 ^ _10303;
  wire _21936 = _7446 ^ _6837;
  wire _21937 = _21935 ^ _21936;
  wire _21938 = _21934 ^ _21937;
  wire _21939 = _2571 ^ _5524;
  wire _21940 = _21939 ^ _15162;
  wire _21941 = _4826 ^ _1002;
  wire _21942 = uncoded_block[314] ^ uncoded_block[320];
  wire _21943 = _21942 ^ _15677;
  wire _21944 = _21941 ^ _21943;
  wire _21945 = _21940 ^ _21944;
  wire _21946 = _21938 ^ _21945;
  wire _21947 = uncoded_block[325] ^ uncoded_block[327];
  wire _21948 = _21947 ^ _11983;
  wire _21949 = _7463 ^ _4129;
  wire _21950 = _21948 ^ _21949;
  wire _21951 = _4841 ^ _7465;
  wire _21952 = _4845 ^ _2602;
  wire _21953 = _21951 ^ _21952;
  wire _21954 = _21950 ^ _21953;
  wire _21955 = uncoded_block[364] ^ uncoded_block[369];
  wire _21956 = _21030 ^ _21955;
  wire _21957 = uncoded_block[370] ^ uncoded_block[374];
  wire _21958 = _21957 ^ _8079;
  wire _21959 = _21956 ^ _21958;
  wire _21960 = _14150 ^ _17661;
  wire _21961 = _4151 ^ _10910;
  wire _21962 = _21960 ^ _21961;
  wire _21963 = _21959 ^ _21962;
  wire _21964 = _21954 ^ _21963;
  wire _21965 = _21946 ^ _21964;
  wire _21966 = _1048 ^ _11471;
  wire _21967 = _9810 ^ _1853;
  wire _21968 = _21966 ^ _21967;
  wire _21969 = _194 ^ _11479;
  wire _21970 = _16184 ^ _13117;
  wire _21971 = _21969 ^ _21970;
  wire _21972 = _21968 ^ _21971;
  wire _21973 = _5574 ^ _5577;
  wire _21974 = uncoded_block[442] ^ uncoded_block[444];
  wire _21975 = _21974 ^ _3409;
  wire _21976 = _21973 ^ _21975;
  wire _21977 = _1076 ^ _1873;
  wire _21978 = _14171 ^ _21977;
  wire _21979 = _21976 ^ _21978;
  wire _21980 = _21972 ^ _21979;
  wire _21981 = _3416 ^ _4186;
  wire _21982 = _1082 ^ _11494;
  wire _21983 = _21981 ^ _21982;
  wire _21984 = _8688 ^ _1085;
  wire _21985 = _21984 ^ _21529;
  wire _21986 = _21983 ^ _21985;
  wire _21987 = uncoded_block[492] ^ uncoded_block[496];
  wire _21988 = _21987 ^ _4905;
  wire _21989 = _19135 ^ _5607;
  wire _21990 = _21988 ^ _21989;
  wire _21991 = _8701 ^ _9295;
  wire _21992 = uncoded_block[517] ^ uncoded_block[520];
  wire _21993 = _21992 ^ _3445;
  wire _21994 = _21991 ^ _21993;
  wire _21995 = _21990 ^ _21994;
  wire _21996 = _21986 ^ _21995;
  wire _21997 = _21980 ^ _21996;
  wire _21998 = _21965 ^ _21997;
  wire _21999 = _21930 ^ _21998;
  wire _22000 = _6289 ^ _20602;
  wire _22001 = uncoded_block[529] ^ uncoded_block[537];
  wire _22002 = _22001 ^ _4217;
  wire _22003 = _22000 ^ _22002;
  wire _22004 = uncoded_block[549] ^ uncoded_block[554];
  wire _22005 = _22004 ^ _8724;
  wire _22006 = _17214 ^ _22005;
  wire _22007 = _22003 ^ _22006;
  wire _22008 = _6305 ^ _9320;
  wire _22009 = _3467 ^ _14208;
  wire _22010 = _22008 ^ _22009;
  wire _22011 = _6945 ^ _1133;
  wire _22012 = uncoded_block[583] ^ uncoded_block[585];
  wire _22013 = _1138 ^ _22012;
  wire _22014 = _22011 ^ _22013;
  wire _22015 = _22010 ^ _22014;
  wire _22016 = _22007 ^ _22015;
  wire _22017 = _270 ^ _13705;
  wire _22018 = _3480 ^ _10408;
  wire _22019 = _22017 ^ _22018;
  wire _22020 = _5646 ^ _4957;
  wire _22021 = _20626 ^ _21098;
  wire _22022 = _22020 ^ _22021;
  wire _22023 = _22019 ^ _22022;
  wire _22024 = uncoded_block[620] ^ uncoded_block[624];
  wire _22025 = _6959 ^ _22024;
  wire _22026 = _4964 ^ _5658;
  wire _22027 = _22025 ^ _22026;
  wire _22028 = uncoded_block[631] ^ uncoded_block[636];
  wire _22029 = _22028 ^ _11543;
  wire _22030 = uncoded_block[644] ^ uncoded_block[649];
  wire _22031 = _16241 ^ _22030;
  wire _22032 = _22029 ^ _22031;
  wire _22033 = _22027 ^ _22032;
  wire _22034 = _22023 ^ _22033;
  wire _22035 = _22016 ^ _22034;
  wire _22036 = _20134 ^ _2738;
  wire _22037 = uncoded_block[662] ^ uncoded_block[667];
  wire _22038 = _8172 ^ _22037;
  wire _22039 = _22036 ^ _22038;
  wire _22040 = _311 ^ _2748;
  wire _22041 = _22040 ^ _19190;
  wire _22042 = _22039 ^ _22041;
  wire _22043 = uncoded_block[682] ^ uncoded_block[691];
  wire _22044 = _22043 ^ _3532;
  wire _22045 = uncoded_block[702] ^ uncoded_block[706];
  wire _22046 = _22045 ^ _16761;
  wire _22047 = _22044 ^ _22046;
  wire _22048 = _337 ^ _340;
  wire _22049 = uncoded_block[722] ^ uncoded_block[727];
  wire _22050 = _341 ^ _22049;
  wire _22051 = _22048 ^ _22050;
  wire _22052 = _22047 ^ _22051;
  wire _22053 = _22042 ^ _22052;
  wire _22054 = _3547 ^ _1206;
  wire _22055 = _9372 ^ _22054;
  wire _22056 = _1996 ^ _352;
  wire _22057 = _1998 ^ _4295;
  wire _22058 = _22056 ^ _22057;
  wire _22059 = _22055 ^ _22058;
  wire _22060 = _2778 ^ _3559;
  wire _22061 = _364 ^ _12113;
  wire _22062 = _22060 ^ _22061;
  wire _22063 = uncoded_block[773] ^ uncoded_block[782];
  wire _22064 = _6382 ^ _22063;
  wire _22065 = _7622 ^ _7626;
  wire _22066 = _22064 ^ _22065;
  wire _22067 = _22062 ^ _22066;
  wire _22068 = _22059 ^ _22067;
  wire _22069 = _22053 ^ _22068;
  wire _22070 = _22035 ^ _22069;
  wire _22071 = uncoded_block[802] ^ uncoded_block[805];
  wire _22072 = _1233 ^ _22071;
  wire _22073 = _16791 ^ _15318;
  wire _22074 = _22072 ^ _22073;
  wire _22075 = _11030 ^ _7634;
  wire _22076 = _7037 ^ _4328;
  wire _22077 = _22075 ^ _22076;
  wire _22078 = _22074 ^ _22077;
  wire _22079 = _2812 ^ _4331;
  wire _22080 = _2035 ^ _5057;
  wire _22081 = _22079 ^ _22080;
  wire _22082 = _1256 ^ _3599;
  wire _22083 = _22082 ^ _12147;
  wire _22084 = _22081 ^ _22083;
  wire _22085 = _22078 ^ _22084;
  wire _22086 = _5066 ^ _9948;
  wire _22087 = _9949 ^ _2827;
  wire _22088 = _22086 ^ _22087;
  wire _22089 = _5072 ^ _2831;
  wire _22090 = _2835 ^ _8820;
  wire _22091 = _22089 ^ _22090;
  wire _22092 = _22088 ^ _22091;
  wire _22093 = _2059 ^ _16819;
  wire _22094 = _2841 ^ _5089;
  wire _22095 = _22093 ^ _22094;
  wire _22096 = uncoded_block[903] ^ uncoded_block[908];
  wire _22097 = _22096 ^ _2071;
  wire _22098 = _22097 ^ _3630;
  wire _22099 = _22095 ^ _22098;
  wire _22100 = _22092 ^ _22099;
  wire _22101 = _22085 ^ _22100;
  wire _22102 = _15840 ^ _2857;
  wire _22103 = _21649 ^ _452;
  wire _22104 = _22102 ^ _22103;
  wire _22105 = uncoded_block[939] ^ uncoded_block[943];
  wire _22106 = _22105 ^ _2086;
  wire _22107 = uncoded_block[952] ^ uncoded_block[956];
  wire _22108 = _4381 ^ _22107;
  wire _22109 = _22106 ^ _22108;
  wire _22110 = _22104 ^ _22109;
  wire _22111 = _2090 ^ _1308;
  wire _22112 = uncoded_block[964] ^ uncoded_block[967];
  wire _22113 = uncoded_block[968] ^ uncoded_block[975];
  wire _22114 = _22112 ^ _22113;
  wire _22115 = _22111 ^ _22114;
  wire _22116 = uncoded_block[983] ^ uncoded_block[987];
  wire _22117 = _476 ^ _22116;
  wire _22118 = _480 ^ _7691;
  wire _22119 = _22117 ^ _22118;
  wire _22120 = _22115 ^ _22119;
  wire _22121 = _22110 ^ _22120;
  wire _22122 = uncoded_block[1002] ^ uncoded_block[1004];
  wire _22123 = _22122 ^ _2114;
  wire _22124 = uncoded_block[1009] ^ uncoded_block[1013];
  wire _22125 = _22124 ^ _5134;
  wire _22126 = _22123 ^ _22125;
  wire _22127 = _16853 ^ _5137;
  wire _22128 = _22127 ^ _12753;
  wire _22129 = _22126 ^ _22128;
  wire _22130 = _5806 ^ _2908;
  wire _22131 = uncoded_block[1038] ^ uncoded_block[1043];
  wire _22132 = uncoded_block[1044] ^ uncoded_block[1046];
  wire _22133 = _22131 ^ _22132;
  wire _22134 = _22130 ^ _22133;
  wire _22135 = uncoded_block[1048] ^ uncoded_block[1052];
  wire _22136 = uncoded_block[1053] ^ uncoded_block[1057];
  wire _22137 = _22135 ^ _22136;
  wire _22138 = _22137 ^ _8320;
  wire _22139 = _22134 ^ _22138;
  wire _22140 = _22129 ^ _22139;
  wire _22141 = _22121 ^ _22140;
  wire _22142 = _22101 ^ _22141;
  wire _22143 = _22070 ^ _22142;
  wire _22144 = _21999 ^ _22143;
  wire _22145 = uncoded_block[1068] ^ uncoded_block[1075];
  wire _22146 = _22145 ^ _2147;
  wire _22147 = _8890 ^ _22146;
  wire _22148 = _530 ^ _2928;
  wire _22149 = uncoded_block[1086] ^ uncoded_block[1088];
  wire _22150 = _22149 ^ _536;
  wire _22151 = _22148 ^ _22150;
  wire _22152 = _22147 ^ _22151;
  wire _22153 = _10026 ^ _13316;
  wire _22154 = _2161 ^ _8915;
  wire _22155 = _22153 ^ _22154;
  wire _22156 = _2165 ^ _553;
  wire _22157 = _557 ^ _18832;
  wire _22158 = _22156 ^ _22157;
  wire _22159 = _22155 ^ _22158;
  wire _22160 = _22152 ^ _22159;
  wire _22161 = _4460 ^ _561;
  wire _22162 = uncoded_block[1135] ^ uncoded_block[1141];
  wire _22163 = _22162 ^ _568;
  wire _22164 = _22161 ^ _22163;
  wire _22165 = _4466 ^ _577;
  wire _22166 = _12239 ^ _22165;
  wire _22167 = _22164 ^ _22166;
  wire _22168 = _9500 ^ _578;
  wire _22169 = _3734 ^ _17390;
  wire _22170 = _22168 ^ _22169;
  wire _22171 = _17392 ^ _16898;
  wire _22172 = _11162 ^ _22171;
  wire _22173 = _22170 ^ _22172;
  wire _22174 = _22167 ^ _22173;
  wire _22175 = _22160 ^ _22174;
  wire _22176 = _590 ^ _592;
  wire _22177 = _4486 ^ _5203;
  wire _22178 = _22176 ^ _22177;
  wire _22179 = uncoded_block[1195] ^ uncoded_block[1196];
  wire _22180 = _1420 ^ _22179;
  wire _22181 = _22180 ^ _14909;
  wire _22182 = _22178 ^ _22181;
  wire _22183 = uncoded_block[1204] ^ uncoded_block[1209];
  wire _22184 = _22183 ^ _4496;
  wire _22185 = _2219 ^ _4502;
  wire _22186 = _22184 ^ _22185;
  wire _22187 = _1435 ^ _8377;
  wire _22188 = uncoded_block[1230] ^ uncoded_block[1234];
  wire _22189 = _22188 ^ _3771;
  wire _22190 = _22187 ^ _22189;
  wire _22191 = _22186 ^ _22190;
  wire _22192 = _22182 ^ _22191;
  wire _22193 = uncoded_block[1239] ^ uncoded_block[1249];
  wire _22194 = _22193 ^ _7778;
  wire _22195 = _3001 ^ _7780;
  wire _22196 = _22194 ^ _22195;
  wire _22197 = uncoded_block[1264] ^ uncoded_block[1267];
  wire _22198 = _7781 ^ _22197;
  wire _22199 = _19834 ^ _7792;
  wire _22200 = _22198 ^ _22199;
  wire _22201 = _22196 ^ _22200;
  wire _22202 = _5241 ^ _3797;
  wire _22203 = _639 ^ _8399;
  wire _22204 = _22202 ^ _22203;
  wire _22205 = _3017 ^ _6564;
  wire _22206 = _2254 ^ _8991;
  wire _22207 = _22205 ^ _22206;
  wire _22208 = _22204 ^ _22207;
  wire _22209 = _22201 ^ _22208;
  wire _22210 = _22192 ^ _22209;
  wire _22211 = _22175 ^ _22210;
  wire _22212 = _6572 ^ _1482;
  wire _22213 = _9552 ^ _4540;
  wire _22214 = _22212 ^ _22213;
  wire _22215 = _8997 ^ _5931;
  wire _22216 = _9556 ^ _22215;
  wire _22217 = _22214 ^ _22216;
  wire _22218 = _5932 ^ _14440;
  wire _22219 = uncoded_block[1344] ^ uncoded_block[1349];
  wire _22220 = _22219 ^ _3041;
  wire _22221 = _22218 ^ _22220;
  wire _22222 = _672 ^ _6587;
  wire _22223 = uncoded_block[1359] ^ uncoded_block[1363];
  wire _22224 = uncoded_block[1368] ^ uncoded_block[1374];
  wire _22225 = _22223 ^ _22224;
  wire _22226 = _22222 ^ _22225;
  wire _22227 = _22221 ^ _22226;
  wire _22228 = _22217 ^ _22227;
  wire _22229 = uncoded_block[1375] ^ uncoded_block[1379];
  wire _22230 = _22229 ^ _7219;
  wire _22231 = _3059 ^ _11782;
  wire _22232 = _22230 ^ _22231;
  wire _22233 = _4568 ^ _694;
  wire _22234 = _2296 ^ _3841;
  wire _22235 = _22233 ^ _22234;
  wire _22236 = _22232 ^ _22235;
  wire _22237 = uncoded_block[1409] ^ uncoded_block[1415];
  wire _22238 = _9585 ^ _22237;
  wire _22239 = _11792 ^ _7842;
  wire _22240 = _22238 ^ _22239;
  wire _22241 = _3074 ^ _10684;
  wire _22242 = uncoded_block[1434] ^ uncoded_block[1436];
  wire _22243 = _3081 ^ _22242;
  wire _22244 = _22241 ^ _22243;
  wire _22245 = _22240 ^ _22244;
  wire _22246 = _22236 ^ _22245;
  wire _22247 = _22228 ^ _22246;
  wire _22248 = uncoded_block[1437] ^ uncoded_block[1445];
  wire _22249 = _22248 ^ _3865;
  wire _22250 = _2326 ^ _2328;
  wire _22251 = _22249 ^ _22250;
  wire _22252 = uncoded_block[1455] ^ uncoded_block[1458];
  wire _22253 = _22252 ^ _724;
  wire _22254 = uncoded_block[1465] ^ uncoded_block[1470];
  wire _22255 = _3871 ^ _22254;
  wire _22256 = _22253 ^ _22255;
  wire _22257 = _22251 ^ _22256;
  wire _22258 = _735 ^ _4607;
  wire _22259 = _9609 ^ _22258;
  wire _22260 = _739 ^ _9614;
  wire _22261 = _22260 ^ _9047;
  wire _22262 = _22259 ^ _22261;
  wire _22263 = _22257 ^ _22262;
  wire _22264 = _8466 ^ _4618;
  wire _22265 = _9059 ^ _1581;
  wire _22266 = uncoded_block[1527] ^ uncoded_block[1532];
  wire _22267 = uncoded_block[1534] ^ uncoded_block[1542];
  wire _22268 = _22266 ^ _22267;
  wire _22269 = _22265 ^ _22268;
  wire _22270 = _22264 ^ _22269;
  wire _22271 = _8482 ^ _16501;
  wire _22272 = _770 ^ _4638;
  wire _22273 = _22271 ^ _22272;
  wire _22274 = _4640 ^ _2372;
  wire _22275 = _6019 ^ _7285;
  wire _22276 = _22274 ^ _22275;
  wire _22277 = _22273 ^ _22276;
  wire _22278 = _22270 ^ _22277;
  wire _22279 = _22263 ^ _22278;
  wire _22280 = _22247 ^ _22279;
  wire _22281 = _22211 ^ _22280;
  wire _22282 = uncoded_block[1574] ^ uncoded_block[1580];
  wire _22283 = _9080 ^ _22282;
  wire _22284 = _10171 ^ _5368;
  wire _22285 = _22283 ^ _22284;
  wire _22286 = _13486 ^ _797;
  wire _22287 = _10174 ^ _22286;
  wire _22288 = _22285 ^ _22287;
  wire _22289 = _798 ^ _2396;
  wire _22290 = _5380 ^ _7908;
  wire _22291 = _22289 ^ _22290;
  wire _22292 = uncoded_block[1623] ^ uncoded_block[1626];
  wire _22293 = _7912 ^ _22292;
  wire _22294 = _17021 ^ _22293;
  wire _22295 = _22291 ^ _22294;
  wire _22296 = _22288 ^ _22295;
  wire _22297 = _14525 ^ _3166;
  wire _22298 = _22297 ^ _15556;
  wire _22299 = uncoded_block[1652] ^ uncoded_block[1661];
  wire _22300 = _3172 ^ _22299;
  wire _22301 = _3170 ^ _22300;
  wire _22302 = _22298 ^ _22301;
  wire _22303 = uncoded_block[1663] ^ uncoded_block[1667];
  wire _22304 = _22303 ^ _16052;
  wire _22305 = _8521 ^ _13513;
  wire _22306 = _22304 ^ _22305;
  wire _22307 = _13517 ^ _14543;
  wire _22308 = uncoded_block[1692] ^ uncoded_block[1698];
  wire _22309 = _13519 ^ _22308;
  wire _22310 = _22307 ^ _22309;
  wire _22311 = _22306 ^ _22310;
  wire _22312 = _22302 ^ _22311;
  wire _22313 = _22296 ^ _22312;
  wire _22314 = uncoded_block[1703] ^ uncoded_block[1705];
  wire _22315 = _3973 ^ _22314;
  wire _22316 = uncoded_block[1711] ^ uncoded_block[1713];
  wire _22317 = _848 ^ _22316;
  wire _22318 = _22315 ^ _22317;
  wire _22319 = _854 ^ _13528;
  wire _22320 = _22319 ^ uncoded_block[1721];
  wire _22321 = _22318 ^ _22320;
  wire _22322 = _22313 ^ _22321;
  wire _22323 = _22281 ^ _22322;
  wire _22324 = _22144 ^ _22323;
  wire _22325 = _21407 ^ _6080;
  wire _22326 = uncoded_block[9] ^ uncoded_block[13];
  wire _22327 = _22326 ^ _8545;
  wire _22328 = _22325 ^ _22327;
  wire _22329 = _13537 ^ _3220;
  wire _22330 = _9143 ^ _11;
  wire _22331 = _22329 ^ _22330;
  wire _22332 = _22328 ^ _22331;
  wire _22333 = uncoded_block[32] ^ uncoded_block[35];
  wire _22334 = _22333 ^ _18549;
  wire _22335 = _22334 ^ _24;
  wire _22336 = _3233 ^ _5436;
  wire _22337 = _889 ^ _13553;
  wire _22338 = _22336 ^ _22337;
  wire _22339 = _22335 ^ _22338;
  wire _22340 = _22332 ^ _22339;
  wire _22341 = _32 ^ _11357;
  wire _22342 = _14583 ^ _2481;
  wire _22343 = _22341 ^ _22342;
  wire _22344 = _6750 ^ _19980;
  wire _22345 = uncoded_block[94] ^ uncoded_block[98];
  wire _22346 = _907 ^ _22345;
  wire _22347 = _22344 ^ _22346;
  wire _22348 = _22343 ^ _22347;
  wire _22349 = _4745 ^ _7986;
  wire _22350 = _20957 ^ _4034;
  wire _22351 = _22349 ^ _22350;
  wire _22352 = _16589 ^ _9721;
  wire _22353 = _4751 ^ _1733;
  wire _22354 = _22352 ^ _22353;
  wire _22355 = _22351 ^ _22354;
  wire _22356 = _22348 ^ _22355;
  wire _22357 = _22340 ^ _22356;
  wire _22358 = _923 ^ _1735;
  wire _22359 = _22358 ^ _9181;
  wire _22360 = _6138 ^ _67;
  wire _22361 = _1744 ^ _1748;
  wire _22362 = _22360 ^ _22361;
  wire _22363 = _22359 ^ _22362;
  wire _22364 = _19998 ^ _8589;
  wire _22365 = _11390 ^ _938;
  wire _22366 = _22364 ^ _22365;
  wire _22367 = _3278 ^ _11933;
  wire _22368 = uncoded_block[186] ^ uncoded_block[189];
  wire _22369 = _2528 ^ _22368;
  wire _22370 = _22367 ^ _22369;
  wire _22371 = _22366 ^ _22370;
  wire _22372 = _22363 ^ _22371;
  wire _22373 = _6155 ^ _9745;
  wire _22374 = _6805 ^ _11405;
  wire _22375 = _22373 ^ _22374;
  wire _22376 = _17116 ^ _102;
  wire _22377 = _5497 ^ _109;
  wire _22378 = _22376 ^ _22377;
  wire _22379 = _22375 ^ _22378;
  wire _22380 = uncoded_block[231] ^ uncoded_block[233];
  wire _22381 = _1774 ^ _22380;
  wire _22382 = _968 ^ _10292;
  wire _22383 = _22381 ^ _22382;
  wire _22384 = _6172 ^ _116;
  wire _22385 = _4800 ^ _11419;
  wire _22386 = _22384 ^ _22385;
  wire _22387 = _22383 ^ _22386;
  wire _22388 = _22379 ^ _22387;
  wire _22389 = _22372 ^ _22388;
  wire _22390 = _22357 ^ _22389;
  wire _22391 = _2559 ^ _4095;
  wire _22392 = uncoded_block[268] ^ uncoded_block[271];
  wire _22393 = _21932 ^ _22392;
  wire _22394 = _22391 ^ _22393;
  wire _22395 = _21479 ^ _4105;
  wire _22396 = _992 ^ _10876;
  wire _22397 = _22395 ^ _22396;
  wire _22398 = _22394 ^ _22397;
  wire _22399 = _5524 ^ _2577;
  wire _22400 = _4111 ^ _1000;
  wire _22401 = _22399 ^ _22400;
  wire _22402 = _20536 ^ _16648;
  wire _22403 = _22402 ^ _2581;
  wire _22404 = _22401 ^ _22403;
  wire _22405 = _22398 ^ _22404;
  wire _22406 = _9240 ^ _11984;
  wire _22407 = _4124 ^ _22406;
  wire _22408 = _6217 ^ _11450;
  wire _22409 = _3359 ^ _15179;
  wire _22410 = _22408 ^ _22409;
  wire _22411 = _22407 ^ _22410;
  wire _22412 = _2601 ^ _2606;
  wire _22413 = _3366 ^ _3368;
  wire _22414 = _22412 ^ _22413;
  wire _22415 = _3369 ^ _1838;
  wire _22416 = _13094 ^ _4854;
  wire _22417 = _22415 ^ _22416;
  wire _22418 = _22414 ^ _22417;
  wire _22419 = _22411 ^ _22418;
  wire _22420 = _22405 ^ _22419;
  wire _22421 = _6239 ^ _10908;
  wire _22422 = _3384 ^ _10911;
  wire _22423 = _22421 ^ _22422;
  wire _22424 = _13106 ^ _2629;
  wire _22425 = _4868 ^ _1055;
  wire _22426 = _22424 ^ _22425;
  wire _22427 = _22423 ^ _22426;
  wire _22428 = _8672 ^ _8674;
  wire _22429 = _195 ^ _22428;
  wire _22430 = _6255 ^ _1863;
  wire _22431 = _21052 ^ _3409;
  wire _22432 = _22430 ^ _22431;
  wire _22433 = _22429 ^ _22432;
  wire _22434 = _22427 ^ _22433;
  wire _22435 = _2645 ^ _212;
  wire _22436 = _4885 ^ _15715;
  wire _22437 = _22435 ^ _22436;
  wire _22438 = _4186 ^ _5590;
  wire _22439 = _12567 ^ _22438;
  wire _22440 = _22437 ^ _22439;
  wire _22441 = uncoded_block[484] ^ uncoded_block[491];
  wire _22442 = _8110 ^ _22441;
  wire _22443 = _3432 ^ _13139;
  wire _22444 = _22442 ^ _22443;
  wire _22445 = uncoded_block[503] ^ uncoded_block[509];
  wire _22446 = _3434 ^ _22445;
  wire _22447 = _232 ^ _20598;
  wire _22448 = _22446 ^ _22447;
  wire _22449 = _22444 ^ _22448;
  wire _22450 = _22440 ^ _22449;
  wire _22451 = _22434 ^ _22450;
  wire _22452 = _22420 ^ _22451;
  wire _22453 = _22390 ^ _22452;
  wire _22454 = uncoded_block[522] ^ uncoded_block[525];
  wire _22455 = _1107 ^ _22454;
  wire _22456 = _18208 ^ _12589;
  wire _22457 = _22455 ^ _22456;
  wire _22458 = _4217 ^ _3453;
  wire _22459 = _8134 ^ _6304;
  wire _22460 = _22458 ^ _22459;
  wire _22461 = _22457 ^ _22460;
  wire _22462 = _17710 ^ _1129;
  wire _22463 = _4941 ^ _10967;
  wire _22464 = _22462 ^ _22463;
  wire _22465 = _3475 ^ _19656;
  wire _22466 = _3480 ^ _8149;
  wire _22467 = _22465 ^ _22466;
  wire _22468 = _22464 ^ _22467;
  wire _22469 = _22461 ^ _22468;
  wire _22470 = _14218 ^ _8739;
  wire _22471 = _10410 ^ _22470;
  wire _22472 = _1945 ^ _4243;
  wire _22473 = _1946 ^ _4963;
  wire _22474 = _22472 ^ _22473;
  wire _22475 = _22471 ^ _22474;
  wire _22476 = _4964 ^ _289;
  wire _22477 = _3501 ^ _11543;
  wire _22478 = _22476 ^ _22477;
  wire _22479 = uncoded_block[639] ^ uncoded_block[642];
  wire _22480 = _22479 ^ _4972;
  wire _22481 = _22480 ^ _19673;
  wire _22482 = _22478 ^ _22481;
  wire _22483 = _22475 ^ _22482;
  wire _22484 = _22469 ^ _22483;
  wire _22485 = _3507 ^ _3513;
  wire _22486 = _22485 ^ _19183;
  wire _22487 = _1180 ^ _10440;
  wire _22488 = _7587 ^ _22487;
  wire _22489 = _22486 ^ _22488;
  wire _22490 = _3522 ^ _321;
  wire _22491 = _322 ^ _325;
  wire _22492 = _22490 ^ _22491;
  wire _22493 = uncoded_block[691] ^ uncoded_block[698];
  wire _22494 = _22493 ^ _3532;
  wire _22495 = _18721 ^ _10448;
  wire _22496 = _22494 ^ _22495;
  wire _22497 = _22492 ^ _22496;
  wire _22498 = _22489 ^ _22497;
  wire _22499 = uncoded_block[710] ^ uncoded_block[713];
  wire _22500 = _22499 ^ _1194;
  wire _22501 = _22500 ^ _20147;
  wire _22502 = _10456 ^ _9372;
  wire _22503 = _22501 ^ _22502;
  wire _22504 = uncoded_block[736] ^ uncoded_block[742];
  wire _22505 = _3547 ^ _22504;
  wire _22506 = _5702 ^ _356;
  wire _22507 = _22505 ^ _22506;
  wire _22508 = _11012 ^ _359;
  wire _22509 = _17276 ^ _22508;
  wire _22510 = _22507 ^ _22509;
  wire _22511 = _22503 ^ _22510;
  wire _22512 = _22498 ^ _22511;
  wire _22513 = _22484 ^ _22512;
  wire _22514 = _2783 ^ _365;
  wire _22515 = uncoded_block[769] ^ uncoded_block[774];
  wire _22516 = _22515 ^ _14278;
  wire _22517 = _22514 ^ _22516;
  wire _22518 = _17284 ^ _1224;
  wire _22519 = _12675 ^ _3574;
  wire _22520 = _22518 ^ _22519;
  wire _22521 = _22517 ^ _22520;
  wire _22522 = _5035 ^ _8793;
  wire _22523 = _15814 ^ _11029;
  wire _22524 = _22522 ^ _22523;
  wire _22525 = uncoded_block[817] ^ uncoded_block[819];
  wire _22526 = _2808 ^ _22525;
  wire _22527 = _11600 ^ _4328;
  wire _22528 = _22526 ^ _22527;
  wire _22529 = _22524 ^ _22528;
  wire _22530 = _22521 ^ _22529;
  wire _22531 = _6401 ^ _12137;
  wire _22532 = uncoded_block[837] ^ uncoded_block[841];
  wire _22533 = _22532 ^ _3597;
  wire _22534 = _22531 ^ _22533;
  wire _22535 = uncoded_block[848] ^ uncoded_block[855];
  wire _22536 = _22535 ^ _8812;
  wire _22537 = _5066 ^ _413;
  wire _22538 = _22536 ^ _22537;
  wire _22539 = _22534 ^ _22538;
  wire _22540 = uncoded_block[866] ^ uncoded_block[868];
  wire _22541 = _5069 ^ _22540;
  wire _22542 = _6415 ^ _2831;
  wire _22543 = _22541 ^ _22542;
  wire _22544 = _420 ^ _5079;
  wire _22545 = _2838 ^ _7660;
  wire _22546 = _22544 ^ _22545;
  wire _22547 = _22543 ^ _22546;
  wire _22548 = _22539 ^ _22547;
  wire _22549 = _22530 ^ _22548;
  wire _22550 = _4356 ^ _14315;
  wire _22551 = _6425 ^ _2070;
  wire _22552 = _19252 ^ _3628;
  wire _22553 = _22551 ^ _22552;
  wire _22554 = _22550 ^ _22553;
  wire _22555 = _3629 ^ _17820;
  wire _22556 = _13261 ^ _18316;
  wire _22557 = _22555 ^ _22556;
  wire _22558 = _8262 ^ _8268;
  wire _22559 = uncoded_block[941] ^ uncoded_block[947];
  wire _22560 = _22559 ^ _5777;
  wire _22561 = _22558 ^ _22560;
  wire _22562 = _22557 ^ _22561;
  wire _22563 = _22554 ^ _22562;
  wire _22564 = uncoded_block[953] ^ uncoded_block[956];
  wire _22565 = _1303 ^ _22564;
  wire _22566 = _2090 ^ _2871;
  wire _22567 = _22565 ^ _22566;
  wire _22568 = _1310 ^ _11646;
  wire _22569 = _11087 ^ _7088;
  wire _22570 = _22568 ^ _22569;
  wire _22571 = _22567 ^ _22570;
  wire _22572 = _1315 ^ _5114;
  wire _22573 = _5790 ^ _3659;
  wire _22574 = _22572 ^ _22573;
  wire _22575 = uncoded_block[992] ^ uncoded_block[995];
  wire _22576 = _16338 ^ _22575;
  wire _22577 = _18331 ^ _22576;
  wire _22578 = _22574 ^ _22577;
  wire _22579 = _22571 ^ _22578;
  wire _22580 = _22563 ^ _22579;
  wire _22581 = _22549 ^ _22580;
  wire _22582 = _22513 ^ _22581;
  wire _22583 = _22453 ^ _22582;
  wire _22584 = uncoded_block[997] ^ uncoded_block[1000];
  wire _22585 = uncoded_block[1001] ^ uncoded_block[1004];
  wire _22586 = _22584 ^ _22585;
  wire _22587 = _2886 ^ _5129;
  wire _22588 = _22586 ^ _22587;
  wire _22589 = _13283 ^ _8296;
  wire _22590 = _2891 ^ _5135;
  wire _22591 = _22589 ^ _22590;
  wire _22592 = _22588 ^ _22591;
  wire _22593 = _9454 ^ _18801;
  wire _22594 = _22593 ^ _20232;
  wire _22595 = uncoded_block[1033] ^ uncoded_block[1036];
  wire _22596 = _22595 ^ _1346;
  wire _22597 = uncoded_block[1044] ^ uncoded_block[1048];
  wire _22598 = _512 ^ _22597;
  wire _22599 = _22596 ^ _22598;
  wire _22600 = _22594 ^ _22599;
  wire _22601 = _22592 ^ _22600;
  wire _22602 = uncoded_block[1054] ^ uncoded_block[1061];
  wire _22603 = uncoded_block[1062] ^ uncoded_block[1068];
  wire _22604 = _22602 ^ _22603;
  wire _22605 = _1366 ^ _5832;
  wire _22606 = _22604 ^ _22605;
  wire _22607 = _533 ^ _11687;
  wire _22608 = _12773 ^ _22607;
  wire _22609 = _22606 ^ _22608;
  wire _22610 = uncoded_block[1091] ^ uncoded_block[1093];
  wire _22611 = _12774 ^ _22610;
  wire _22612 = _1380 ^ _545;
  wire _22613 = _22611 ^ _22612;
  wire _22614 = uncoded_block[1115] ^ uncoded_block[1119];
  wire _22615 = _4451 ^ _22614;
  wire _22616 = _19312 ^ _22615;
  wire _22617 = _22613 ^ _22616;
  wire _22618 = _22609 ^ _22617;
  wire _22619 = _22601 ^ _22618;
  wire _22620 = _14376 ^ _8343;
  wire _22621 = _14887 ^ _8929;
  wire _22622 = _22620 ^ _22621;
  wire _22623 = _5859 ^ _8932;
  wire _22624 = _2956 ^ _578;
  wire _22625 = _22623 ^ _22624;
  wire _22626 = _22622 ^ _22625;
  wire _22627 = uncoded_block[1162] ^ uncoded_block[1163];
  wire _22628 = _7748 ^ _22627;
  wire _22629 = _22628 ^ _14896;
  wire _22630 = _11161 ^ _1410;
  wire _22631 = _22630 ^ _5196;
  wire _22632 = _22629 ^ _22631;
  wire _22633 = _22626 ^ _22632;
  wire _22634 = uncoded_block[1184] ^ uncoded_block[1194];
  wire _22635 = _22634 ^ _5882;
  wire _22636 = _18389 ^ _2978;
  wire _22637 = _22635 ^ _22636;
  wire _22638 = _17407 ^ _2982;
  wire _22639 = _606 ^ _5215;
  wire _22640 = _22638 ^ _22639;
  wire _22641 = _22637 ^ _22640;
  wire _22642 = _7168 ^ _12819;
  wire _22643 = _18400 ^ _18404;
  wire _22644 = _22642 ^ _22643;
  wire _22645 = _8962 ^ _13365;
  wire _22646 = _3773 ^ _22645;
  wire _22647 = _22644 ^ _22646;
  wire _22648 = _22641 ^ _22647;
  wire _22649 = _22633 ^ _22648;
  wire _22650 = _22619 ^ _22649;
  wire _22651 = uncoded_block[1253] ^ uncoded_block[1256];
  wire _22652 = _1451 ^ _22651;
  wire _22653 = uncoded_block[1262] ^ uncoded_block[1267];
  wire _22654 = _1456 ^ _22653;
  wire _22655 = _22652 ^ _22654;
  wire _22656 = _2245 ^ _16419;
  wire _22657 = uncoded_block[1279] ^ uncoded_block[1285];
  wire _22658 = _2247 ^ _22657;
  wire _22659 = _22656 ^ _22658;
  wire _22660 = _22655 ^ _22659;
  wire _22661 = _5913 ^ _8399;
  wire _22662 = uncoded_block[1297] ^ uncoded_block[1301];
  wire _22663 = _3015 ^ _22662;
  wire _22664 = _22661 ^ _22663;
  wire _22665 = uncoded_block[1303] ^ uncoded_block[1305];
  wire _22666 = _22665 ^ _8991;
  wire _22667 = _6572 ^ _8407;
  wire _22668 = _22666 ^ _22667;
  wire _22669 = _22664 ^ _22668;
  wire _22670 = _22660 ^ _22669;
  wire _22671 = _14433 ^ _11206;
  wire _22672 = uncoded_block[1332] ^ uncoded_block[1337];
  wire _22673 = _1494 ^ _22672;
  wire _22674 = _13399 ^ _1497;
  wire _22675 = _22673 ^ _22674;
  wire _22676 = _22671 ^ _22675;
  wire _22677 = _5266 ^ _5268;
  wire _22678 = uncoded_block[1352] ^ uncoded_block[1357];
  wire _22679 = _22678 ^ _5273;
  wire _22680 = _22677 ^ _22679;
  wire _22681 = _3045 ^ _10665;
  wire _22682 = _12302 ^ _3832;
  wire _22683 = _22681 ^ _22682;
  wire _22684 = _22680 ^ _22683;
  wire _22685 = _22676 ^ _22684;
  wire _22686 = _22670 ^ _22685;
  wire _22687 = uncoded_block[1381] ^ uncoded_block[1384];
  wire _22688 = _2290 ^ _22687;
  wire _22689 = _18444 ^ _7828;
  wire _22690 = _22688 ^ _22689;
  wire _22691 = _694 ^ _4572;
  wire _22692 = _3847 ^ _9585;
  wire _22693 = _22691 ^ _22692;
  wire _22694 = _22690 ^ _22693;
  wire _22695 = _14460 ^ _5965;
  wire _22696 = _17465 ^ _1535;
  wire _22697 = _22695 ^ _22696;
  wire _22698 = _22694 ^ _22697;
  wire _22699 = _13432 ^ _1541;
  wire _22700 = _9033 ^ _2325;
  wire _22701 = _22699 ^ _22700;
  wire _22702 = _2326 ^ _3868;
  wire _22703 = uncoded_block[1461] ^ uncoded_block[1467];
  wire _22704 = _724 ^ _22703;
  wire _22705 = _22702 ^ _22704;
  wire _22706 = _22701 ^ _22705;
  wire _22707 = uncoded_block[1472] ^ uncoded_block[1475];
  wire _22708 = _5983 ^ _22707;
  wire _22709 = _9610 ^ _1558;
  wire _22710 = _22708 ^ _22709;
  wire _22711 = uncoded_block[1483] ^ uncoded_block[1487];
  wire _22712 = _22711 ^ _1563;
  wire _22713 = _5329 ^ _10712;
  wire _22714 = _22712 ^ _22713;
  wire _22715 = _22710 ^ _22714;
  wire _22716 = _22706 ^ _22715;
  wire _22717 = _22698 ^ _22716;
  wire _22718 = _22686 ^ _22717;
  wire _22719 = _22650 ^ _22718;
  wire _22720 = _1571 ^ _7259;
  wire _22721 = _4616 ^ _9053;
  wire _22722 = _22720 ^ _22721;
  wire _22723 = uncoded_block[1520] ^ uncoded_block[1523];
  wire _22724 = _3117 ^ _22723;
  wire _22725 = _6001 ^ _3905;
  wire _22726 = _22724 ^ _22725;
  wire _22727 = _22722 ^ _22726;
  wire _22728 = _12915 ^ _5350;
  wire _22729 = _20387 ^ _18492;
  wire _22730 = _22728 ^ _22729;
  wire _22731 = uncoded_block[1555] ^ uncoded_block[1556];
  wire _22732 = _767 ^ _22731;
  wire _22733 = _22732 ^ _775;
  wire _22734 = _22730 ^ _22733;
  wire _22735 = _22727 ^ _22734;
  wire _22736 = uncoded_block[1563] ^ uncoded_block[1569];
  wire _22737 = _22736 ^ _5363;
  wire _22738 = _22737 ^ _18950;
  wire _22739 = _2383 ^ _1612;
  wire _22740 = _16515 ^ _791;
  wire _22741 = _22739 ^ _22740;
  wire _22742 = _22738 ^ _22741;
  wire _22743 = _4654 ^ _13486;
  wire _22744 = _5373 ^ _6039;
  wire _22745 = _22743 ^ _22744;
  wire _22746 = uncoded_block[1607] ^ uncoded_block[1612];
  wire _22747 = _3153 ^ _22746;
  wire _22748 = _10181 ^ _7912;
  wire _22749 = _22747 ^ _22748;
  wire _22750 = _22745 ^ _22749;
  wire _22751 = _22742 ^ _22750;
  wire _22752 = _22735 ^ _22751;
  wire _22753 = _10185 ^ _14525;
  wire _22754 = _15551 ^ _2405;
  wire _22755 = _22753 ^ _22754;
  wire _22756 = uncoded_block[1644] ^ uncoded_block[1649];
  wire _22757 = _2408 ^ _22756;
  wire _22758 = _4677 ^ _14011;
  wire _22759 = _22757 ^ _22758;
  wire _22760 = _22755 ^ _22759;
  wire _22761 = uncoded_block[1663] ^ uncoded_block[1665];
  wire _22762 = _10196 ^ _22761;
  wire _22763 = uncoded_block[1670] ^ uncoded_block[1673];
  wire _22764 = _5399 ^ _22763;
  wire _22765 = _22762 ^ _22764;
  wire _22766 = _3962 ^ _10766;
  wire _22767 = _3187 ^ _20429;
  wire _22768 = _22766 ^ _22767;
  wire _22769 = _22765 ^ _22768;
  wire _22770 = _22760 ^ _22769;
  wire _22771 = _840 ^ _9677;
  wire _22772 = uncoded_block[1698] ^ uncoded_block[1701];
  wire _22773 = uncoded_block[1702] ^ uncoded_block[1705];
  wire _22774 = _22772 ^ _22773;
  wire _22775 = _22771 ^ _22774;
  wire _22776 = _2435 ^ _10778;
  wire _22777 = _852 ^ _6072;
  wire _22778 = _22776 ^ _22777;
  wire _22779 = _22775 ^ _22778;
  wire _22780 = _22779 ^ _21402;
  wire _22781 = _22770 ^ _22780;
  wire _22782 = _22752 ^ _22781;
  wire _22783 = _22719 ^ _22782;
  wire _22784 = _22583 ^ _22783;
  wire _22785 = _3209 ^ _1;
  wire _22786 = _22785 ^ _6725;
  wire _22787 = _1686 ^ _868;
  wire _22788 = _22787 ^ _20450;
  wire _22789 = _22786 ^ _22788;
  wire _22790 = uncoded_block[24] ^ uncoded_block[26];
  wire _22791 = _4000 ^ _22790;
  wire _22792 = _11344 ^ _2461;
  wire _22793 = _22791 ^ _22792;
  wire _22794 = _6095 ^ _11347;
  wire _22795 = uncoded_block[46] ^ uncoded_block[49];
  wire _22796 = _17065 ^ _22795;
  wire _22797 = _22794 ^ _22796;
  wire _22798 = _22793 ^ _22797;
  wire _22799 = _22789 ^ _22798;
  wire _22800 = _5435 ^ _16572;
  wire _22801 = _889 ^ _2474;
  wire _22802 = _22800 ^ _22801;
  wire _22803 = uncoded_block[68] ^ uncoded_block[72];
  wire _22804 = _22803 ^ _4020;
  wire _22805 = uncoded_block[79] ^ uncoded_block[83];
  wire _22806 = _22805 ^ _17578;
  wire _22807 = _22804 ^ _22806;
  wire _22808 = _22802 ^ _22807;
  wire _22809 = _4026 ^ _7375;
  wire _22810 = _15096 ^ _22809;
  wire _22811 = _21889 ^ _50;
  wire _22812 = _1726 ^ _18090;
  wire _22813 = _22811 ^ _22812;
  wire _22814 = _22810 ^ _22813;
  wire _22815 = _22808 ^ _22814;
  wire _22816 = _22799 ^ _22815;
  wire _22817 = uncoded_block[127] ^ uncoded_block[130];
  wire _22818 = _10819 ^ _22817;
  wire _22819 = uncoded_block[134] ^ uncoded_block[137];
  wire _22820 = _1735 ^ _22819;
  wire _22821 = _22818 ^ _22820;
  wire _22822 = _64 ^ _4043;
  wire _22823 = _1742 ^ _6780;
  wire _22824 = _22822 ^ _22823;
  wire _22825 = _22821 ^ _22824;
  wire _22826 = _3268 ^ _9186;
  wire _22827 = _1748 ^ _15118;
  wire _22828 = _22826 ^ _22827;
  wire _22829 = uncoded_block[162] ^ uncoded_block[170];
  wire _22830 = _22829 ^ _19539;
  wire _22831 = _6149 ^ _11933;
  wire _22832 = _22830 ^ _22831;
  wire _22833 = _22828 ^ _22832;
  wire _22834 = _22825 ^ _22833;
  wire _22835 = _8009 ^ _86;
  wire _22836 = _22835 ^ _20983;
  wire _22837 = uncoded_block[196] ^ uncoded_block[200];
  wire _22838 = _1763 ^ _22837;
  wire _22839 = _3289 ^ _1764;
  wire _22840 = _22838 ^ _22839;
  wire _22841 = _22836 ^ _22840;
  wire _22842 = _11405 ^ _1767;
  wire _22843 = _22842 ^ _8607;
  wire _22844 = _4788 ^ _17617;
  wire _22845 = uncoded_block[228] ^ uncoded_block[232];
  wire _22846 = _22845 ^ _2550;
  wire _22847 = _22844 ^ _22846;
  wire _22848 = _22843 ^ _22847;
  wire _22849 = _22841 ^ _22848;
  wire _22850 = _22834 ^ _22849;
  wire _22851 = _22816 ^ _22850;
  wire _22852 = _10289 ^ _6172;
  wire _22853 = _6179 ^ _7434;
  wire _22854 = _22852 ^ _22853;
  wire _22855 = uncoded_block[260] ^ uncoded_block[264];
  wire _22856 = _22855 ^ _127;
  wire _22857 = _11420 ^ _22856;
  wire _22858 = _22854 ^ _22857;
  wire _22859 = _14124 ^ _6833;
  wire _22860 = _22859 ^ _9771;
  wire _22861 = _9226 ^ _4819;
  wire _22862 = _4820 ^ _3332;
  wire _22863 = _22861 ^ _22862;
  wire _22864 = _22860 ^ _22863;
  wire _22865 = _22858 ^ _22864;
  wire _22866 = uncoded_block[309] ^ uncoded_block[311];
  wire _22867 = _4824 ^ _22866;
  wire _22868 = _145 ^ _20539;
  wire _22869 = _22867 ^ _22868;
  wire _22870 = _6850 ^ _15677;
  wire _22871 = _22870 ^ _11982;
  wire _22872 = _22869 ^ _22871;
  wire _22873 = uncoded_block[332] ^ uncoded_block[336];
  wire _22874 = _2586 ^ _22873;
  wire _22875 = _6217 ^ _4841;
  wire _22876 = _22874 ^ _22875;
  wire _22877 = _8652 ^ _5541;
  wire _22878 = _1024 ^ _2601;
  wire _22879 = _22877 ^ _22878;
  wire _22880 = _22876 ^ _22879;
  wire _22881 = _22872 ^ _22880;
  wire _22882 = _22865 ^ _22881;
  wire _22883 = uncoded_block[357] ^ uncoded_block[361];
  wire _22884 = _22883 ^ _21030;
  wire _22885 = _168 ^ _16662;
  wire _22886 = _22884 ^ _22885;
  wire _22887 = _19596 ^ _12539;
  wire _22888 = _22886 ^ _22887;
  wire _22889 = _3380 ^ _6239;
  wire _22890 = _5554 ^ _4152;
  wire _22891 = _22889 ^ _22890;
  wire _22892 = _3384 ^ _1048;
  wire _22893 = _22892 ^ _20565;
  wire _22894 = _22891 ^ _22893;
  wire _22895 = _22888 ^ _22894;
  wire _22896 = _190 ^ _3394;
  wire _22897 = _6249 ^ _14160;
  wire _22898 = _22896 ^ _22897;
  wire _22899 = _8671 ^ _16184;
  wire _22900 = _200 ^ _6255;
  wire _22901 = _22899 ^ _22900;
  wire _22902 = _22898 ^ _22901;
  wire _22903 = uncoded_block[448] ^ uncoded_block[452];
  wire _22904 = _13122 ^ _22903;
  wire _22905 = _16681 ^ _22904;
  wire _22906 = _1867 ^ _20078;
  wire _22907 = uncoded_block[461] ^ uncoded_block[466];
  wire _22908 = _22907 ^ _3418;
  wire _22909 = _22906 ^ _22908;
  wire _22910 = _22905 ^ _22909;
  wire _22911 = _22902 ^ _22910;
  wire _22912 = _22895 ^ _22911;
  wire _22913 = _22882 ^ _22912;
  wire _22914 = _22851 ^ _22913;
  wire _22915 = _4188 ^ _13132;
  wire _22916 = _16693 ^ _1086;
  wire _22917 = _22915 ^ _22916;
  wire _22918 = uncoded_block[494] ^ uncoded_block[500];
  wire _22919 = _3424 ^ _22918;
  wire _22920 = _16697 ^ _22919;
  wire _22921 = _22917 ^ _22920;
  wire _22922 = _7521 ^ _5607;
  wire _22923 = _22922 ^ _21991;
  wire _22924 = uncoded_block[522] ^ uncoded_block[528];
  wire _22925 = _14193 ^ _22924;
  wire _22926 = uncoded_block[533] ^ uncoded_block[538];
  wire _22927 = _1901 ^ _22926;
  wire _22928 = _22925 ^ _22927;
  wire _22929 = _22923 ^ _22928;
  wire _22930 = _22921 ^ _22929;
  wire _22931 = _8718 ^ _7541;
  wire _22932 = _6300 ^ _4933;
  wire _22933 = _22931 ^ _22932;
  wire _22934 = uncoded_block[551] ^ uncoded_block[555];
  wire _22935 = _22934 ^ _1916;
  wire _22936 = uncoded_block[569] ^ uncoded_block[580];
  wire _22937 = _9320 ^ _22936;
  wire _22938 = _22935 ^ _22937;
  wire _22939 = _22933 ^ _22938;
  wire _22940 = _4946 ^ _270;
  wire _22941 = _4950 ^ _20618;
  wire _22942 = _22940 ^ _22941;
  wire _22943 = _15247 ^ _12066;
  wire _22944 = _22943 ^ _15253;
  wire _22945 = _22942 ^ _22944;
  wire _22946 = _22939 ^ _22945;
  wire _22947 = _22930 ^ _22946;
  wire _22948 = uncoded_block[608] ^ uncoded_block[620];
  wire _22949 = _22948 ^ _2719;
  wire _22950 = uncoded_block[631] ^ uncoded_block[633];
  wire _22951 = _8159 ^ _22950;
  wire _22952 = _22949 ^ _22951;
  wire _22953 = _6331 ^ _4249;
  wire _22954 = uncoded_block[643] ^ uncoded_block[648];
  wire _22955 = _22954 ^ _1960;
  wire _22956 = _22953 ^ _22955;
  wire _22957 = _22952 ^ _22956;
  wire _22958 = uncoded_block[653] ^ uncoded_block[658];
  wire _22959 = _22958 ^ _20638;
  wire _22960 = uncoded_block[663] ^ uncoded_block[668];
  wire _22961 = _22960 ^ _311;
  wire _22962 = _22959 ^ _22961;
  wire _22963 = uncoded_block[681] ^ uncoded_block[685];
  wire _22964 = _17747 ^ _22963;
  wire _22965 = _322 ^ _2754;
  wire _22966 = _22964 ^ _22965;
  wire _22967 = _22962 ^ _22966;
  wire _22968 = _22957 ^ _22967;
  wire _22969 = _8186 ^ _12641;
  wire _22970 = _18721 ^ _336;
  wire _22971 = _22969 ^ _22970;
  wire _22972 = _1194 ^ _6367;
  wire _22973 = _22972 ^ _21130;
  wire _22974 = _22971 ^ _22973;
  wire _22975 = uncoded_block[733] ^ uncoded_block[737];
  wire _22976 = _13749 ^ _22975;
  wire _22977 = _1996 ^ _5010;
  wire _22978 = _22976 ^ _22977;
  wire _22979 = _1998 ^ _5704;
  wire _22980 = _22979 ^ _4296;
  wire _22981 = _22978 ^ _22980;
  wire _22982 = _22974 ^ _22981;
  wire _22983 = _22968 ^ _22982;
  wire _22984 = _22947 ^ _22983;
  wire _22985 = _4298 ^ _3559;
  wire _22986 = _22985 ^ _14782;
  wire _22987 = _10470 ^ _1221;
  wire _22988 = _5711 ^ _3567;
  wire _22989 = _22987 ^ _22988;
  wire _22990 = _22986 ^ _22989;
  wire _22991 = uncoded_block[780] ^ uncoded_block[783];
  wire _22992 = _22991 ^ _4311;
  wire _22993 = _7626 ^ _11024;
  wire _22994 = _22992 ^ _22993;
  wire _22995 = _382 ^ _386;
  wire _22996 = _389 ^ _8228;
  wire _22997 = _22995 ^ _22996;
  wire _22998 = _22994 ^ _22997;
  wire _22999 = _22990 ^ _22998;
  wire _23000 = _10485 ^ _4325;
  wire _23001 = _1242 ^ _6399;
  wire _23002 = _23000 ^ _23001;
  wire _23003 = uncoded_block[829] ^ uncoded_block[834];
  wire _23004 = _1247 ^ _23003;
  wire _23005 = _5054 ^ _5057;
  wire _23006 = _23004 ^ _23005;
  wire _23007 = _23002 ^ _23006;
  wire _23008 = _5741 ^ _2821;
  wire _23009 = _1258 ^ _23008;
  wire _23010 = uncoded_block[858] ^ uncoded_block[861];
  wire _23011 = _3600 ^ _23010;
  wire _23012 = _413 ^ _2827;
  wire _23013 = _23011 ^ _23012;
  wire _23014 = _23009 ^ _23013;
  wire _23015 = _23007 ^ _23014;
  wire _23016 = _22999 ^ _23015;
  wire _23017 = _12150 ^ _1269;
  wire _23018 = _23017 ^ _19730;
  wire _23019 = _18770 ^ _4354;
  wire _23020 = _23019 ^ _15834;
  wire _23021 = _23018 ^ _23020;
  wire _23022 = uncoded_block[908] ^ uncoded_block[913];
  wire _23023 = _2844 ^ _23022;
  wire _23024 = _9959 ^ _23023;
  wire _23025 = _12712 ^ _15350;
  wire _23026 = uncoded_block[927] ^ uncoded_block[934];
  wire _23027 = _16315 ^ _23026;
  wire _23028 = _23025 ^ _23027;
  wire _23029 = _23024 ^ _23028;
  wire _23030 = _23021 ^ _23029;
  wire _23031 = _7674 ^ _16834;
  wire _23032 = _22107 ^ _9979;
  wire _23033 = _10529 ^ _11646;
  wire _23034 = _23032 ^ _23033;
  wire _23035 = _23031 ^ _23034;
  wire _23036 = _5785 ^ _470;
  wire _23037 = _23036 ^ _21199;
  wire _23038 = uncoded_block[982] ^ uncoded_block[985];
  wire _23039 = _23038 ^ _8856;
  wire _23040 = uncoded_block[990] ^ uncoded_block[995];
  wire _23041 = _23040 ^ _480;
  wire _23042 = _23039 ^ _23041;
  wire _23043 = _23037 ^ _23042;
  wire _23044 = _23035 ^ _23043;
  wire _23045 = _23030 ^ _23044;
  wire _23046 = _23016 ^ _23045;
  wire _23047 = _22984 ^ _23046;
  wire _23048 = _22914 ^ _23047;
  wire _23049 = _484 ^ _486;
  wire _23050 = _18335 ^ _23049;
  wire _23051 = _487 ^ _4412;
  wire _23052 = _8871 ^ _1338;
  wire _23053 = _23051 ^ _23052;
  wire _23054 = _23050 ^ _23053;
  wire _23055 = uncoded_block[1031] ^ uncoded_block[1037];
  wire _23056 = _23055 ^ _6475;
  wire _23057 = _2899 ^ _23056;
  wire _23058 = _1357 ^ _12762;
  wire _23059 = _22598 ^ _23058;
  wire _23060 = _23057 ^ _23059;
  wire _23061 = _23054 ^ _23060;
  wire _23062 = uncoded_block[1055] ^ uncoded_block[1058];
  wire _23063 = _23062 ^ _6483;
  wire _23064 = _2917 ^ _11122;
  wire _23065 = _23063 ^ _23064;
  wire _23066 = _527 ^ _2146;
  wire _23067 = _2147 ^ _21228;
  wire _23068 = _23066 ^ _23067;
  wire _23069 = _23065 ^ _23068;
  wire _23070 = _12774 ^ _5840;
  wire _23071 = uncoded_block[1094] ^ uncoded_block[1098];
  wire _23072 = _23071 ^ _2160;
  wire _23073 = _23070 ^ _23072;
  wire _23074 = _2161 ^ _6494;
  wire _23075 = uncoded_block[1113] ^ uncoded_block[1115];
  wire _23076 = _4451 ^ _23075;
  wire _23077 = _23074 ^ _23076;
  wire _23078 = _23073 ^ _23077;
  wire _23079 = _23069 ^ _23078;
  wire _23080 = _23061 ^ _23079;
  wire _23081 = _2944 ^ _4459;
  wire _23082 = _21699 ^ _23081;
  wire _23083 = _18371 ^ _1393;
  wire _23084 = _10591 ^ _8929;
  wire _23085 = _23083 ^ _23084;
  wire _23086 = _23082 ^ _23085;
  wire _23087 = _565 ^ _567;
  wire _23088 = _568 ^ _9499;
  wire _23089 = _23087 ^ _23088;
  wire _23090 = _7143 ^ _11711;
  wire _23091 = _2964 ^ _4476;
  wire _23092 = _23090 ^ _23091;
  wire _23093 = _23089 ^ _23092;
  wire _23094 = _23086 ^ _23093;
  wire _23095 = _11161 ^ _17392;
  wire _23096 = _23095 ^ _8943;
  wire _23097 = uncoded_block[1186] ^ uncoded_block[1190];
  wire _23098 = _4486 ^ _23097;
  wire _23099 = _3749 ^ _22179;
  wire _23100 = _23098 ^ _23099;
  wire _23101 = _23096 ^ _23100;
  wire _23102 = _7758 ^ _1425;
  wire _23103 = _2216 ^ _2981;
  wire _23104 = _23102 ^ _23103;
  wire _23105 = uncoded_block[1216] ^ uncoded_block[1220];
  wire _23106 = _2982 ^ _23105;
  wire _23107 = uncoded_block[1226] ^ uncoded_block[1232];
  wire _23108 = _23107 ^ _1442;
  wire _23109 = _23106 ^ _23108;
  wire _23110 = _23104 ^ _23109;
  wire _23111 = _23101 ^ _23110;
  wire _23112 = _23094 ^ _23111;
  wire _23113 = _23080 ^ _23112;
  wire _23114 = uncoded_block[1241] ^ uncoded_block[1246];
  wire _23115 = _23114 ^ _1451;
  wire _23116 = _5222 ^ _23115;
  wire _23117 = _8385 ^ _2236;
  wire _23118 = _3784 ^ _3004;
  wire _23119 = _23117 ^ _23118;
  wire _23120 = _23116 ^ _23119;
  wire _23121 = _21737 ^ _21280;
  wire _23122 = _10635 ^ _23121;
  wire _23123 = uncoded_block[1280] ^ uncoded_block[1282];
  wire _23124 = uncoded_block[1285] ^ uncoded_block[1288];
  wire _23125 = _23123 ^ _23124;
  wire _23126 = _4529 ^ _8399;
  wire _23127 = _23125 ^ _23126;
  wire _23128 = _23122 ^ _23127;
  wire _23129 = _23120 ^ _23128;
  wire _23130 = _19369 ^ _6564;
  wire _23131 = uncoded_block[1303] ^ uncoded_block[1307];
  wire _23132 = _16424 ^ _23131;
  wire _23133 = _23130 ^ _23132;
  wire _23134 = uncoded_block[1317] ^ uncoded_block[1319];
  wire _23135 = _1483 ^ _23134;
  wire _23136 = _22667 ^ _23135;
  wire _23137 = _23133 ^ _23136;
  wire _23138 = _21749 ^ _656;
  wire _23139 = uncoded_block[1328] ^ uncoded_block[1331];
  wire _23140 = _23139 ^ _21753;
  wire _23141 = _23138 ^ _23140;
  wire _23142 = _5259 ^ _5261;
  wire _23143 = _5262 ^ _7206;
  wire _23144 = _23142 ^ _23143;
  wire _23145 = _23141 ^ _23144;
  wire _23146 = _23137 ^ _23145;
  wire _23147 = _23129 ^ _23146;
  wire _23148 = uncoded_block[1360] ^ uncoded_block[1365];
  wire _23149 = _15477 ^ _23148;
  wire _23150 = _15474 ^ _23149;
  wire _23151 = _5281 ^ _8423;
  wire _23152 = _23151 ^ _2291;
  wire _23153 = _23150 ^ _23152;
  wire _23154 = uncoded_block[1384] ^ uncoded_block[1389];
  wire _23155 = _23154 ^ _13412;
  wire _23156 = _7827 ^ _23155;
  wire _23157 = uncoded_block[1392] ^ uncoded_block[1394];
  wire _23158 = _23157 ^ _13938;
  wire _23159 = _6600 ^ _9016;
  wire _23160 = _23158 ^ _23159;
  wire _23161 = _23156 ^ _23160;
  wire _23162 = _23153 ^ _23161;
  wire _23163 = uncoded_block[1408] ^ uncoded_block[1412];
  wire _23164 = _23163 ^ _4583;
  wire _23165 = uncoded_block[1424] ^ uncoded_block[1429];
  wire _23166 = _7842 ^ _23165;
  wire _23167 = _23164 ^ _23166;
  wire _23168 = uncoded_block[1430] ^ uncoded_block[1434];
  wire _23169 = uncoded_block[1437] ^ uncoded_block[1441];
  wire _23170 = _23168 ^ _23169;
  wire _23171 = _3864 ^ _5976;
  wire _23172 = _23170 ^ _23171;
  wire _23173 = _23167 ^ _23172;
  wire _23174 = uncoded_block[1456] ^ uncoded_block[1459];
  wire _23175 = _6622 ^ _23174;
  wire _23176 = uncoded_block[1460] ^ uncoded_block[1467];
  wire _23177 = _23176 ^ _18919;
  wire _23178 = _23175 ^ _23177;
  wire _23179 = uncoded_block[1474] ^ uncoded_block[1477];
  wire _23180 = _11255 ^ _23179;
  wire _23181 = uncoded_block[1480] ^ uncoded_block[1484];
  wire _23182 = _23181 ^ _17489;
  wire _23183 = _23180 ^ _23182;
  wire _23184 = _23178 ^ _23183;
  wire _23185 = _23173 ^ _23184;
  wire _23186 = _23162 ^ _23185;
  wire _23187 = _23147 ^ _23186;
  wire _23188 = _23113 ^ _23187;
  wire _23189 = _11260 ^ _1571;
  wire _23190 = uncoded_block[1504] ^ uncoded_block[1509];
  wire _23191 = _23190 ^ _9053;
  wire _23192 = _23189 ^ _23191;
  wire _23193 = _751 ^ _3898;
  wire _23194 = uncoded_block[1524] ^ uncoded_block[1527];
  wire _23195 = _9059 ^ _23194;
  wire _23196 = _23193 ^ _23195;
  wire _23197 = _23192 ^ _23196;
  wire _23198 = _1582 ^ _6002;
  wire _23199 = _6005 ^ _12915;
  wire _23200 = _23198 ^ _23199;
  wire _23201 = _3128 ^ _4634;
  wire _23202 = _6013 ^ _5358;
  wire _23203 = _23201 ^ _23202;
  wire _23204 = _23200 ^ _23203;
  wire _23205 = _23197 ^ _23204;
  wire _23206 = _13991 ^ _3918;
  wire _23207 = _1598 ^ _23206;
  wire _23208 = _11838 ^ _15031;
  wire _23209 = _15028 ^ _23208;
  wire _23210 = _23207 ^ _23209;
  wire _23211 = _3146 ^ _1620;
  wire _23212 = _11847 ^ _10742;
  wire _23213 = _23211 ^ _23212;
  wire _23214 = _7906 ^ _7908;
  wire _23215 = _23214 ^ _18021;
  wire _23216 = _23213 ^ _23215;
  wire _23217 = _23210 ^ _23216;
  wire _23218 = _23205 ^ _23217;
  wire _23219 = _16524 ^ _18964;
  wire _23220 = _4667 ^ _10754;
  wire _23221 = _23220 ^ _7310;
  wire _23222 = _23219 ^ _23221;
  wire _23223 = _3169 ^ _18969;
  wire _23224 = _10757 ^ _18030;
  wire _23225 = _23223 ^ _23224;
  wire _23226 = uncoded_block[1654] ^ uncoded_block[1659];
  wire _23227 = _23226 ^ _3175;
  wire _23228 = _7319 ^ _6058;
  wire _23229 = _23227 ^ _23228;
  wire _23230 = _23225 ^ _23229;
  wire _23231 = _23222 ^ _23230;
  wire _23232 = uncoded_block[1686] ^ uncoded_block[1693];
  wire _23233 = _23232 ^ _6068;
  wire _23234 = _13518 ^ _23233;
  wire _23235 = _8535 ^ _15063;
  wire _23236 = _7335 ^ _22316;
  wire _23237 = _23235 ^ _23236;
  wire _23238 = _23234 ^ _23237;
  wire _23239 = _2441 ^ _2444;
  wire _23240 = _23239 ^ uncoded_block[1722];
  wire _23241 = _23238 ^ _23240;
  wire _23242 = _23231 ^ _23241;
  wire _23243 = _23218 ^ _23242;
  wire _23244 = _23188 ^ _23243;
  wire _23245 = _23048 ^ _23244;
  wire _23246 = _866 ^ _6724;
  wire _23247 = _868 ^ _5426;
  wire _23248 = _23246 ^ _23247;
  wire _23249 = uncoded_block[26] ^ uncoded_block[28];
  wire _23250 = _3220 ^ _23249;
  wire _23251 = _2461 ^ _18548;
  wire _23252 = _23250 ^ _23251;
  wire _23253 = _23248 ^ _23252;
  wire _23254 = _18 ^ _4723;
  wire _23255 = uncoded_block[51] ^ uncoded_block[55];
  wire _23256 = uncoded_block[56] ^ uncoded_block[59];
  wire _23257 = _23255 ^ _23256;
  wire _23258 = _23254 ^ _23257;
  wire _23259 = uncoded_block[80] ^ uncoded_block[84];
  wire _23260 = _23259 ^ _14065;
  wire _23261 = _10240 ^ _23260;
  wire _23262 = _23258 ^ _23261;
  wire _23263 = _23253 ^ _23262;
  wire _23264 = _17580 ^ _18082;
  wire _23265 = _7377 ^ _6120;
  wire _23266 = _23265 ^ _22350;
  wire _23267 = _23264 ^ _23266;
  wire _23268 = _10816 ^ _2497;
  wire _23269 = uncoded_block[120] ^ uncoded_block[123];
  wire _23270 = _23269 ^ _2502;
  wire _23271 = _23268 ^ _23270;
  wire _23272 = _924 ^ _2510;
  wire _23273 = _11918 ^ _6138;
  wire _23274 = _23272 ^ _23273;
  wire _23275 = _23271 ^ _23274;
  wire _23276 = _23267 ^ _23275;
  wire _23277 = _23263 ^ _23276;
  wire _23278 = _17097 ^ _14082;
  wire _23279 = _70 ^ _9186;
  wire _23280 = _23278 ^ _23279;
  wire _23281 = uncoded_block[156] ^ uncoded_block[159];
  wire _23282 = _23281 ^ _74;
  wire _23283 = _78 ^ _8591;
  wire _23284 = _23282 ^ _23283;
  wire _23285 = _23280 ^ _23284;
  wire _23286 = uncoded_block[172] ^ uncoded_block[182];
  wire _23287 = _23286 ^ _944;
  wire _23288 = _5483 ^ _89;
  wire _23289 = _23287 ^ _23288;
  wire _23290 = _9745 ^ _14622;
  wire _23291 = _1764 ^ _955;
  wire _23292 = _23290 ^ _23291;
  wire _23293 = _23289 ^ _23292;
  wire _23294 = _23285 ^ _23293;
  wire _23295 = _956 ^ _9750;
  wire _23296 = uncoded_block[216] ^ uncoded_block[221];
  wire _23297 = _23296 ^ _7419;
  wire _23298 = _23295 ^ _23297;
  wire _23299 = _6814 ^ _4081;
  wire _23300 = uncoded_block[232] ^ uncoded_block[236];
  wire _23301 = _23300 ^ _2552;
  wire _23302 = _23299 ^ _23301;
  wire _23303 = _23298 ^ _23302;
  wire _23304 = _116 ^ _4800;
  wire _23305 = _11953 ^ _23304;
  wire _23306 = uncoded_block[260] ^ uncoded_block[265];
  wire _23307 = _14639 ^ _23306;
  wire _23308 = _7440 ^ _3321;
  wire _23309 = _23307 ^ _23308;
  wire _23310 = _23305 ^ _23309;
  wire _23311 = _23303 ^ _23310;
  wire _23312 = _23294 ^ _23311;
  wire _23313 = _23277 ^ _23312;
  wire _23314 = _10303 ^ _12506;
  wire _23315 = _11424 ^ _11428;
  wire _23316 = _23314 ^ _23315;
  wire _23317 = _21014 ^ _8636;
  wire _23318 = _13614 ^ _23317;
  wire _23319 = _23316 ^ _23318;
  wire _23320 = _8637 ^ _17642;
  wire _23321 = _23320 ^ _11978;
  wire _23322 = _9780 ^ _11444;
  wire _23323 = _1015 ^ _15173;
  wire _23324 = _23322 ^ _23323;
  wire _23325 = _23321 ^ _23324;
  wire _23326 = _23319 ^ _23325;
  wire _23327 = _11987 ^ _159;
  wire _23328 = _23327 ^ _3360;
  wire _23329 = _6863 ^ _6227;
  wire _23330 = uncoded_block[361] ^ uncoded_block[366];
  wire _23331 = _23330 ^ _8076;
  wire _23332 = _23329 ^ _23331;
  wire _23333 = _23328 ^ _23332;
  wire _23334 = _4141 ^ _1841;
  wire _23335 = _10901 ^ _10907;
  wire _23336 = _23334 ^ _23335;
  wire _23337 = uncoded_block[390] ^ uncoded_block[397];
  wire _23338 = _23337 ^ _8087;
  wire _23339 = uncoded_block[403] ^ uncoded_block[409];
  wire _23340 = _23339 ^ _11473;
  wire _23341 = _23338 ^ _23340;
  wire _23342 = _23336 ^ _23341;
  wire _23343 = _23333 ^ _23342;
  wire _23344 = _23326 ^ _23343;
  wire _23345 = _9266 ^ _4871;
  wire _23346 = _4872 ^ _4164;
  wire _23347 = _23345 ^ _23346;
  wire _23348 = uncoded_block[432] ^ uncoded_block[437];
  wire _23349 = uncoded_block[439] ^ uncoded_block[443];
  wire _23350 = _23348 ^ _23349;
  wire _23351 = _14688 ^ _23350;
  wire _23352 = _23347 ^ _23351;
  wire _23353 = _12559 ^ _2645;
  wire _23354 = _17185 ^ _8681;
  wire _23355 = _23353 ^ _23354;
  wire _23356 = _13662 ^ _4890;
  wire _23357 = uncoded_block[466] ^ uncoded_block[469];
  wire _23358 = _23357 ^ _4188;
  wire _23359 = _23356 ^ _23358;
  wire _23360 = _23355 ^ _23359;
  wire _23361 = _23352 ^ _23360;
  wire _23362 = uncoded_block[474] ^ uncoded_block[480];
  wire _23363 = _23362 ^ _15212;
  wire _23364 = _2660 ^ _5600;
  wire _23365 = _23363 ^ _23364;
  wire _23366 = _6919 ^ _228;
  wire _23367 = _12034 ^ _17694;
  wire _23368 = _23366 ^ _23367;
  wire _23369 = _23365 ^ _23368;
  wire _23370 = uncoded_block[514] ^ uncoded_block[516];
  wire _23371 = _23370 ^ _20598;
  wire _23372 = _4919 ^ _3447;
  wire _23373 = _23371 ^ _23372;
  wire _23374 = _9850 ^ _3451;
  wire _23375 = _8132 ^ _5628;
  wire _23376 = _23374 ^ _23375;
  wire _23377 = _23373 ^ _23376;
  wire _23378 = _23369 ^ _23377;
  wire _23379 = _23361 ^ _23378;
  wire _23380 = _23344 ^ _23379;
  wire _23381 = _23313 ^ _23380;
  wire _23382 = uncoded_block[548] ^ uncoded_block[553];
  wire _23383 = _23382 ^ _1122;
  wire _23384 = _1916 ^ _10395;
  wire _23385 = _23383 ^ _23384;
  wire _23386 = _18682 ^ _4223;
  wire _23387 = uncoded_block[572] ^ uncoded_block[576];
  wire _23388 = _23387 ^ _263;
  wire _23389 = _23386 ^ _23388;
  wire _23390 = _23385 ^ _23389;
  wire _23391 = uncoded_block[584] ^ uncoded_block[590];
  wire _23392 = _9325 ^ _23391;
  wire _23393 = _2700 ^ _4952;
  wire _23394 = _23392 ^ _23393;
  wire _23395 = _9332 ^ _2710;
  wire _23396 = _4240 ^ _2713;
  wire _23397 = _23395 ^ _23396;
  wire _23398 = _23394 ^ _23397;
  wire _23399 = _23390 ^ _23398;
  wire _23400 = uncoded_block[611] ^ uncoded_block[614];
  wire _23401 = _23400 ^ _4243;
  wire _23402 = _1946 ^ _6966;
  wire _23403 = _23401 ^ _23402;
  wire _23404 = _8161 ^ _3502;
  wire _23405 = _23404 ^ _18237;
  wire _23406 = _23403 ^ _23405;
  wire _23407 = _8166 ^ _2738;
  wire _23408 = _308 ^ _13190;
  wire _23409 = _23407 ^ _23408;
  wire _23410 = uncoded_block[676] ^ uncoded_block[679];
  wire _23411 = _16752 ^ _23410;
  wire _23412 = uncoded_block[680] ^ uncoded_block[684];
  wire _23413 = _23412 ^ _3527;
  wire _23414 = _23411 ^ _23413;
  wire _23415 = _23409 ^ _23414;
  wire _23416 = _23406 ^ _23415;
  wire _23417 = _23399 ^ _23416;
  wire _23418 = _6985 ^ _9896;
  wire _23419 = _3535 ^ _337;
  wire _23420 = _23418 ^ _23419;
  wire _23421 = _9902 ^ _6374;
  wire _23422 = _5693 ^ _8200;
  wire _23423 = _23421 ^ _23422;
  wire _23424 = _23420 ^ _23423;
  wire _23425 = uncoded_block[736] ^ uncoded_block[738];
  wire _23426 = _8201 ^ _23425;
  wire _23427 = _1207 ^ _10464;
  wire _23428 = _23426 ^ _23427;
  wire _23429 = _16775 ^ _7013;
  wire _23430 = _7015 ^ _3559;
  wire _23431 = _23429 ^ _23430;
  wire _23432 = _23428 ^ _23431;
  wire _23433 = _23424 ^ _23432;
  wire _23434 = _12113 ^ _2012;
  wire _23435 = _366 ^ _23434;
  wire _23436 = _2014 ^ _2794;
  wire _23437 = _4309 ^ _5032;
  wire _23438 = _23436 ^ _23437;
  wire _23439 = _23435 ^ _23438;
  wire _23440 = _8223 ^ _16790;
  wire _23441 = _3575 ^ _23440;
  wire _23442 = uncoded_block[805] ^ uncoded_block[810];
  wire _23443 = _23442 ^ _2026;
  wire _23444 = _6398 ^ _15320;
  wire _23445 = _23443 ^ _23444;
  wire _23446 = _23441 ^ _23445;
  wire _23447 = _23439 ^ _23446;
  wire _23448 = _23433 ^ _23447;
  wire _23449 = _23417 ^ _23448;
  wire _23450 = uncoded_block[824] ^ uncoded_block[826];
  wire _23451 = _23450 ^ _10490;
  wire _23452 = _1250 ^ _2035;
  wire _23453 = _23451 ^ _23452;
  wire _23454 = uncoded_block[843] ^ uncoded_block[848];
  wire _23455 = _5737 ^ _23454;
  wire _23456 = _2044 ^ _8237;
  wire _23457 = _23455 ^ _23456;
  wire _23458 = _23453 ^ _23457;
  wire _23459 = _8812 ^ _15824;
  wire _23460 = _5069 ^ _5749;
  wire _23461 = _23459 ^ _23460;
  wire _23462 = uncoded_block[879] ^ uncoded_block[884];
  wire _23463 = _11620 ^ _23462;
  wire _23464 = uncoded_block[885] ^ uncoded_block[889];
  wire _23465 = _23464 ^ _5085;
  wire _23466 = _23463 ^ _23465;
  wire _23467 = _23461 ^ _23466;
  wire _23468 = _23458 ^ _23467;
  wire _23469 = _8826 ^ _3623;
  wire _23470 = _23469 ^ _15349;
  wire _23471 = uncoded_block[921] ^ uncoded_block[925];
  wire _23472 = _23471 ^ _18316;
  wire _23473 = _12713 ^ _23472;
  wire _23474 = _23470 ^ _23473;
  wire _23475 = uncoded_block[933] ^ uncoded_block[938];
  wire _23476 = _23475 ^ _12723;
  wire _23477 = _12725 ^ _1303;
  wire _23478 = _23476 ^ _23477;
  wire _23479 = _8275 ^ _9979;
  wire _23480 = _5783 ^ _7088;
  wire _23481 = _23479 ^ _23480;
  wire _23482 = _23478 ^ _23481;
  wire _23483 = _23474 ^ _23482;
  wire _23484 = _23468 ^ _23483;
  wire _23485 = _20219 ^ _5789;
  wire _23486 = _476 ^ _12734;
  wire _23487 = _23485 ^ _23486;
  wire _23488 = _6453 ^ _4404;
  wire _23489 = _484 ^ _4405;
  wire _23490 = _23488 ^ _23489;
  wire _23491 = _23487 ^ _23490;
  wire _23492 = _4409 ^ _1331;
  wire _23493 = _492 ^ _5137;
  wire _23494 = _23492 ^ _23493;
  wire _23495 = _8302 ^ _8305;
  wire _23496 = _23494 ^ _23495;
  wire _23497 = _23491 ^ _23496;
  wire _23498 = uncoded_block[1041] ^ uncoded_block[1045];
  wire _23499 = _23498 ^ _2913;
  wire _23500 = _5144 ^ _23499;
  wire _23501 = _2136 ^ _9465;
  wire _23502 = _522 ^ _8888;
  wire _23503 = _23501 ^ _23502;
  wire _23504 = _23500 ^ _23503;
  wire _23505 = uncoded_block[1068] ^ uncoded_block[1077];
  wire _23506 = uncoded_block[1078] ^ uncoded_block[1087];
  wire _23507 = _23505 ^ _23506;
  wire _23508 = uncoded_block[1091] ^ uncoded_block[1094];
  wire _23509 = _4440 ^ _23508;
  wire _23510 = _23507 ^ _23509;
  wire _23511 = _1380 ^ _19794;
  wire _23512 = _8336 ^ _4450;
  wire _23513 = _23511 ^ _23512;
  wire _23514 = _23510 ^ _23513;
  wire _23515 = _23504 ^ _23514;
  wire _23516 = _23497 ^ _23515;
  wire _23517 = _23484 ^ _23516;
  wire _23518 = _23449 ^ _23517;
  wire _23519 = _23381 ^ _23518;
  wire _23520 = _8917 ^ _5175;
  wire _23521 = _16376 ^ _5854;
  wire _23522 = _23520 ^ _23521;
  wire _23523 = uncoded_block[1127] ^ uncoded_block[1129];
  wire _23524 = _23523 ^ _1393;
  wire _23525 = uncoded_block[1136] ^ uncoded_block[1141];
  wire _23526 = _10591 ^ _23525;
  wire _23527 = _23524 ^ _23526;
  wire _23528 = _23522 ^ _23527;
  wire _23529 = _568 ^ _8932;
  wire _23530 = _4465 ^ _2185;
  wire _23531 = _23529 ^ _23530;
  wire _23532 = uncoded_block[1162] ^ uncoded_block[1167];
  wire _23533 = _23532 ^ _10046;
  wire _23534 = _5191 ^ _23533;
  wire _23535 = _23531 ^ _23534;
  wire _23536 = _23528 ^ _23535;
  wire _23537 = _4482 ^ _16901;
  wire _23538 = _5201 ^ _2971;
  wire _23539 = _23537 ^ _23538;
  wire _23540 = _17898 ^ _11721;
  wire _23541 = _8370 ^ _16399;
  wire _23542 = _23540 ^ _23541;
  wire _23543 = _23539 ^ _23542;
  wire _23544 = uncoded_block[1208] ^ uncoded_block[1210];
  wire _23545 = _23544 ^ _12813;
  wire _23546 = _2220 ^ _4502;
  wire _23547 = _23545 ^ _23546;
  wire _23548 = uncoded_block[1230] ^ uncoded_block[1235];
  wire _23549 = _609 ^ _23548;
  wire _23550 = uncoded_block[1241] ^ uncoded_block[1245];
  wire _23551 = _23550 ^ _1449;
  wire _23552 = _23549 ^ _23551;
  wire _23553 = _23547 ^ _23552;
  wire _23554 = _23543 ^ _23553;
  wire _23555 = _23536 ^ _23554;
  wire _23556 = _3779 ^ _8388;
  wire _23557 = _3783 ^ _7781;
  wire _23558 = _23556 ^ _23557;
  wire _23559 = uncoded_block[1266] ^ uncoded_block[1270];
  wire _23560 = _23559 ^ _628;
  wire _23561 = _3005 ^ _23560;
  wire _23562 = _23558 ^ _23561;
  wire _23563 = _16419 ^ _7792;
  wire _23564 = _23563 ^ _13911;
  wire _23565 = _3800 ^ _9547;
  wire _23566 = _16421 ^ _23565;
  wire _23567 = _23564 ^ _23566;
  wire _23568 = _23562 ^ _23567;
  wire _23569 = _18870 ^ _22665;
  wire _23570 = _8991 ^ _6572;
  wire _23571 = _23569 ^ _23570;
  wire _23572 = _20314 ^ _9552;
  wire _23573 = _19375 ^ _4545;
  wire _23574 = _23572 ^ _23573;
  wire _23575 = _23571 ^ _23574;
  wire _23576 = uncoded_block[1336] ^ uncoded_block[1339];
  wire _23577 = _5256 ^ _23576;
  wire _23578 = _1497 ^ _14950;
  wire _23579 = _23577 ^ _23578;
  wire _23580 = _11771 ^ _18434;
  wire _23581 = uncoded_block[1357] ^ uncoded_block[1359];
  wire _23582 = _18436 ^ _23581;
  wire _23583 = _23580 ^ _23582;
  wire _23584 = _23579 ^ _23583;
  wire _23585 = _23575 ^ _23584;
  wire _23586 = _23568 ^ _23585;
  wire _23587 = _23555 ^ _23586;
  wire _23588 = _16444 ^ _679;
  wire _23589 = uncoded_block[1374] ^ uncoded_block[1377];
  wire _23590 = _17945 ^ _23589;
  wire _23591 = _23588 ^ _23590;
  wire _23592 = _2290 ^ _7219;
  wire _23593 = _3059 ^ _12311;
  wire _23594 = _23592 ^ _23593;
  wire _23595 = _23591 ^ _23594;
  wire _23596 = _1513 ^ _4568;
  wire _23597 = _23596 ^ _9015;
  wire _23598 = _695 ^ _14968;
  wire _23599 = _9585 ^ _12877;
  wire _23600 = _23598 ^ _23599;
  wire _23601 = _23597 ^ _23600;
  wire _23602 = _23595 ^ _23601;
  wire _23603 = _2306 ^ _11792;
  wire _23604 = uncoded_block[1427] ^ uncoded_block[1430];
  wire _23605 = _9588 ^ _23604;
  wire _23606 = _23603 ^ _23605;
  wire _23607 = _9591 ^ _9595;
  wire _23608 = uncoded_block[1441] ^ uncoded_block[1448];
  wire _23609 = _23608 ^ _5976;
  wire _23610 = _23607 ^ _23609;
  wire _23611 = _23606 ^ _23610;
  wire _23612 = _726 ^ _8455;
  wire _23613 = _23175 ^ _23612;
  wire _23614 = uncoded_block[1468] ^ uncoded_block[1472];
  wire _23615 = _10136 ^ _23614;
  wire _23616 = _4603 ^ _3100;
  wire _23617 = _23615 ^ _23616;
  wire _23618 = _23613 ^ _23617;
  wire _23619 = _23611 ^ _23618;
  wire _23620 = _23602 ^ _23619;
  wire _23621 = _22711 ^ _740;
  wire _23622 = _17489 ^ _12896;
  wire _23623 = _23621 ^ _23622;
  wire _23624 = uncoded_block[1507] ^ uncoded_block[1510];
  wire _23625 = _18478 ^ _23624;
  wire _23626 = _12345 ^ _23625;
  wire _23627 = _23623 ^ _23626;
  wire _23628 = _1575 ^ _1578;
  wire _23629 = uncoded_block[1524] ^ uncoded_block[1528];
  wire _23630 = _9059 ^ _23629;
  wire _23631 = _23628 ^ _23630;
  wire _23632 = _3125 ^ _6648;
  wire _23633 = _2365 ^ _3129;
  wire _23634 = _23632 ^ _23633;
  wire _23635 = _23631 ^ _23634;
  wire _23636 = _23627 ^ _23635;
  wire _23637 = _9067 ^ _6657;
  wire _23638 = _9070 ^ _3914;
  wire _23639 = _23637 ^ _23638;
  wire _23640 = uncoded_block[1561] ^ uncoded_block[1564];
  wire _23641 = _23640 ^ _16510;
  wire _23642 = _14506 ^ _1609;
  wire _23643 = _23641 ^ _23642;
  wire _23644 = _23639 ^ _23643;
  wire _23645 = _17009 ^ _3145;
  wire _23646 = _14512 ^ _4654;
  wire _23647 = _23645 ^ _23646;
  wire _23648 = uncoded_block[1597] ^ uncoded_block[1602];
  wire _23649 = _23648 ^ _8502;
  wire _23650 = _23649 ^ _2399;
  wire _23651 = _23647 ^ _23650;
  wire _23652 = _23644 ^ _23651;
  wire _23653 = _23636 ^ _23652;
  wire _23654 = _23620 ^ _23653;
  wire _23655 = _23587 ^ _23654;
  wire _23656 = _18021 ^ _18024;
  wire _23657 = _14525 ^ _4667;
  wire _23658 = uncoded_block[1632] ^ uncoded_block[1634];
  wire _23659 = _23658 ^ _7309;
  wire _23660 = _23657 ^ _23659;
  wire _23661 = _23656 ^ _23660;
  wire _23662 = _4673 ^ _2412;
  wire _23663 = _23662 ^ _19936;
  wire _23664 = _3174 ^ _10196;
  wire _23665 = uncoded_block[1667] ^ uncoded_block[1673];
  wire _23666 = _17032 ^ _23665;
  wire _23667 = _23664 ^ _23666;
  wire _23668 = _23663 ^ _23667;
  wire _23669 = _23661 ^ _23668;
  wire _23670 = _3183 ^ _20427;
  wire _23671 = uncoded_block[1681] ^ uncoded_block[1684];
  wire _23672 = _23671 ^ _14543;
  wire _23673 = _23670 ^ _23672;
  wire _23674 = _3968 ^ _21394;
  wire _23675 = _9671 ^ _23674;
  wire _23676 = _23673 ^ _23675;
  wire _23677 = _15063 ^ _3200;
  wire _23678 = _17545 ^ _23677;
  wire _23679 = _14552 ^ _3988;
  wire _23680 = _23679 ^ uncoded_block[1720];
  wire _23681 = _23678 ^ _23680;
  wire _23682 = _23676 ^ _23681;
  wire _23683 = _23669 ^ _23682;
  wire _23684 = _23655 ^ _23683;
  wire _23685 = _23519 ^ _23684;
  wire _23686 = _4712 ^ _4;
  wire _23687 = _2 ^ _23686;
  wire _23688 = uncoded_block[12] ^ uncoded_block[19];
  wire _23689 = _23688 ^ _1690;
  wire _23690 = _5427 ^ _9144;
  wire _23691 = _23689 ^ _23690;
  wire _23692 = _23687 ^ _23691;
  wire _23693 = uncoded_block[36] ^ uncoded_block[40];
  wire _23694 = _16 ^ _23693;
  wire _23695 = _23694 ^ _21873;
  wire _23696 = _3232 ^ _1700;
  wire _23697 = uncoded_block[55] ^ uncoded_block[60];
  wire _23698 = uncoded_block[62] ^ uncoded_block[65];
  wire _23699 = _23697 ^ _23698;
  wire _23700 = _23696 ^ _23699;
  wire _23701 = _23695 ^ _23700;
  wire _23702 = _23692 ^ _23701;
  wire _23703 = _11357 ^ _10244;
  wire _23704 = _39 ^ _6750;
  wire _23705 = _23703 ^ _23704;
  wire _23706 = uncoded_block[86] ^ uncoded_block[91];
  wire _23707 = _23706 ^ _8567;
  wire _23708 = _14068 ^ _4745;
  wire _23709 = _23707 ^ _23708;
  wire _23710 = _23705 ^ _23709;
  wire _23711 = _49 ^ _13011;
  wire _23712 = _5453 ^ _915;
  wire _23713 = _23711 ^ _23712;
  wire _23714 = _4750 ^ _12451;
  wire _23715 = _917 ^ _923;
  wire _23716 = _23714 ^ _23715;
  wire _23717 = _23713 ^ _23716;
  wire _23718 = _23710 ^ _23717;
  wire _23719 = _23702 ^ _23718;
  wire _23720 = uncoded_block[133] ^ uncoded_block[138];
  wire _23721 = _23720 ^ _15114;
  wire _23722 = uncoded_block[146] ^ uncoded_block[150];
  wire _23723 = _7392 ^ _23722;
  wire _23724 = _23721 ^ _23723;
  wire _23725 = _15623 ^ _1748;
  wire _23726 = _15118 ^ _74;
  wire _23727 = _23725 ^ _23726;
  wire _23728 = _23724 ^ _23727;
  wire _23729 = uncoded_block[170] ^ uncoded_block[173];
  wire _23730 = _23729 ^ _1756;
  wire _23731 = _13580 ^ _23730;
  wire _23732 = _18110 ^ _22368;
  wire _23733 = _89 ^ _10277;
  wire _23734 = _23732 ^ _23733;
  wire _23735 = _23731 ^ _23734;
  wire _23736 = _23728 ^ _23735;
  wire _23737 = _15135 ^ _3289;
  wire _23738 = _23737 ^ _18117;
  wire _23739 = uncoded_block[222] ^ uncoded_block[226];
  wire _23740 = _4787 ^ _23739;
  wire _23741 = uncoded_block[227] ^ uncoded_block[235];
  wire _23742 = _23741 ^ _5500;
  wire _23743 = _23740 ^ _23742;
  wire _23744 = _23738 ^ _23743;
  wire _23745 = _8032 ^ _3309;
  wire _23746 = uncoded_block[255] ^ uncoded_block[257];
  wire _23747 = _23746 ^ _1788;
  wire _23748 = _23745 ^ _23747;
  wire _23749 = _120 ^ _20523;
  wire _23750 = uncoded_block[271] ^ uncoded_block[281];
  wire _23751 = _14642 ^ _23750;
  wire _23752 = _23749 ^ _23751;
  wire _23753 = _23748 ^ _23752;
  wire _23754 = _23744 ^ _23753;
  wire _23755 = _23736 ^ _23754;
  wire _23756 = _23719 ^ _23755;
  wire _23757 = _1803 ^ _6837;
  wire _23758 = _10876 ^ _4819;
  wire _23759 = _23757 ^ _23758;
  wire _23760 = uncoded_block[294] ^ uncoded_block[299];
  wire _23761 = _23760 ^ _17144;
  wire _23762 = _23761 ^ _10314;
  wire _23763 = _23759 ^ _23762;
  wire _23764 = uncoded_block[313] ^ uncoded_block[316];
  wire _23765 = _21017 ^ _23764;
  wire _23766 = _23765 ^ _15676;
  wire _23767 = _3346 ^ _9780;
  wire _23768 = _6853 ^ _13629;
  wire _23769 = _23767 ^ _23768;
  wire _23770 = _23766 ^ _23769;
  wire _23771 = _23763 ^ _23770;
  wire _23772 = _3356 ^ _16657;
  wire _23773 = _19092 ^ _3361;
  wire _23774 = _6866 ^ _15183;
  wire _23775 = _23773 ^ _23774;
  wire _23776 = _23772 ^ _23775;
  wire _23777 = uncoded_block[376] ^ uncoded_block[383];
  wire _23778 = _169 ^ _23777;
  wire _23779 = uncoded_block[387] ^ uncoded_block[390];
  wire _23780 = _23779 ^ _19604;
  wire _23781 = _23778 ^ _23780;
  wire _23782 = _3384 ^ _2622;
  wire _23783 = _10341 ^ _1051;
  wire _23784 = _23782 ^ _23783;
  wire _23785 = _23781 ^ _23784;
  wire _23786 = _23776 ^ _23785;
  wire _23787 = _23771 ^ _23786;
  wire _23788 = uncoded_block[415] ^ uncoded_block[418];
  wire _23789 = _1052 ^ _23788;
  wire _23790 = _4872 ^ _12551;
  wire _23791 = _23789 ^ _23790;
  wire _23792 = _13115 ^ _1857;
  wire _23793 = uncoded_block[435] ^ uncoded_block[441];
  wire _23794 = _23793 ^ _5580;
  wire _23795 = _23792 ^ _23794;
  wire _23796 = _23791 ^ _23795;
  wire _23797 = _1070 ^ _1076;
  wire _23798 = _8681 ^ _1873;
  wire _23799 = _23797 ^ _23798;
  wire _23800 = uncoded_block[467] ^ uncoded_block[470];
  wire _23801 = _8683 ^ _23800;
  wire _23802 = _221 ^ _8110;
  wire _23803 = _23801 ^ _23802;
  wire _23804 = _23799 ^ _23803;
  wire _23805 = _23796 ^ _23804;
  wire _23806 = _21528 ^ _6276;
  wire _23807 = uncoded_block[495] ^ uncoded_block[500];
  wire _23808 = _10937 ^ _23807;
  wire _23809 = _23806 ^ _23808;
  wire _23810 = _19135 ^ _1892;
  wire _23811 = uncoded_block[514] ^ uncoded_block[522];
  wire _23812 = _9295 ^ _23811;
  wire _23813 = _23810 ^ _23812;
  wire _23814 = _23809 ^ _23813;
  wire _23815 = _6290 ^ _1114;
  wire _23816 = _15228 ^ _23815;
  wire _23817 = _6293 ^ _9854;
  wire _23818 = _1117 ^ _4931;
  wire _23819 = _23817 ^ _23818;
  wire _23820 = _23816 ^ _23819;
  wire _23821 = _23814 ^ _23820;
  wire _23822 = _23805 ^ _23821;
  wire _23823 = _23787 ^ _23822;
  wire _23824 = _23756 ^ _23823;
  wire _23825 = _4933 ^ _3459;
  wire _23826 = uncoded_block[559] ^ uncoded_block[563];
  wire _23827 = _14204 ^ _23826;
  wire _23828 = _23825 ^ _23827;
  wire _23829 = uncoded_block[567] ^ uncoded_block[571];
  wire _23830 = _3465 ^ _23829;
  wire _23831 = _4224 ^ _1931;
  wire _23832 = _23830 ^ _23831;
  wire _23833 = _23828 ^ _23832;
  wire _23834 = _15747 ^ _1933;
  wire _23835 = uncoded_block[590] ^ uncoded_block[594];
  wire _23836 = _1934 ^ _23835;
  wire _23837 = _23834 ^ _23836;
  wire _23838 = _6952 ^ _1142;
  wire _23839 = _23838 ^ _2711;
  wire _23840 = _23837 ^ _23839;
  wire _23841 = _23833 ^ _23840;
  wire _23842 = uncoded_block[609] ^ uncoded_block[614];
  wire _23843 = _277 ^ _23842;
  wire _23844 = _5653 ^ _4960;
  wire _23845 = _23843 ^ _23844;
  wire _23846 = uncoded_block[624] ^ uncoded_block[633];
  wire _23847 = _23846 ^ _13717;
  wire _23848 = _16241 ^ _3505;
  wire _23849 = _23847 ^ _23848;
  wire _23850 = _23845 ^ _23849;
  wire _23851 = _16247 ^ _4975;
  wire _23852 = _14755 ^ _4261;
  wire _23853 = _23851 ^ _23852;
  wire _23854 = uncoded_block[670] ^ uncoded_block[674];
  wire _23855 = _2742 ^ _23854;
  wire _23856 = uncoded_block[681] ^ uncoded_block[688];
  wire _23857 = _12634 ^ _23856;
  wire _23858 = _23855 ^ _23857;
  wire _23859 = _23853 ^ _23858;
  wire _23860 = _23850 ^ _23859;
  wire _23861 = _23841 ^ _23860;
  wire _23862 = _21121 ^ _330;
  wire _23863 = uncoded_block[707] ^ uncoded_block[709];
  wire _23864 = _23863 ^ _2762;
  wire _23865 = _15286 ^ _23864;
  wire _23866 = _23862 ^ _23865;
  wire _23867 = uncoded_block[713] ^ uncoded_block[719];
  wire _23868 = _23867 ^ _12648;
  wire _23869 = _23868 ^ _3545;
  wire _23870 = uncoded_block[739] ^ uncoded_block[740];
  wire _23871 = _23870 ^ _2774;
  wire _23872 = _21599 ^ _23871;
  wire _23873 = _23869 ^ _23872;
  wire _23874 = _23866 ^ _23873;
  wire _23875 = _5012 ^ _4293;
  wire _23876 = uncoded_block[752] ^ uncoded_block[754];
  wire _23877 = _23876 ^ _2778;
  wire _23878 = _23875 ^ _23877;
  wire _23879 = uncoded_block[758] ^ uncoded_block[760];
  wire _23880 = _23879 ^ _13761;
  wire _23881 = _11018 ^ _5027;
  wire _23882 = _23880 ^ _23881;
  wire _23883 = _23878 ^ _23882;
  wire _23884 = _6382 ^ _13766;
  wire _23885 = _3568 ^ _4311;
  wire _23886 = _23884 ^ _23885;
  wire _23887 = _2019 ^ _1233;
  wire _23888 = _383 ^ _4317;
  wire _23889 = _23887 ^ _23888;
  wire _23890 = _23886 ^ _23889;
  wire _23891 = _23883 ^ _23890;
  wire _23892 = _23874 ^ _23891;
  wire _23893 = _23861 ^ _23892;
  wire _23894 = _11596 ^ _1241;
  wire _23895 = _19227 ^ _23894;
  wire _23896 = uncoded_block[826] ^ uncoded_block[829];
  wire _23897 = _11600 ^ _23896;
  wire _23898 = _10490 ^ _401;
  wire _23899 = _23897 ^ _23898;
  wire _23900 = _23895 ^ _23899;
  wire _23901 = uncoded_block[837] ^ uncoded_block[846];
  wire _23902 = _23901 ^ _4340;
  wire _23903 = _11048 ^ _3600;
  wire _23904 = _23902 ^ _23903;
  wire _23905 = _14300 ^ _2824;
  wire _23906 = uncoded_block[874] ^ uncoded_block[877];
  wire _23907 = _8243 ^ _23906;
  wire _23908 = _23905 ^ _23907;
  wire _23909 = _23904 ^ _23908;
  wire _23910 = _23900 ^ _23909;
  wire _23911 = _23464 ^ _2061;
  wire _23912 = _23911 ^ _15834;
  wire _23913 = _8250 ^ _429;
  wire _23914 = _23913 ^ _1282;
  wire _23915 = _23912 ^ _23914;
  wire _23916 = _1284 ^ _14317;
  wire _23917 = uncoded_block[916] ^ uncoded_block[918];
  wire _23918 = _23917 ^ _445;
  wire _23919 = _23916 ^ _23918;
  wire _23920 = _2857 ^ _21649;
  wire _23921 = _453 ^ _8271;
  wire _23922 = _23920 ^ _23921;
  wire _23923 = _23919 ^ _23922;
  wire _23924 = _23915 ^ _23923;
  wire _23925 = _23910 ^ _23924;
  wire _23926 = uncoded_block[946] ^ uncoded_block[948];
  wire _23927 = _23926 ^ _21191;
  wire _23928 = _8275 ^ _4384;
  wire _23929 = _23927 ^ _23928;
  wire _23930 = _8277 ^ _5107;
  wire _23931 = _14844 ^ _11087;
  wire _23932 = _23930 ^ _23931;
  wire _23933 = _23929 ^ _23932;
  wire _23934 = uncoded_block[974] ^ uncoded_block[978];
  wire _23935 = _2877 ^ _23934;
  wire _23936 = _12733 ^ _6451;
  wire _23937 = _23935 ^ _23936;
  wire _23938 = uncoded_block[988] ^ uncoded_block[989];
  wire _23939 = uncoded_block[990] ^ uncoded_block[992];
  wire _23940 = _23938 ^ _23939;
  wire _23941 = _10543 ^ _6453;
  wire _23942 = _23940 ^ _23941;
  wire _23943 = _23937 ^ _23942;
  wire _23944 = _23933 ^ _23943;
  wire _23945 = uncoded_block[999] ^ uncoded_block[1001];
  wire _23946 = _11101 ^ _23945;
  wire _23947 = _4404 ^ _2114;
  wire _23948 = _23946 ^ _23947;
  wire _23949 = _1330 ^ _2117;
  wire _23950 = _2893 ^ _7108;
  wire _23951 = _23949 ^ _23950;
  wire _23952 = _23948 ^ _23951;
  wire _23953 = _1338 ^ _18801;
  wire _23954 = _23953 ^ _8305;
  wire _23955 = _7707 ^ _3678;
  wire _23956 = _2130 ^ _2133;
  wire _23957 = _23955 ^ _23956;
  wire _23958 = _23954 ^ _23957;
  wire _23959 = _23952 ^ _23958;
  wire _23960 = _23944 ^ _23959;
  wire _23961 = _23925 ^ _23960;
  wire _23962 = _23893 ^ _23961;
  wire _23963 = _23824 ^ _23962;
  wire _23964 = uncoded_block[1047] ^ uncoded_block[1049];
  wire _23965 = _23964 ^ _7714;
  wire _23966 = uncoded_block[1054] ^ uncoded_block[1057];
  wire _23967 = _23966 ^ _6483;
  wire _23968 = _23965 ^ _23967;
  wire _23969 = uncoded_block[1066] ^ uncoded_block[1069];
  wire _23970 = _23969 ^ _2924;
  wire _23971 = _8895 ^ _5163;
  wire _23972 = _23970 ^ _23971;
  wire _23973 = _23968 ^ _23972;
  wire _23974 = _534 ^ _5840;
  wire _23975 = _23974 ^ _5844;
  wire _23976 = _3707 ^ _549;
  wire _23977 = _23976 ^ _4452;
  wire _23978 = _23975 ^ _23977;
  wire _23979 = _23973 ^ _23978;
  wire _23980 = _19313 ^ _2168;
  wire _23981 = uncoded_block[1129] ^ uncoded_block[1132];
  wire _23982 = _13327 ^ _23981;
  wire _23983 = _23980 ^ _23982;
  wire _23984 = _5859 ^ _10597;
  wire _23985 = _15897 ^ _23984;
  wire _23986 = _23983 ^ _23985;
  wire _23987 = _6505 ^ _17386;
  wire _23988 = _8356 ^ _6511;
  wire _23989 = _23987 ^ _23988;
  wire _23990 = _5193 ^ _17392;
  wire _23991 = _5872 ^ _590;
  wire _23992 = _23990 ^ _23991;
  wire _23993 = _23989 ^ _23992;
  wire _23994 = _23986 ^ _23993;
  wire _23995 = _23979 ^ _23994;
  wire _23996 = uncoded_block[1187] ^ uncoded_block[1189];
  wire _23997 = _13882 ^ _23996;
  wire _23998 = _23997 ^ _7757;
  wire _23999 = uncoded_block[1197] ^ uncoded_block[1200];
  wire _24000 = _23999 ^ _11722;
  wire _24001 = uncoded_block[1208] ^ uncoded_block[1211];
  wire _24002 = _24001 ^ _4502;
  wire _24003 = _24000 ^ _24002;
  wire _24004 = _23998 ^ _24003;
  wire _24005 = _8958 ^ _612;
  wire _24006 = _13357 ^ _15927;
  wire _24007 = _24005 ^ _24006;
  wire _24008 = uncoded_block[1244] ^ uncoded_block[1249];
  wire _24009 = _2230 ^ _24008;
  wire _24010 = uncoded_block[1250] ^ uncoded_block[1254];
  wire _24011 = _24010 ^ _7780;
  wire _24012 = _24009 ^ _24011;
  wire _24013 = _24007 ^ _24012;
  wire _24014 = _24004 ^ _24013;
  wire _24015 = _7781 ^ _3003;
  wire _24016 = _3004 ^ _627;
  wire _24017 = _24015 ^ _24016;
  wire _24018 = uncoded_block[1267] ^ uncoded_block[1274];
  wire _24019 = _24018 ^ _5908;
  wire _24020 = _631 ^ _12837;
  wire _24021 = _24019 ^ _24020;
  wire _24022 = _24017 ^ _24021;
  wire _24023 = uncoded_block[1285] ^ uncoded_block[1287];
  wire _24024 = _24023 ^ _13380;
  wire _24025 = _24024 ^ _1470;
  wire _24026 = _9547 ^ _4532;
  wire _24027 = _8984 ^ _3025;
  wire _24028 = _24026 ^ _24027;
  wire _24029 = _24025 ^ _24028;
  wire _24030 = _24022 ^ _24029;
  wire _24031 = _24014 ^ _24030;
  wire _24032 = _23995 ^ _24031;
  wire _24033 = _1480 ^ _1482;
  wire _24034 = _24033 ^ _14944;
  wire _24035 = _4543 ^ _11764;
  wire _24036 = uncoded_block[1334] ^ uncoded_block[1337];
  wire _24037 = _5931 ^ _24036;
  wire _24038 = _24035 ^ _24037;
  wire _24039 = _24034 ^ _24038;
  wire _24040 = uncoded_block[1346] ^ uncoded_block[1350];
  wire _24041 = _24040 ^ _3042;
  wire _24042 = _5934 ^ _24041;
  wire _24043 = _5940 ^ _12300;
  wire _24044 = _2283 ^ _14960;
  wire _24045 = _24043 ^ _24044;
  wire _24046 = _24042 ^ _24045;
  wire _24047 = _24039 ^ _24046;
  wire _24048 = _5284 ^ _2290;
  wire _24049 = _16451 ^ _3061;
  wire _24050 = _24048 ^ _24049;
  wire _24051 = _11782 ^ _13412;
  wire _24052 = _7834 ^ _2297;
  wire _24053 = _24051 ^ _24052;
  wire _24054 = _24050 ^ _24053;
  wire _24055 = _2299 ^ _3849;
  wire _24056 = _10681 ^ _705;
  wire _24057 = _24055 ^ _24056;
  wire _24058 = uncoded_block[1423] ^ uncoded_block[1426];
  wire _24059 = _13428 ^ _24058;
  wire _24060 = _10684 ^ _10690;
  wire _24061 = _24059 ^ _24060;
  wire _24062 = _24057 ^ _24061;
  wire _24063 = _24054 ^ _24062;
  wire _24064 = _24047 ^ _24063;
  wire _24065 = uncoded_block[1439] ^ uncoded_block[1441];
  wire _24066 = _24065 ^ _716;
  wire _24067 = _2322 ^ _6620;
  wire _24068 = _24066 ^ _24067;
  wire _24069 = _6622 ^ _11249;
  wire _24070 = uncoded_block[1462] ^ uncoded_block[1465];
  wire _24071 = uncoded_block[1467] ^ uncoded_block[1470];
  wire _24072 = _24070 ^ _24071;
  wire _24073 = _24069 ^ _24072;
  wire _24074 = _24068 ^ _24073;
  wire _24075 = _10701 ^ _3884;
  wire _24076 = _739 ^ _13966;
  wire _24077 = _24075 ^ _24076;
  wire _24078 = uncoded_block[1494] ^ uncoded_block[1496];
  wire _24079 = _1565 ^ _24078;
  wire _24080 = _2352 ^ _7258;
  wire _24081 = _24079 ^ _24080;
  wire _24082 = _24077 ^ _24081;
  wire _24083 = _24074 ^ _24082;
  wire _24084 = uncoded_block[1503] ^ uncoded_block[1506];
  wire _24085 = _24084 ^ _5333;
  wire _24086 = _24085 ^ _9622;
  wire _24087 = _22723 ^ _17499;
  wire _24088 = _4624 ^ _5347;
  wire _24089 = _24087 ^ _24088;
  wire _24090 = _24086 ^ _24089;
  wire _24091 = _5348 ^ _5350;
  wire _24092 = _5355 ^ _7275;
  wire _24093 = _24091 ^ _24092;
  wire _24094 = uncoded_block[1556] ^ uncoded_block[1559];
  wire _24095 = _24094 ^ _13991;
  wire _24096 = _14497 ^ _24095;
  wire _24097 = _24093 ^ _24096;
  wire _24098 = _24090 ^ _24097;
  wire _24099 = _24083 ^ _24098;
  wire _24100 = _24064 ^ _24099;
  wire _24101 = _24032 ^ _24100;
  wire _24102 = uncoded_block[1565] ^ uncoded_block[1570];
  wire _24103 = uncoded_block[1574] ^ uncoded_block[1577];
  wire _24104 = _24102 ^ _24103;
  wire _24105 = _13479 ^ _1612;
  wire _24106 = _24104 ^ _24105;
  wire _24107 = _10172 ^ _4653;
  wire _24108 = _21827 ^ _11295;
  wire _24109 = _24107 ^ _24108;
  wire _24110 = _24106 ^ _24109;
  wire _24111 = _3151 ^ _20406;
  wire _24112 = _2396 ^ _4662;
  wire _24113 = _24111 ^ _24112;
  wire _24114 = _7908 ^ _10181;
  wire _24115 = uncoded_block[1617] ^ uncoded_block[1620];
  wire _24116 = _24115 ^ _7300;
  wire _24117 = _24114 ^ _24116;
  wire _24118 = _24113 ^ _24117;
  wire _24119 = _24110 ^ _24118;
  wire _24120 = _12947 ^ _4667;
  wire _24121 = _5388 ^ _7914;
  wire _24122 = _24120 ^ _24121;
  wire _24123 = _7306 ^ _12383;
  wire _24124 = _24123 ^ _13507;
  wire _24125 = _24122 ^ _24124;
  wire _24126 = _12390 ^ _3958;
  wire _24127 = _19939 ^ _6700;
  wire _24128 = _24126 ^ _24127;
  wire _24129 = _11319 ^ _7933;
  wire _24130 = uncoded_block[1686] ^ uncoded_block[1687];
  wire _24131 = _24130 ^ _11325;
  wire _24132 = _24129 ^ _24131;
  wire _24133 = _24128 ^ _24132;
  wire _24134 = _24125 ^ _24133;
  wire _24135 = _24119 ^ _24134;
  wire _24136 = _21394 ^ _11327;
  wire _24137 = uncoded_block[1701] ^ uncoded_block[1702];
  wire _24138 = _24137 ^ _8535;
  wire _24139 = _24136 ^ _24138;
  wire _24140 = _851 ^ _2443;
  wire _24141 = _15064 ^ _24140;
  wire _24142 = _24139 ^ _24141;
  wire _24143 = _24142 ^ uncoded_block[1722];
  wire _24144 = _24135 ^ _24143;
  wire _24145 = _24101 ^ _24144;
  wire _24146 = _23963 ^ _24145;
  wire _24147 = uncoded_block[4] ^ uncoded_block[7];
  wire _24148 = _21407 ^ _24147;
  wire _24149 = _24148 ^ _13535;
  wire _24150 = uncoded_block[25] ^ uncoded_block[29];
  wire _24151 = _24150 ^ _6095;
  wire _24152 = _4717 ^ _24151;
  wire _24153 = _24149 ^ _24152;
  wire _24154 = _21871 ^ _17065;
  wire _24155 = _3232 ^ _5435;
  wire _24156 = _24154 ^ _24155;
  wire _24157 = _23697 ^ _1705;
  wire _24158 = _4728 ^ _897;
  wire _24159 = _24157 ^ _24158;
  wire _24160 = _24156 ^ _24159;
  wire _24161 = _24153 ^ _24160;
  wire _24162 = _11363 ^ _10249;
  wire _24163 = _6757 ^ _4026;
  wire _24164 = _24162 ^ _24163;
  wire _24165 = _12443 ^ _4745;
  wire _24166 = _49 ^ _14595;
  wire _24167 = _24165 ^ _24166;
  wire _24168 = _24164 ^ _24167;
  wire _24169 = _6123 ^ _4034;
  wire _24170 = _24169 ^ _6770;
  wire _24171 = _12451 ^ _7386;
  wire _24172 = _6774 ^ _21898;
  wire _24173 = _24171 ^ _24172;
  wire _24174 = _24170 ^ _24173;
  wire _24175 = _24168 ^ _24174;
  wire _24176 = _24161 ^ _24175;
  wire _24177 = _926 ^ _7391;
  wire _24178 = uncoded_block[144] ^ uncoded_block[146];
  wire _24179 = _24178 ^ _14082;
  wire _24180 = _24177 ^ _24179;
  wire _24181 = _70 ^ _3271;
  wire _24182 = uncoded_block[157] ^ uncoded_block[160];
  wire _24183 = _24182 ^ _4053;
  wire _24184 = _24181 ^ _24183;
  wire _24185 = _24180 ^ _24184;
  wire _24186 = _5473 ^ _4057;
  wire _24187 = _4770 ^ _11935;
  wire _24188 = _24186 ^ _24187;
  wire _24189 = _2529 ^ _1763;
  wire _24190 = _5485 ^ _19546;
  wire _24191 = _24189 ^ _24190;
  wire _24192 = _24188 ^ _24191;
  wire _24193 = _24185 ^ _24192;
  wire _24194 = uncoded_block[214] ^ uncoded_block[219];
  wire _24195 = _956 ^ _24194;
  wire _24196 = _14102 ^ _24195;
  wire _24197 = _5492 ^ _17118;
  wire _24198 = _4081 ^ _967;
  wire _24199 = _24197 ^ _24198;
  wire _24200 = _24196 ^ _24199;
  wire _24201 = _21465 ^ _6180;
  wire _24202 = _22382 ^ _24201;
  wire _24203 = _14633 ^ _10298;
  wire _24204 = _24202 ^ _24203;
  wire _24205 = _24200 ^ _24204;
  wire _24206 = _24193 ^ _24205;
  wire _24207 = _24176 ^ _24206;
  wire _24208 = _6187 ^ _14122;
  wire _24209 = _130 ^ _1795;
  wire _24210 = _24208 ^ _24209;
  wire _24211 = _7445 ^ _11967;
  wire _24212 = uncoded_block[283] ^ uncoded_block[286];
  wire _24213 = _24212 ^ _2571;
  wire _24214 = _24211 ^ _24213;
  wire _24215 = _24210 ^ _24214;
  wire _24216 = uncoded_block[293] ^ uncoded_block[297];
  wire _24217 = _24216 ^ _15163;
  wire _24218 = _8056 ^ _3340;
  wire _24219 = _24217 ^ _24218;
  wire _24220 = uncoded_block[316] ^ uncoded_block[321];
  wire _24221 = _24220 ^ _11441;
  wire _24222 = _24221 ^ _7461;
  wire _24223 = _24219 ^ _24222;
  wire _24224 = _24215 ^ _24223;
  wire _24225 = _3352 ^ _8646;
  wire _24226 = uncoded_block[341] ^ uncoded_block[350];
  wire _24227 = _9242 ^ _24226;
  wire _24228 = _24225 ^ _24227;
  wire _24229 = uncoded_block[352] ^ uncoded_block[357];
  wire _24230 = _24229 ^ _6864;
  wire _24231 = _6866 ^ _168;
  wire _24232 = _24230 ^ _24231;
  wire _24233 = _24228 ^ _24232;
  wire _24234 = _1835 ^ _17658;
  wire _24235 = _6233 ^ _7476;
  wire _24236 = _24234 ^ _24235;
  wire _24237 = uncoded_block[390] ^ uncoded_block[394];
  wire _24238 = _17661 ^ _24237;
  wire _24239 = _24238 ^ _9808;
  wire _24240 = _24236 ^ _24239;
  wire _24241 = _24233 ^ _24240;
  wire _24242 = _24224 ^ _24241;
  wire _24243 = uncoded_block[409] ^ uncoded_block[411];
  wire _24244 = _184 ^ _24243;
  wire _24245 = uncoded_block[414] ^ uncoded_block[420];
  wire _24246 = _24245 ^ _194;
  wire _24247 = _24244 ^ _24246;
  wire _24248 = uncoded_block[424] ^ uncoded_block[427];
  wire _24249 = _24248 ^ _16184;
  wire _24250 = _13117 ^ _3405;
  wire _24251 = _24249 ^ _24250;
  wire _24252 = _24247 ^ _24251;
  wire _24253 = _21974 ^ _9275;
  wire _24254 = uncoded_block[447] ^ uncoded_block[450];
  wire _24255 = _24254 ^ _2645;
  wire _24256 = _24253 ^ _24255;
  wire _24257 = _6261 ^ _213;
  wire _24258 = _2653 ^ _1874;
  wire _24259 = _24257 ^ _24258;
  wire _24260 = _24256 ^ _24259;
  wire _24261 = _24252 ^ _24260;
  wire _24262 = _5592 ^ _2659;
  wire _24263 = _12024 ^ _24262;
  wire _24264 = _2660 ^ _3424;
  wire _24265 = _24264 ^ _13140;
  wire _24266 = _24263 ^ _24265;
  wire _24267 = _3434 ^ _6921;
  wire _24268 = _13674 ^ _9295;
  wire _24269 = _24267 ^ _24268;
  wire _24270 = uncoded_block[525] ^ uncoded_block[531];
  wire _24271 = _1108 ^ _24270;
  wire _24272 = _17206 ^ _24271;
  wire _24273 = _24269 ^ _24272;
  wire _24274 = _24266 ^ _24273;
  wire _24275 = _24261 ^ _24274;
  wire _24276 = _24242 ^ _24275;
  wire _24277 = _24207 ^ _24276;
  wire _24278 = _9309 ^ _1905;
  wire _24279 = uncoded_block[537] ^ uncoded_block[539];
  wire _24280 = _24279 ^ _1908;
  wire _24281 = _24278 ^ _24280;
  wire _24282 = uncoded_block[545] ^ uncoded_block[548];
  wire _24283 = _24282 ^ _8724;
  wire _24284 = uncoded_block[558] ^ uncoded_block[561];
  wire _24285 = _24284 ^ _3465;
  wire _24286 = _24283 ^ _24285;
  wire _24287 = _24281 ^ _24286;
  wire _24288 = _3467 ^ _1928;
  wire _24289 = uncoded_block[582] ^ uncoded_block[585];
  wire _24290 = _6947 ^ _24289;
  wire _24291 = _24288 ^ _24290;
  wire _24292 = _1141 ^ _6316;
  wire _24293 = _1939 ^ _12066;
  wire _24294 = _24292 ^ _24293;
  wire _24295 = _24291 ^ _24294;
  wire _24296 = _24287 ^ _24295;
  wire _24297 = _14218 ^ _12609;
  wire _24298 = _7559 ^ _24297;
  wire _24299 = uncoded_block[615] ^ uncoded_block[620];
  wire _24300 = _5652 ^ _24299;
  wire _24301 = _24300 ^ _13716;
  wire _24302 = _24298 ^ _24301;
  wire _24303 = _22950 ^ _5661;
  wire _24304 = _1161 ^ _2727;
  wire _24305 = _24303 ^ _24304;
  wire _24306 = _19181 ^ _2738;
  wire _24307 = _12626 ^ _24306;
  wire _24308 = _24305 ^ _24307;
  wire _24309 = _24302 ^ _24308;
  wire _24310 = _24296 ^ _24309;
  wire _24311 = _15273 ^ _17742;
  wire _24312 = _19185 ^ _8177;
  wire _24313 = _24311 ^ _24312;
  wire _24314 = uncoded_block[680] ^ uncoded_block[683];
  wire _24315 = _24314 ^ _1972;
  wire _24316 = _2751 ^ _326;
  wire _24317 = _24315 ^ _24316;
  wire _24318 = _24313 ^ _24317;
  wire _24319 = _11557 ^ _14250;
  wire _24320 = uncoded_block[705] ^ uncoded_block[709];
  wire _24321 = _24320 ^ _1192;
  wire _24322 = _24319 ^ _24321;
  wire _24323 = _10452 ^ _17762;
  wire _24324 = _9369 ^ _6374;
  wire _24325 = _24323 ^ _24324;
  wire _24326 = _24322 ^ _24325;
  wire _24327 = _24318 ^ _24326;
  wire _24328 = _7603 ^ _7005;
  wire _24329 = _11572 ^ _24328;
  wire _24330 = _4289 ^ _5699;
  wire _24331 = uncoded_block[750] ^ uncoded_block[754];
  wire _24332 = _24331 ^ _2778;
  wire _24333 = _24330 ^ _24332;
  wire _24334 = _24329 ^ _24333;
  wire _24335 = uncoded_block[760] ^ uncoded_block[769];
  wire _24336 = _4298 ^ _24335;
  wire _24337 = _6382 ^ _2792;
  wire _24338 = _24336 ^ _24337;
  wire _24339 = _7021 ^ _18277;
  wire _24340 = _24339 ^ _16284;
  wire _24341 = _24338 ^ _24340;
  wire _24342 = _24334 ^ _24341;
  wire _24343 = _24327 ^ _24342;
  wire _24344 = _24310 ^ _24343;
  wire _24345 = uncoded_block[800] ^ uncoded_block[804];
  wire _24346 = _383 ^ _24345;
  wire _24347 = _12127 ^ _10483;
  wire _24348 = _24346 ^ _24347;
  wire _24349 = _5046 ^ _2029;
  wire _24350 = uncoded_block[828] ^ uncoded_block[832];
  wire _24351 = _6399 ^ _24350;
  wire _24352 = _24349 ^ _24351;
  wire _24353 = _24348 ^ _24352;
  wire _24354 = _1250 ^ _5057;
  wire _24355 = _1256 ^ _2820;
  wire _24356 = _24354 ^ _24355;
  wire _24357 = uncoded_block[852] ^ uncoded_block[856];
  wire _24358 = _7643 ^ _24357;
  wire _24359 = _6410 ^ _5069;
  wire _24360 = _24358 ^ _24359;
  wire _24361 = _24356 ^ _24360;
  wire _24362 = _24353 ^ _24361;
  wire _24363 = uncoded_block[872] ^ uncoded_block[876];
  wire _24364 = _2828 ^ _24363;
  wire _24365 = _24364 ^ _16816;
  wire _24366 = _11056 ^ _11059;
  wire _24367 = uncoded_block[888] ^ uncoded_block[895];
  wire _24368 = _24367 ^ _1278;
  wire _24369 = _24366 ^ _24368;
  wire _24370 = _24365 ^ _24369;
  wire _24371 = _429 ^ _12159;
  wire _24372 = uncoded_block[907] ^ uncoded_block[911];
  wire _24373 = _24372 ^ _17818;
  wire _24374 = _24371 ^ _24373;
  wire _24375 = uncoded_block[916] ^ uncoded_block[920];
  wire _24376 = _24375 ^ _23471;
  wire _24377 = uncoded_block[926] ^ uncoded_block[929];
  wire _24378 = _24377 ^ _448;
  wire _24379 = _24376 ^ _24378;
  wire _24380 = _24374 ^ _24379;
  wire _24381 = _24370 ^ _24380;
  wire _24382 = _24362 ^ _24381;
  wire _24383 = uncoded_block[936] ^ uncoded_block[940];
  wire _24384 = _12717 ^ _24383;
  wire _24385 = _455 ^ _5777;
  wire _24386 = _24384 ^ _24385;
  wire _24387 = _4381 ^ _1307;
  wire _24388 = uncoded_block[963] ^ uncoded_block[967];
  wire _24389 = _10528 ^ _24388;
  wire _24390 = _24387 ^ _24389;
  wire _24391 = _24386 ^ _24390;
  wire _24392 = _13272 ^ _18329;
  wire _24393 = _13271 ^ _24392;
  wire _24394 = _12186 ^ _1318;
  wire _24395 = _24394 ^ _16340;
  wire _24396 = _24393 ^ _24395;
  wire _24397 = _24391 ^ _24396;
  wire _24398 = uncoded_block[997] ^ uncoded_block[1002];
  wire _24399 = _6453 ^ _24398;
  wire _24400 = uncoded_block[1004] ^ uncoded_block[1007];
  wire _24401 = _24400 ^ _5129;
  wire _24402 = _24399 ^ _24401;
  wire _24403 = _2891 ^ _2894;
  wire _24404 = _22589 ^ _24403;
  wire _24405 = _24402 ^ _24404;
  wire _24406 = _22593 ^ _4419;
  wire _24407 = _501 ^ _21218;
  wire _24408 = uncoded_block[1040] ^ uncoded_block[1042];
  wire _24409 = _24408 ^ _514;
  wire _24410 = _24407 ^ _24409;
  wire _24411 = _24406 ^ _24410;
  wire _24412 = _24405 ^ _24411;
  wire _24413 = _24397 ^ _24412;
  wire _24414 = _24382 ^ _24413;
  wire _24415 = _24344 ^ _24414;
  wire _24416 = _24277 ^ _24415;
  wire _24417 = uncoded_block[1049] ^ uncoded_block[1052];
  wire _24418 = _3681 ^ _24417;
  wire _24419 = _9465 ^ _11120;
  wire _24420 = _24418 ^ _24419;
  wire _24421 = _5153 ^ _9475;
  wire _24422 = _8893 ^ _6486;
  wire _24423 = _24421 ^ _24422;
  wire _24424 = _24420 ^ _24423;
  wire _24425 = _5834 ^ _1371;
  wire _24426 = _24425 ^ _1375;
  wire _24427 = _536 ^ _3698;
  wire _24428 = _11139 ^ _12224;
  wire _24429 = _24427 ^ _24428;
  wire _24430 = _24426 ^ _24429;
  wire _24431 = _24424 ^ _24430;
  wire _24432 = _8336 ^ _4451;
  wire _24433 = _23075 ^ _13322;
  wire _24434 = _24432 ^ _24433;
  wire _24435 = _5853 ^ _2944;
  wire _24436 = _24435 ^ _15895;
  wire _24437 = _24434 ^ _24436;
  wire _24438 = _1393 ^ _8345;
  wire _24439 = uncoded_block[1143] ^ uncoded_block[1146];
  wire _24440 = _24439 ^ _3725;
  wire _24441 = _24438 ^ _24440;
  wire _24442 = uncoded_block[1158] ^ uncoded_block[1162];
  wire _24443 = _577 ^ _24442;
  wire _24444 = _2964 ^ _17390;
  wire _24445 = _24443 ^ _24444;
  wire _24446 = _24441 ^ _24445;
  wire _24447 = _24437 ^ _24446;
  wire _24448 = _24431 ^ _24447;
  wire _24449 = _5870 ^ _1410;
  wire _24450 = _585 ^ _6519;
  wire _24451 = _24449 ^ _24450;
  wire _24452 = _2195 ^ _4486;
  wire _24453 = _2200 ^ _1420;
  wire _24454 = _24452 ^ _24453;
  wire _24455 = _24451 ^ _24454;
  wire _24456 = uncoded_block[1203] ^ uncoded_block[1207];
  wire _24457 = _17400 ^ _24456;
  wire _24458 = _6526 ^ _24457;
  wire _24459 = uncoded_block[1218] ^ uncoded_block[1222];
  wire _24460 = _3762 ^ _24459;
  wire _24461 = _5210 ^ _24460;
  wire _24462 = _24458 ^ _24461;
  wire _24463 = _24455 ^ _24462;
  wire _24464 = _8958 ^ _12819;
  wire _24465 = _18404 ^ _15927;
  wire _24466 = _24464 ^ _24465;
  wire _24467 = _4509 ^ _13365;
  wire _24468 = _2232 ^ _8388;
  wire _24469 = _24467 ^ _24468;
  wire _24470 = _24466 ^ _24469;
  wire _24471 = uncoded_block[1255] ^ uncoded_block[1258];
  wire _24472 = _24471 ^ _4514;
  wire _24473 = _5235 ^ _1458;
  wire _24474 = _24472 ^ _24473;
  wire _24475 = _11188 ^ _13374;
  wire _24476 = _24475 ^ _11748;
  wire _24477 = _24474 ^ _24476;
  wire _24478 = _24470 ^ _24477;
  wire _24479 = _24463 ^ _24478;
  wire _24480 = _24448 ^ _24479;
  wire _24481 = _12837 ^ _5243;
  wire _24482 = uncoded_block[1287] ^ uncoded_block[1288];
  wire _24483 = _24482 ^ _10646;
  wire _24484 = _24481 ^ _24483;
  wire _24485 = _2255 ^ _8991;
  wire _24486 = _21743 ^ _24485;
  wire _24487 = _24484 ^ _24486;
  wire _24488 = _8992 ^ _14430;
  wire _24489 = _14432 ^ _2262;
  wire _24490 = _24488 ^ _24489;
  wire _24491 = _9555 ^ _3814;
  wire _24492 = _8411 ^ _1489;
  wire _24493 = _24491 ^ _24492;
  wire _24494 = _24490 ^ _24493;
  wire _24495 = _24487 ^ _24494;
  wire _24496 = _13922 ^ _4551;
  wire _24497 = _2276 ^ _7815;
  wire _24498 = _24496 ^ _24497;
  wire _24499 = uncoded_block[1348] ^ uncoded_block[1351];
  wire _24500 = _3039 ^ _24499;
  wire _24501 = _3042 ^ _12857;
  wire _24502 = _24500 ^ _24501;
  wire _24503 = _24498 ^ _24502;
  wire _24504 = _16444 ^ _17945;
  wire _24505 = _16443 ^ _24504;
  wire _24506 = _12305 ^ _3055;
  wire _24507 = _24506 ^ _7220;
  wire _24508 = _24505 ^ _24507;
  wire _24509 = _24503 ^ _24508;
  wire _24510 = _24495 ^ _24509;
  wire _24511 = uncoded_block[1389] ^ uncoded_block[1391];
  wire _24512 = _24511 ^ _4569;
  wire _24513 = _24512 ^ _3067;
  wire _24514 = _9016 ^ _18452;
  wire _24515 = _8436 ^ _4580;
  wire _24516 = _24514 ^ _24515;
  wire _24517 = _24513 ^ _24516;
  wire _24518 = _20347 ^ _17960;
  wire _24519 = _3074 ^ _14977;
  wire _24520 = _24518 ^ _24519;
  wire _24521 = uncoded_block[1437] ^ uncoded_block[1439];
  wire _24522 = _24521 ^ _5304;
  wire _24523 = _716 ^ _6619;
  wire _24524 = _24522 ^ _24523;
  wire _24525 = _24520 ^ _24524;
  wire _24526 = _24517 ^ _24525;
  wire _24527 = _6620 ^ _3088;
  wire _24528 = uncoded_block[1463] ^ uncoded_block[1468];
  wire _24529 = _24528 ^ _18919;
  wire _24530 = _24527 ^ _24529;
  wire _24531 = uncoded_block[1474] ^ uncoded_block[1484];
  wire _24532 = _9608 ^ _24531;
  wire _24533 = _17980 ^ _1563;
  wire _24534 = _24532 ^ _24533;
  wire _24535 = _24530 ^ _24534;
  wire _24536 = _4610 ^ _12896;
  wire _24537 = _3890 ^ _7258;
  wire _24538 = _24536 ^ _24537;
  wire _24539 = uncoded_block[1507] ^ uncoded_block[1509];
  wire _24540 = _1572 ^ _24539;
  wire _24541 = _5334 ^ _3115;
  wire _24542 = _24540 ^ _24541;
  wire _24543 = _24538 ^ _24542;
  wire _24544 = _24535 ^ _24543;
  wire _24545 = _24526 ^ _24544;
  wire _24546 = _24510 ^ _24545;
  wire _24547 = _24480 ^ _24546;
  wire _24548 = _11267 ^ _3900;
  wire _24549 = uncoded_block[1532] ^ uncoded_block[1538];
  wire _24550 = _15007 ^ _24549;
  wire _24551 = _24548 ^ _24550;
  wire _24552 = _6651 ^ _1589;
  wire _24553 = _7274 ^ _6013;
  wire _24554 = _24552 ^ _24553;
  wire _24555 = _24551 ^ _24554;
  wire _24556 = _767 ^ _770;
  wire _24557 = uncoded_block[1558] ^ uncoded_block[1565];
  wire _24558 = _24557 ^ _1606;
  wire _24559 = _24556 ^ _24558;
  wire _24560 = _15026 ^ _4651;
  wire _24561 = _18952 ^ _16515;
  wire _24562 = _24560 ^ _24561;
  wire _24563 = _24559 ^ _24562;
  wire _24564 = _24555 ^ _24563;
  wire _24565 = uncoded_block[1593] ^ uncoded_block[1596];
  wire _24566 = _3146 ^ _24565;
  wire _24567 = _4659 ^ _6039;
  wire _24568 = _24566 ^ _24567;
  wire _24569 = _4660 ^ _4662;
  wire _24570 = _6042 ^ _16032;
  wire _24571 = _24569 ^ _24570;
  wire _24572 = _24568 ^ _24571;
  wire _24573 = _7912 ^ _6046;
  wire _24574 = _9656 ^ _7306;
  wire _24575 = _24573 ^ _24574;
  wire _24576 = uncoded_block[1639] ^ uncoded_block[1644];
  wire _24577 = _24576 ^ _6691;
  wire _24578 = uncoded_block[1650] ^ uncoded_block[1652];
  wire _24579 = uncoded_block[1653] ^ uncoded_block[1663];
  wire _24580 = _24578 ^ _24579;
  wire _24581 = _24577 ^ _24580;
  wire _24582 = _24575 ^ _24581;
  wire _24583 = _24572 ^ _24582;
  wire _24584 = _24564 ^ _24583;
  wire _24585 = _3179 ^ _4687;
  wire _24586 = uncoded_block[1669] ^ uncoded_block[1674];
  wire _24587 = _24586 ^ _12398;
  wire _24588 = _24585 ^ _24587;
  wire _24589 = _833 ^ _6061;
  wire _24590 = _24589 ^ _14544;
  wire _24591 = _24588 ^ _24590;
  wire _24592 = _1666 ^ _844;
  wire _24593 = _20436 ^ _16551;
  wire _24594 = _24592 ^ _24593;
  wire _24595 = _851 ^ _18531;
  wire _24596 = _24595 ^ uncoded_block[1721];
  wire _24597 = _24594 ^ _24596;
  wire _24598 = _24591 ^ _24597;
  wire _24599 = _24584 ^ _24598;
  wire _24600 = _24547 ^ _24599;
  wire _24601 = _24416 ^ _24600;
  wire _24602 = _0 ^ _21861;
  wire _24603 = _3995 ^ _3216;
  wire _24604 = _24602 ^ _24603;
  wire _24605 = _6087 ^ _10;
  wire _24606 = uncoded_block[25] ^ uncoded_block[31];
  wire _24607 = _24606 ^ _6095;
  wire _24608 = _24605 ^ _24607;
  wire _24609 = _24604 ^ _24608;
  wire _24610 = _8549 ^ _21871;
  wire _24611 = _7965 ^ _8554;
  wire _24612 = _24610 ^ _24611;
  wire _24613 = uncoded_block[51] ^ uncoded_block[58];
  wire _24614 = _9150 ^ _24613;
  wire _24615 = _10801 ^ _12435;
  wire _24616 = _24614 ^ _24615;
  wire _24617 = _24612 ^ _24616;
  wire _24618 = _24609 ^ _24617;
  wire _24619 = _5440 ^ _900;
  wire _24620 = _7979 ^ _6750;
  wire _24621 = _24619 ^ _24620;
  wire _24622 = _17077 ^ _14065;
  wire _24623 = _4739 ^ _4026;
  wire _24624 = _24622 ^ _24623;
  wire _24625 = _24621 ^ _24624;
  wire _24626 = _14069 ^ _17083;
  wire _24627 = _14595 ^ _2491;
  wire _24628 = uncoded_block[110] ^ uncoded_block[115];
  wire _24629 = _24628 ^ _54;
  wire _24630 = _24627 ^ _24629;
  wire _24631 = _24626 ^ _24630;
  wire _24632 = _24625 ^ _24631;
  wire _24633 = _24618 ^ _24632;
  wire _24634 = _2498 ^ _2502;
  wire _24635 = _4753 ^ _1735;
  wire _24636 = _24634 ^ _24635;
  wire _24637 = uncoded_block[134] ^ uncoded_block[141];
  wire _24638 = _24637 ^ _6138;
  wire _24639 = _17097 ^ _70;
  wire _24640 = _24638 ^ _24639;
  wire _24641 = _24636 ^ _24640;
  wire _24642 = uncoded_block[152] ^ uncoded_block[156];
  wire _24643 = _24642 ^ _4049;
  wire _24644 = _4053 ^ _81;
  wire _24645 = _24643 ^ _24644;
  wire _24646 = _13583 ^ _1759;
  wire _24647 = _3279 ^ _24646;
  wire _24648 = _24645 ^ _24647;
  wire _24649 = _24641 ^ _24648;
  wire _24650 = _945 ^ _19544;
  wire _24651 = _7411 ^ _15135;
  wire _24652 = _24650 ^ _24651;
  wire _24653 = _18586 ^ _10853;
  wire _24654 = _24652 ^ _24653;
  wire _24655 = uncoded_block[212] ^ uncoded_block[216];
  wire _24656 = _24655 ^ _2543;
  wire _24657 = uncoded_block[223] ^ uncoded_block[228];
  wire _24658 = _24657 ^ _2549;
  wire _24659 = _24656 ^ _24658;
  wire _24660 = uncoded_block[233] ^ uncoded_block[235];
  wire _24661 = _24660 ^ _970;
  wire _24662 = _2553 ^ _6180;
  wire _24663 = _24661 ^ _24662;
  wire _24664 = _24659 ^ _24663;
  wire _24665 = _24654 ^ _24664;
  wire _24666 = _24649 ^ _24665;
  wire _24667 = _24633 ^ _24666;
  wire _24668 = _11954 ^ _13053;
  wire _24669 = _20999 ^ _13055;
  wire _24670 = _24668 ^ _24669;
  wire _24671 = _7438 ^ _4096;
  wire _24672 = _3321 ^ _6833;
  wire _24673 = _24671 ^ _24672;
  wire _24674 = _24670 ^ _24673;
  wire _24675 = _10303 ^ _3325;
  wire _24676 = _24675 ^ _22396;
  wire _24677 = _4110 ^ _13071;
  wire _24678 = _4821 ^ _24677;
  wire _24679 = _24676 ^ _24678;
  wire _24680 = _24674 ^ _24679;
  wire _24681 = _12515 ^ _3338;
  wire _24682 = _3340 ^ _1814;
  wire _24683 = _24681 ^ _24682;
  wire _24684 = _1009 ^ _152;
  wire _24685 = uncoded_block[331] ^ uncoded_block[338];
  wire _24686 = _9235 ^ _24685;
  wire _24687 = _24684 ^ _24686;
  wire _24688 = _24683 ^ _24687;
  wire _24689 = _158 ^ _20547;
  wire _24690 = _5541 ^ _162;
  wire _24691 = _24689 ^ _24690;
  wire _24692 = _20554 ^ _6228;
  wire _24693 = _15183 ^ _13094;
  wire _24694 = _24692 ^ _24693;
  wire _24695 = _24691 ^ _24694;
  wire _24696 = _24688 ^ _24695;
  wire _24697 = _24680 ^ _24696;
  wire _24698 = _1036 ^ _13101;
  wire _24699 = _3380 ^ _10907;
  wire _24700 = _24698 ^ _24699;
  wire _24701 = uncoded_block[396] ^ uncoded_block[400];
  wire _24702 = _5554 ^ _24701;
  wire _24703 = uncoded_block[403] ^ uncoded_block[408];
  wire _24704 = _5559 ^ _24703;
  wire _24705 = _24702 ^ _24704;
  wire _24706 = _24700 ^ _24705;
  wire _24707 = uncoded_block[420] ^ uncoded_block[424];
  wire _24708 = _13112 ^ _24707;
  wire _24709 = _14683 ^ _24708;
  wire _24710 = _197 ^ _1857;
  wire _24711 = uncoded_block[438] ^ uncoded_block[442];
  wire _24712 = _10919 ^ _24711;
  wire _24713 = _24710 ^ _24712;
  wire _24714 = _24709 ^ _24713;
  wire _24715 = _24706 ^ _24714;
  wire _24716 = uncoded_block[444] ^ uncoded_block[448];
  wire _24717 = uncoded_block[449] ^ uncoded_block[452];
  wire _24718 = _24716 ^ _24717;
  wire _24719 = _5586 ^ _1874;
  wire _24720 = _24718 ^ _24719;
  wire _24721 = uncoded_block[472] ^ uncoded_block[475];
  wire _24722 = _6906 ^ _24721;
  wire _24723 = uncoded_block[476] ^ uncoded_block[479];
  wire _24724 = _24723 ^ _224;
  wire _24725 = _24722 ^ _24724;
  wire _24726 = _24720 ^ _24725;
  wire _24727 = uncoded_block[489] ^ uncoded_block[494];
  wire _24728 = _24727 ^ _5603;
  wire _24729 = _24728 ^ _18200;
  wire _24730 = _8705 ^ _19638;
  wire _24731 = _6923 ^ _24730;
  wire _24732 = _24729 ^ _24731;
  wire _24733 = _24726 ^ _24732;
  wire _24734 = _24715 ^ _24733;
  wire _24735 = _24697 ^ _24734;
  wire _24736 = _24667 ^ _24735;
  wire _24737 = _13684 ^ _20602;
  wire _24738 = _1109 ^ _24737;
  wire _24739 = _16215 ^ _7536;
  wire _24740 = _8132 ^ _1909;
  wire _24741 = _24739 ^ _24740;
  wire _24742 = _24738 ^ _24741;
  wire _24743 = _1915 ^ _23826;
  wire _24744 = _7543 ^ _24743;
  wire _24745 = uncoded_block[565] ^ uncoded_block[569];
  wire _24746 = _24745 ^ _262;
  wire _24747 = uncoded_block[576] ^ uncoded_block[581];
  wire _24748 = _24747 ^ _8733;
  wire _24749 = _24746 ^ _24748;
  wire _24750 = _24744 ^ _24749;
  wire _24751 = _24742 ^ _24750;
  wire _24752 = _20618 ^ _4953;
  wire _24753 = _2710 ^ _16233;
  wire _24754 = _24752 ^ _24753;
  wire _24755 = _17232 ^ _7564;
  wire _24756 = _13713 ^ _1946;
  wire _24757 = _24755 ^ _24756;
  wire _24758 = _24754 ^ _24757;
  wire _24759 = _12618 ^ _8159;
  wire _24760 = _12071 ^ _22950;
  wire _24761 = _24759 ^ _24760;
  wire _24762 = _17241 ^ _23848;
  wire _24763 = _24761 ^ _24762;
  wire _24764 = _24758 ^ _24763;
  wire _24765 = _24751 ^ _24764;
  wire _24766 = _14235 ^ _1961;
  wire _24767 = _3508 ^ _18705;
  wire _24768 = _24767 ^ _6345;
  wire _24769 = _24766 ^ _24768;
  wire _24770 = _1174 ^ _1177;
  wire _24771 = _19185 ^ _8761;
  wire _24772 = _24770 ^ _24771;
  wire _24773 = _3522 ^ _3526;
  wire _24774 = _15281 ^ _17753;
  wire _24775 = _24773 ^ _24774;
  wire _24776 = _24772 ^ _24775;
  wire _24777 = _24769 ^ _24776;
  wire _24778 = _8186 ^ _20143;
  wire _24779 = _14255 ^ _16761;
  wire _24780 = _24778 ^ _24779;
  wire _24781 = _3536 ^ _1983;
  wire _24782 = _24781 ^ _342;
  wire _24783 = _24780 ^ _24782;
  wire _24784 = _343 ^ _3544;
  wire _24785 = _14774 ^ _8200;
  wire _24786 = _24784 ^ _24785;
  wire _24787 = _7002 ^ _23425;
  wire _24788 = _20156 ^ _5012;
  wire _24789 = _24787 ^ _24788;
  wire _24790 = _24786 ^ _24789;
  wire _24791 = _24783 ^ _24790;
  wire _24792 = _24777 ^ _24791;
  wire _24793 = _24765 ^ _24792;
  wire _24794 = uncoded_block[747] ^ uncoded_block[752];
  wire _24795 = _24794 ^ _11012;
  wire _24796 = uncoded_block[760] ^ uncoded_block[764];
  wire _24797 = _359 ^ _24796;
  wire _24798 = _24795 ^ _24797;
  wire _24799 = uncoded_block[775] ^ uncoded_block[785];
  wire _24800 = _11018 ^ _24799;
  wire _24801 = _8215 ^ _374;
  wire _24802 = _24800 ^ _24801;
  wire _24803 = _24798 ^ _24802;
  wire _24804 = uncoded_block[795] ^ uncoded_block[800];
  wire _24805 = _24804 ^ _4317;
  wire _24806 = _24805 ^ _8227;
  wire _24807 = _392 ^ _10483;
  wire _24808 = uncoded_block[814] ^ uncoded_block[820];
  wire _24809 = _24808 ^ _21155;
  wire _24810 = _24807 ^ _24809;
  wire _24811 = _24806 ^ _24810;
  wire _24812 = _24803 ^ _24811;
  wire _24813 = _4328 ^ _12135;
  wire _24814 = _3590 ^ _16801;
  wire _24815 = _24813 ^ _24814;
  wire _24816 = _1254 ^ _5058;
  wire _24817 = _3597 ^ _5741;
  wire _24818 = _24816 ^ _24817;
  wire _24819 = _24815 ^ _24818;
  wire _24820 = _11048 ^ _5069;
  wire _24821 = _22540 ^ _6416;
  wire _24822 = _24820 ^ _24821;
  wire _24823 = _11620 ^ _16304;
  wire _24824 = _2838 ^ _4352;
  wire _24825 = _24823 ^ _24824;
  wire _24826 = _24822 ^ _24825;
  wire _24827 = _24819 ^ _24826;
  wire _24828 = _24812 ^ _24827;
  wire _24829 = _8248 ^ _4355;
  wire _24830 = _8250 ^ _5089;
  wire _24831 = _24829 ^ _24830;
  wire _24832 = uncoded_block[917] ^ uncoded_block[922];
  wire _24833 = _436 ^ _24832;
  wire _24834 = _19253 ^ _24833;
  wire _24835 = _24831 ^ _24834;
  wire _24836 = _2076 ^ _3637;
  wire _24837 = uncoded_block[934] ^ uncoded_block[938];
  wire _24838 = _24837 ^ _16832;
  wire _24839 = _24836 ^ _24838;
  wire _24840 = uncoded_block[946] ^ uncoded_block[949];
  wire _24841 = _2865 ^ _24840;
  wire _24842 = _7083 ^ _4385;
  wire _24843 = _24841 ^ _24842;
  wire _24844 = _24839 ^ _24843;
  wire _24845 = _24835 ^ _24844;
  wire _24846 = _1310 ^ _12180;
  wire _24847 = _11648 ^ _1314;
  wire _24848 = _24846 ^ _24847;
  wire _24849 = _2877 ^ _470;
  wire _24850 = _4391 ^ _2100;
  wire _24851 = _24849 ^ _24850;
  wire _24852 = _24848 ^ _24851;
  wire _24853 = uncoded_block[986] ^ uncoded_block[988];
  wire _24854 = _23038 ^ _24853;
  wire _24855 = uncoded_block[989] ^ uncoded_block[992];
  wire _24856 = _24855 ^ _479;
  wire _24857 = _24854 ^ _24856;
  wire _24858 = uncoded_block[1000] ^ uncoded_block[1003];
  wire _24859 = _480 ^ _24858;
  wire _24860 = _24400 ^ _13283;
  wire _24861 = _24859 ^ _24860;
  wire _24862 = _24857 ^ _24861;
  wire _24863 = _24852 ^ _24862;
  wire _24864 = _24845 ^ _24863;
  wire _24865 = _24828 ^ _24864;
  wire _24866 = _24793 ^ _24865;
  wire _24867 = _24736 ^ _24866;
  wire _24868 = _8296 ^ _9996;
  wire _24869 = _8871 ^ _8299;
  wire _24870 = _24868 ^ _24869;
  wire _24871 = _495 ^ _6472;
  wire _24872 = uncoded_block[1034] ^ uncoded_block[1041];
  wire _24873 = _24872 ^ _2130;
  wire _24874 = _24871 ^ _24873;
  wire _24875 = _24870 ^ _24874;
  wire _24876 = _1356 ^ _13295;
  wire _24877 = uncoded_block[1057] ^ uncoded_block[1063];
  wire _24878 = _24877 ^ _2921;
  wire _24879 = _24876 ^ _24878;
  wire _24880 = _3689 ^ _8892;
  wire _24881 = _8893 ^ _1370;
  wire _24882 = _24880 ^ _24881;
  wire _24883 = _24879 ^ _24882;
  wire _24884 = _24875 ^ _24883;
  wire _24885 = _13857 ^ _542;
  wire _24886 = _17866 ^ _24885;
  wire _24887 = _11139 ^ _3705;
  wire _24888 = _24887 ^ _3709;
  wire _24889 = _24886 ^ _24888;
  wire _24890 = _5175 ^ _3714;
  wire _24891 = _8918 ^ _24890;
  wire _24892 = _4455 ^ _5854;
  wire _24893 = _24892 ^ _10034;
  wire _24894 = _24891 ^ _24893;
  wire _24895 = _24889 ^ _24894;
  wire _24896 = _24884 ^ _24895;
  wire _24897 = _14380 ^ _5182;
  wire _24898 = _2179 ^ _3724;
  wire _24899 = _24897 ^ _24898;
  wire _24900 = _6505 ^ _4466;
  wire _24901 = _3727 ^ _11711;
  wire _24902 = _24900 ^ _24901;
  wire _24903 = _24899 ^ _24902;
  wire _24904 = _7749 ^ _4476;
  wire _24905 = _24904 ^ _8363;
  wire _24906 = _13339 ^ _10608;
  wire _24907 = _24906 ^ _11167;
  wire _24908 = _24905 ^ _24907;
  wire _24909 = _24903 ^ _24908;
  wire _24910 = uncoded_block[1193] ^ uncoded_block[1194];
  wire _24911 = _24910 ^ _22179;
  wire _24912 = _7160 ^ _12258;
  wire _24913 = _24911 ^ _24912;
  wire _24914 = _12813 ^ _605;
  wire _24915 = _24914 ^ _21267;
  wire _24916 = _24913 ^ _24915;
  wire _24917 = _1436 ^ _7169;
  wire _24918 = _24917 ^ _18856;
  wire _24919 = _23550 ^ _6543;
  wire _24920 = _8388 ^ _3001;
  wire _24921 = _24919 ^ _24920;
  wire _24922 = _24918 ^ _24921;
  wire _24923 = _24916 ^ _24922;
  wire _24924 = _24909 ^ _24923;
  wire _24925 = _24896 ^ _24924;
  wire _24926 = _7780 ^ _4514;
  wire _24927 = uncoded_block[1265] ^ uncoded_block[1268];
  wire _24928 = _24927 ^ _1459;
  wire _24929 = _24926 ^ _24928;
  wire _24930 = _628 ^ _9539;
  wire _24931 = _3794 ^ _12837;
  wire _24932 = _24930 ^ _24931;
  wire _24933 = _24929 ^ _24932;
  wire _24934 = _639 ^ _13380;
  wire _24935 = _1469 ^ _3015;
  wire _24936 = _24934 ^ _24935;
  wire _24937 = _4532 ^ _1472;
  wire _24938 = _6572 ^ _3808;
  wire _24939 = _24937 ^ _24938;
  wire _24940 = _24936 ^ _24939;
  wire _24941 = _24933 ^ _24940;
  wire _24942 = uncoded_block[1316] ^ uncoded_block[1320];
  wire _24943 = _14432 ^ _24942;
  wire _24944 = _3032 ^ _4545;
  wire _24945 = _24943 ^ _24944;
  wire _24946 = _1494 ^ _8413;
  wire _24947 = uncoded_block[1335] ^ uncoded_block[1343];
  wire _24948 = _24947 ^ _5268;
  wire _24949 = _24946 ^ _24948;
  wire _24950 = _24945 ^ _24949;
  wire _24951 = uncoded_block[1354] ^ uncoded_block[1360];
  wire _24952 = _670 ^ _24951;
  wire _24953 = _24952 ^ _6590;
  wire _24954 = uncoded_block[1371] ^ uncoded_block[1375];
  wire _24955 = _679 ^ _24954;
  wire _24956 = _3055 ^ _3058;
  wire _24957 = _24955 ^ _24956;
  wire _24958 = _24953 ^ _24957;
  wire _24959 = _24950 ^ _24958;
  wire _24960 = _24941 ^ _24959;
  wire _24961 = _7222 ^ _2293;
  wire _24962 = _3836 ^ _24961;
  wire _24963 = _13416 ^ _1517;
  wire _24964 = uncoded_block[1404] ^ uncoded_block[1408];
  wire _24965 = _24964 ^ _17461;
  wire _24966 = _24963 ^ _24965;
  wire _24967 = _24962 ^ _24966;
  wire _24968 = _13422 ^ _3072;
  wire _24969 = _3074 ^ _7844;
  wire _24970 = _24968 ^ _24969;
  wire _24971 = _8443 ^ _17470;
  wire _24972 = _4590 ^ _2321;
  wire _24973 = _24971 ^ _24972;
  wire _24974 = _24970 ^ _24973;
  wire _24975 = _24967 ^ _24974;
  wire _24976 = _10694 ^ _1544;
  wire _24977 = _24976 ^ _13438;
  wire _24978 = _3870 ^ _24070;
  wire _24979 = _3879 ^ _3097;
  wire _24980 = _24978 ^ _24979;
  wire _24981 = _24977 ^ _24980;
  wire _24982 = _3100 ^ _19887;
  wire _24983 = _740 ^ _17489;
  wire _24984 = _24982 ^ _24983;
  wire _24985 = _7864 ^ _18931;
  wire _24986 = _9053 ^ _6643;
  wire _24987 = _24985 ^ _24986;
  wire _24988 = _24984 ^ _24987;
  wire _24989 = _24981 ^ _24988;
  wire _24990 = _24975 ^ _24989;
  wire _24991 = _24960 ^ _24990;
  wire _24992 = _24925 ^ _24991;
  wire _24993 = _15004 ^ _7269;
  wire _24994 = uncoded_block[1531] ^ uncoded_block[1533];
  wire _24995 = _8473 ^ _24994;
  wire _24996 = _24993 ^ _24995;
  wire _24997 = _6648 ^ _2365;
  wire _24998 = _3129 ^ _7275;
  wire _24999 = _24997 ^ _24998;
  wire _25000 = _24996 ^ _24999;
  wire _25001 = uncoded_block[1552] ^ uncoded_block[1555];
  wire _25002 = _25001 ^ _24094;
  wire _25003 = uncoded_block[1561] ^ uncoded_block[1568];
  wire _25004 = uncoded_block[1572] ^ uncoded_block[1576];
  wire _25005 = _25003 ^ _25004;
  wire _25006 = _25002 ^ _25005;
  wire _25007 = _4651 ^ _2384;
  wire _25008 = uncoded_block[1585] ^ uncoded_block[1588];
  wire _25009 = _25008 ^ _789;
  wire _25010 = _25007 ^ _25009;
  wire _25011 = _25006 ^ _25010;
  wire _25012 = _25000 ^ _25011;
  wire _25013 = uncoded_block[1593] ^ uncoded_block[1600];
  wire _25014 = _25013 ^ _6039;
  wire _25015 = _5380 ^ _10181;
  wire _25016 = _25014 ^ _25015;
  wire _25017 = _18020 ^ _3160;
  wire _25018 = _22292 ^ _11307;
  wire _25019 = _25017 ^ _25018;
  wire _25020 = _25016 ^ _25019;
  wire _25021 = _7305 ^ _9659;
  wire _25022 = _25021 ^ _4672;
  wire _25023 = _5394 ^ _4677;
  wire _25024 = _4678 ^ _10760;
  wire _25025 = _25023 ^ _25024;
  wire _25026 = _25022 ^ _25025;
  wire _25027 = _25020 ^ _25026;
  wire _25028 = _25012 ^ _25027;
  wire _25029 = _4681 ^ _7318;
  wire _25030 = _8521 ^ _7323;
  wire _25031 = _9110 ^ _25030;
  wire _25032 = _25029 ^ _25031;
  wire _25033 = _12398 ^ _10766;
  wire _25034 = _4693 ^ _2429;
  wire _25035 = _25033 ^ _25034;
  wire _25036 = _6707 ^ _6710;
  wire _25037 = uncoded_block[1698] ^ uncoded_block[1700];
  wire _25038 = uncoded_block[1701] ^ uncoded_block[1706];
  wire _25039 = _25037 ^ _25038;
  wire _25040 = _25036 ^ _25039;
  wire _25041 = _25035 ^ _25040;
  wire _25042 = _25032 ^ _25041;
  wire _25043 = _3200 ^ uncoded_block[1719];
  wire _25044 = _3198 ^ _25043;
  wire _25045 = _25042 ^ _25044;
  wire _25046 = _25028 ^ _25045;
  wire _25047 = _24992 ^ _25046;
  wire _25048 = _24867 ^ _25047;
  wire _25049 = _0 ^ _6082;
  wire _25050 = _25049 ^ _10789;
  wire _25051 = _2458 ^ _3220;
  wire _25052 = _2456 ^ _25051;
  wire _25053 = _25050 ^ _25052;
  wire _25054 = uncoded_block[35] ^ uncoded_block[43];
  wire _25055 = _3224 ^ _25054;
  wire _25056 = _22795 ^ _886;
  wire _25057 = _25055 ^ _25056;
  wire _25058 = _2471 ^ _13553;
  wire _25059 = _16577 ^ _38;
  wire _25060 = _25058 ^ _25059;
  wire _25061 = _25057 ^ _25060;
  wire _25062 = _25053 ^ _25061;
  wire _25063 = _21881 ^ _18076;
  wire _25064 = _18077 ^ _15603;
  wire _25065 = _25063 ^ _25064;
  wire _25066 = _1718 ^ _47;
  wire _25067 = _910 ^ _17584;
  wire _25068 = _25066 ^ _25067;
  wire _25069 = _25065 ^ _25068;
  wire _25070 = uncoded_block[119] ^ uncoded_block[122];
  wire _25071 = _2495 ^ _25070;
  wire _25072 = _15104 ^ _25071;
  wire _25073 = uncoded_block[128] ^ uncoded_block[131];
  wire _25074 = _7386 ^ _25073;
  wire _25075 = uncoded_block[135] ^ uncoded_block[138];
  wire _25076 = _9177 ^ _25075;
  wire _25077 = _25074 ^ _25076;
  wire _25078 = _25072 ^ _25077;
  wire _25079 = _25069 ^ _25078;
  wire _25080 = _25062 ^ _25079;
  wire _25081 = _4043 ^ _1742;
  wire _25082 = uncoded_block[147] ^ uncoded_block[151];
  wire _25083 = _25082 ^ _71;
  wire _25084 = _25081 ^ _25083;
  wire _25085 = _2514 ^ _5472;
  wire _25086 = _1751 ^ _938;
  wire _25087 = _25085 ^ _25086;
  wire _25088 = _25084 ^ _25087;
  wire _25089 = _6149 ^ _85;
  wire _25090 = _25089 ^ _5480;
  wire _25091 = uncoded_block[185] ^ uncoded_block[192];
  wire _25092 = _25091 ^ _89;
  wire _25093 = _15135 ^ _6805;
  wire _25094 = _25092 ^ _25093;
  wire _25095 = _25090 ^ _25094;
  wire _25096 = _25088 ^ _25095;
  wire _25097 = _12479 ^ _956;
  wire _25098 = _959 ^ _4074;
  wire _25099 = _25097 ^ _25098;
  wire _25100 = _104 ^ _2545;
  wire _25101 = _109 ^ _6821;
  wire _25102 = _25100 ^ _25101;
  wire _25103 = _25099 ^ _25102;
  wire _25104 = uncoded_block[234] ^ uncoded_block[240];
  wire _25105 = _967 ^ _25104;
  wire _25106 = _6172 ^ _4799;
  wire _25107 = _25105 ^ _25106;
  wire _25108 = uncoded_block[261] ^ uncoded_block[263];
  wire _25109 = _3312 ^ _25108;
  wire _25110 = _17129 ^ _25109;
  wire _25111 = _25107 ^ _25110;
  wire _25112 = _25103 ^ _25111;
  wire _25113 = _25096 ^ _25112;
  wire _25114 = _25080 ^ _25113;
  wire _25115 = _4098 ^ _7440;
  wire _25116 = _3320 ^ _10300;
  wire _25117 = _25115 ^ _25116;
  wire _25118 = _8632 ^ _4819;
  wire _25119 = _13065 ^ _25118;
  wire _25120 = _25117 ^ _25119;
  wire _25121 = _10880 ^ _17144;
  wire _25122 = _4114 ^ _13619;
  wire _25123 = _25121 ^ _25122;
  wire _25124 = _3340 ^ _2580;
  wire _25125 = _11444 ^ _6853;
  wire _25126 = _25124 ^ _25125;
  wire _25127 = _25123 ^ _25126;
  wire _25128 = _25120 ^ _25127;
  wire _25129 = _4129 ^ _20547;
  wire _25130 = _17158 ^ _25129;
  wire _25131 = uncoded_block[356] ^ uncoded_block[363];
  wire _25132 = _19092 ^ _25131;
  wire _25133 = _17163 ^ _8076;
  wire _25134 = _25132 ^ _25133;
  wire _25135 = _25130 ^ _25134;
  wire _25136 = _13094 ^ _1036;
  wire _25137 = uncoded_block[378] ^ uncoded_block[382];
  wire _25138 = _25137 ^ _1039;
  wire _25139 = _25136 ^ _25138;
  wire _25140 = _2613 ^ _5554;
  wire _25141 = uncoded_block[398] ^ uncoded_block[403];
  wire _25142 = _8661 ^ _25141;
  wire _25143 = _25140 ^ _25142;
  wire _25144 = _25139 ^ _25143;
  wire _25145 = _25135 ^ _25144;
  wire _25146 = _25128 ^ _25145;
  wire _25147 = _6244 ^ _3391;
  wire _25148 = _8091 ^ _2630;
  wire _25149 = _25147 ^ _25148;
  wire _25150 = uncoded_block[415] ^ uncoded_block[420];
  wire _25151 = _25150 ^ _4874;
  wire _25152 = _25151 ^ _13116;
  wire _25153 = _25149 ^ _25152;
  wire _25154 = uncoded_block[434] ^ uncoded_block[439];
  wire _25155 = _25154 ^ _16190;
  wire _25156 = _10356 ^ _12562;
  wire _25157 = _25155 ^ _25156;
  wire _25158 = _17185 ^ _22907;
  wire _25159 = _25158 ^ _9284;
  wire _25160 = _25157 ^ _25159;
  wire _25161 = _25153 ^ _25160;
  wire _25162 = _1879 ^ _3421;
  wire _25163 = _25162 ^ _12570;
  wire _25164 = _4897 ^ _17198;
  wire _25165 = _25164 ^ _18661;
  wire _25166 = _25163 ^ _25165;
  wire _25167 = uncoded_block[504] ^ uncoded_block[507];
  wire _25168 = _6279 ^ _25167;
  wire _25169 = _6285 ^ _236;
  wire _25170 = _25168 ^ _25169;
  wire _25171 = uncoded_block[527] ^ uncoded_block[535];
  wire _25172 = _3445 ^ _25171;
  wire _25173 = uncoded_block[541] ^ uncoded_block[543];
  wire _25174 = _14197 ^ _25173;
  wire _25175 = _25172 ^ _25174;
  wire _25176 = _25170 ^ _25175;
  wire _25177 = _25166 ^ _25176;
  wire _25178 = _25161 ^ _25177;
  wire _25179 = _25146 ^ _25178;
  wire _25180 = _25114 ^ _25179;
  wire _25181 = _1117 ^ _1912;
  wire _25182 = uncoded_block[553] ^ uncoded_block[556];
  wire _25183 = _247 ^ _25182;
  wire _25184 = _25181 ^ _25183;
  wire _25185 = _1916 ^ _9319;
  wire _25186 = uncoded_block[570] ^ uncoded_block[572];
  wire _25187 = _20110 ^ _25186;
  wire _25188 = _25185 ^ _25187;
  wire _25189 = _25184 ^ _25188;
  wire _25190 = _3475 ^ _266;
  wire _25191 = _15748 ^ _25190;
  wire _25192 = _19656 ^ _6316;
  wire _25193 = _2706 ^ _4953;
  wire _25194 = _25192 ^ _25193;
  wire _25195 = _25191 ^ _25194;
  wire _25196 = _25189 ^ _25195;
  wire _25197 = _3487 ^ _8738;
  wire _25198 = _12609 ^ _16238;
  wire _25199 = _25197 ^ _25198;
  wire _25200 = _5658 ^ _22950;
  wire _25201 = _17237 ^ _25200;
  wire _25202 = _25199 ^ _25201;
  wire _25203 = _6331 ^ _1160;
  wire _25204 = _5665 ^ _6336;
  wire _25205 = _25203 ^ _25204;
  wire _25206 = uncoded_block[648] ^ uncoded_block[652];
  wire _25207 = _296 ^ _25206;
  wire _25208 = _19181 ^ _3508;
  wire _25209 = _25207 ^ _25208;
  wire _25210 = _25205 ^ _25209;
  wire _25211 = _25202 ^ _25210;
  wire _25212 = _25196 ^ _25211;
  wire _25213 = _3513 ^ _15273;
  wire _25214 = _10990 ^ _23410;
  wire _25215 = _25213 ^ _25214;
  wire _25216 = uncoded_block[680] ^ uncoded_block[691];
  wire _25217 = _25216 ^ _9895;
  wire _25218 = uncoded_block[701] ^ uncoded_block[705];
  wire _25219 = _19195 ^ _25218;
  wire _25220 = _25217 ^ _25219;
  wire _25221 = _25215 ^ _25220;
  wire _25222 = _8198 ^ _9905;
  wire _25223 = _23864 ^ _25222;
  wire _25224 = _3547 ^ _7005;
  wire _25225 = _1207 ^ _21136;
  wire _25226 = _25224 ^ _25225;
  wire _25227 = _25223 ^ _25226;
  wire _25228 = _25221 ^ _25227;
  wire _25229 = _5704 ^ _5016;
  wire _25230 = _4298 ^ _5019;
  wire _25231 = _25229 ^ _25230;
  wire _25232 = uncoded_block[765] ^ uncoded_block[770];
  wire _25233 = _1217 ^ _25232;
  wire _25234 = _12114 ^ _2014;
  wire _25235 = _25233 ^ _25234;
  wire _25236 = _25231 ^ _25235;
  wire _25237 = _2015 ^ _1224;
  wire _25238 = _1225 ^ _12676;
  wire _25239 = _25237 ^ _25238;
  wire _25240 = _5726 ^ _12127;
  wire _25241 = _2802 ^ _25240;
  wire _25242 = _25239 ^ _25241;
  wire _25243 = _25236 ^ _25242;
  wire _25244 = _25228 ^ _25243;
  wire _25245 = _25212 ^ _25244;
  wire _25246 = _5043 ^ _23000;
  wire _25247 = _23450 ^ _12135;
  wire _25248 = _7038 ^ _25247;
  wire _25249 = _25246 ^ _25248;
  wire _25250 = _5054 ^ _1254;
  wire _25251 = _4339 ^ _3599;
  wire _25252 = _25250 ^ _25251;
  wire _25253 = uncoded_block[860] ^ uncoded_block[867];
  wire _25254 = _20692 ^ _25253;
  wire _25255 = _5065 ^ _25254;
  wire _25256 = _25252 ^ _25255;
  wire _25257 = _25249 ^ _25256;
  wire _25258 = _4347 ^ _420;
  wire _25259 = _5079 ^ _8820;
  wire _25260 = _25258 ^ _25259;
  wire _25261 = _2058 ^ _7660;
  wire _25262 = uncoded_block[891] ^ uncoded_block[894];
  wire _25263 = _25262 ^ _3616;
  wire _25264 = _25261 ^ _25263;
  wire _25265 = _25260 ^ _25264;
  wire _25266 = _3617 ^ _1280;
  wire _25267 = _2070 ^ _5762;
  wire _25268 = _25266 ^ _25267;
  wire _25269 = _6434 ^ _2855;
  wire _25270 = _446 ^ _1296;
  wire _25271 = _25269 ^ _25270;
  wire _25272 = _25268 ^ _25271;
  wire _25273 = _25265 ^ _25272;
  wire _25274 = _25257 ^ _25273;
  wire _25275 = _2078 ^ _452;
  wire _25276 = _25275 ^ _6440;
  wire _25277 = _13266 ^ _9437;
  wire _25278 = _16834 ^ _25277;
  wire _25279 = _25276 ^ _25278;
  wire _25280 = _7680 ^ _4385;
  wire _25281 = _11646 ^ _11087;
  wire _25282 = _25280 ^ _25281;
  wire _25283 = uncoded_block[969] ^ uncoded_block[973];
  wire _25284 = _25283 ^ _470;
  wire _25285 = _25284 ^ _5791;
  wire _25286 = _25282 ^ _25285;
  wire _25287 = _25279 ^ _25286;
  wire _25288 = _5792 ^ _6451;
  wire _25289 = uncoded_block[991] ^ uncoded_block[994];
  wire _25290 = _23938 ^ _25289;
  wire _25291 = _25288 ^ _25290;
  wire _25292 = _13277 ^ _2107;
  wire _25293 = _25292 ^ _16850;
  wire _25294 = _25291 ^ _25293;
  wire _25295 = uncoded_block[1011] ^ uncoded_block[1013];
  wire _25296 = _25295 ^ _8871;
  wire _25297 = uncoded_block[1026] ^ uncoded_block[1031];
  wire _25298 = _5137 ^ _25297;
  wire _25299 = _25296 ^ _25298;
  wire _25300 = _9461 ^ _8306;
  wire _25301 = _8309 ^ _19295;
  wire _25302 = _25300 ^ _25301;
  wire _25303 = _25299 ^ _25302;
  wire _25304 = _25294 ^ _25303;
  wire _25305 = _25287 ^ _25304;
  wire _25306 = _25274 ^ _25305;
  wire _25307 = _25245 ^ _25306;
  wire _25308 = _25180 ^ _25307;
  wire _25309 = uncoded_block[1051] ^ uncoded_block[1057];
  wire _25310 = _25309 ^ _10566;
  wire _25311 = uncoded_block[1067] ^ uncoded_block[1072];
  wire _25312 = _14357 ^ _25311;
  wire _25313 = _25310 ^ _25312;
  wire _25314 = _529 ^ _2925;
  wire _25315 = _7724 ^ _8906;
  wire _25316 = _25314 ^ _25315;
  wire _25317 = _25313 ^ _25316;
  wire _25318 = uncoded_block[1097] ^ uncoded_block[1101];
  wire _25319 = _25318 ^ _11142;
  wire _25320 = _11138 ^ _25319;
  wire _25321 = uncoded_block[1104] ^ uncoded_block[1110];
  wire _25322 = _25321 ^ _4451;
  wire _25323 = uncoded_block[1113] ^ uncoded_block[1116];
  wire _25324 = _25323 ^ _8920;
  wire _25325 = _25322 ^ _25324;
  wire _25326 = _25320 ^ _25325;
  wire _25327 = _25317 ^ _25326;
  wire _25328 = _7736 ^ _2942;
  wire _25329 = _2944 ^ _15894;
  wire _25330 = _25328 ^ _25329;
  wire _25331 = _8343 ^ _1395;
  wire _25332 = uncoded_block[1142] ^ uncoded_block[1144];
  wire _25333 = _4462 ^ _25332;
  wire _25334 = _25331 ^ _25333;
  wire _25335 = _25330 ^ _25334;
  wire _25336 = _2180 ^ _8933;
  wire _25337 = _8937 ^ _578;
  wire _25338 = _25336 ^ _25337;
  wire _25339 = _8356 ^ _13335;
  wire _25340 = _4476 ^ _5870;
  wire _25341 = _25339 ^ _25340;
  wire _25342 = _25338 ^ _25341;
  wire _25343 = _25335 ^ _25342;
  wire _25344 = _25327 ^ _25343;
  wire _25345 = _1410 ^ _5195;
  wire _25346 = uncoded_block[1179] ^ uncoded_block[1183];
  wire _25347 = _25346 ^ _23996;
  wire _25348 = _25345 ^ _25347;
  wire _25349 = _2971 ^ _1420;
  wire _25350 = _6525 ^ _7758;
  wire _25351 = _25349 ^ _25350;
  wire _25352 = _25348 ^ _25351;
  wire _25353 = _2974 ^ _4491;
  wire _25354 = _25353 ^ _1429;
  wire _25355 = _2219 ^ _4499;
  wire _25356 = _4502 ^ _10061;
  wire _25357 = _25355 ^ _25356;
  wire _25358 = _25354 ^ _25357;
  wire _25359 = _25352 ^ _25358;
  wire _25360 = _1442 ^ _16915;
  wire _25361 = _14411 ^ _25360;
  wire _25362 = _10627 ^ _3777;
  wire _25363 = _8385 ^ _3780;
  wire _25364 = _25362 ^ _25363;
  wire _25365 = _25361 ^ _25364;
  wire _25366 = uncoded_block[1256] ^ uncoded_block[1261];
  wire _25367 = _25366 ^ _4516;
  wire _25368 = _2244 ^ _5905;
  wire _25369 = _25367 ^ _25368;
  wire _25370 = _1463 ^ _5908;
  wire _25371 = _25370 ^ _9542;
  wire _25372 = _25369 ^ _25371;
  wire _25373 = _25365 ^ _25372;
  wire _25374 = _25359 ^ _25373;
  wire _25375 = _25344 ^ _25374;
  wire _25376 = _6560 ^ _24482;
  wire _25377 = uncoded_block[1290] ^ uncoded_block[1293];
  wire _25378 = _25377 ^ _3801;
  wire _25379 = _25376 ^ _25378;
  wire _25380 = _645 ^ _6564;
  wire _25381 = _15462 ^ _3808;
  wire _25382 = _25380 ^ _25381;
  wire _25383 = _25379 ^ _25382;
  wire _25384 = _5919 ^ _23134;
  wire _25385 = _25384 ^ _24491;
  wire _25386 = _8411 ^ _8998;
  wire _25387 = _25386 ^ _9000;
  wire _25388 = _25385 ^ _25387;
  wire _25389 = _25383 ^ _25388;
  wire _25390 = _664 ^ _670;
  wire _25391 = _1499 ^ _25390;
  wire _25392 = _5272 ^ _6587;
  wire _25393 = uncoded_block[1361] ^ uncoded_block[1363];
  wire _25394 = _4559 ^ _25393;
  wire _25395 = _25392 ^ _25394;
  wire _25396 = _25391 ^ _25395;
  wire _25397 = _10665 ^ _14959;
  wire _25398 = _25397 ^ _20833;
  wire _25399 = uncoded_block[1384] ^ uncoded_block[1387];
  wire _25400 = _687 ^ _25399;
  wire _25401 = _12867 ^ _23157;
  wire _25402 = _25400 ^ _25401;
  wire _25403 = _25398 ^ _25402;
  wire _25404 = _25396 ^ _25403;
  wire _25405 = _25389 ^ _25404;
  wire _25406 = uncoded_block[1401] ^ uncoded_block[1406];
  wire _25407 = _1516 ^ _25406;
  wire _25408 = _9585 ^ _13947;
  wire _25409 = _25407 ^ _25408;
  wire _25410 = uncoded_block[1427] ^ uncoded_block[1435];
  wire _25411 = _4584 ^ _25410;
  wire _25412 = _15493 ^ _25411;
  wire _25413 = _25409 ^ _25412;
  wire _25414 = _1541 ^ _2322;
  wire _25415 = _21785 ^ _25414;
  wire _25416 = uncoded_block[1460] ^ uncoded_block[1465];
  wire _25417 = _3089 ^ _25416;
  wire _25418 = _721 ^ _25417;
  wire _25419 = _25415 ^ _25418;
  wire _25420 = _25413 ^ _25419;
  wire _25421 = _727 ^ _7247;
  wire _25422 = _25421 ^ _19413;
  wire _25423 = uncoded_block[1475] ^ uncoded_block[1478];
  wire _25424 = uncoded_block[1479] ^ uncoded_block[1487];
  wire _25425 = _25423 ^ _25424;
  wire _25426 = uncoded_block[1489] ^ uncoded_block[1491];
  wire _25427 = _25426 ^ _12896;
  wire _25428 = _25425 ^ _25427;
  wire _25429 = _25422 ^ _25428;
  wire _25430 = uncoded_block[1495] ^ uncoded_block[1499];
  wire _25431 = _25430 ^ _1571;
  wire _25432 = uncoded_block[1502] ^ uncoded_block[1506];
  wire _25433 = _25432 ^ _24539;
  wire _25434 = _25431 ^ _25433;
  wire _25435 = _7875 ^ _751;
  wire _25436 = _754 ^ _8473;
  wire _25437 = _25435 ^ _25436;
  wire _25438 = _25434 ^ _25437;
  wire _25439 = _25429 ^ _25438;
  wire _25440 = _25420 ^ _25439;
  wire _25441 = _25405 ^ _25440;
  wire _25442 = _25375 ^ _25441;
  wire _25443 = _6001 ^ _12914;
  wire _25444 = _6006 ^ _16010;
  wire _25445 = _25443 ^ _25444;
  wire _25446 = _4634 ^ _1596;
  wire _25447 = _2372 ^ _2376;
  wire _25448 = _25446 ^ _25447;
  wire _25449 = _25445 ^ _25448;
  wire _25450 = uncoded_block[1571] ^ uncoded_block[1574];
  wire _25451 = _11284 ^ _25450;
  wire _25452 = _25451 ^ _17510;
  wire _25453 = _1612 ^ _2386;
  wire _25454 = uncoded_block[1590] ^ uncoded_block[1593];
  wire _25455 = _14511 ^ _25454;
  wire _25456 = _25453 ^ _25455;
  wire _25457 = _25452 ^ _25456;
  wire _25458 = _25449 ^ _25457;
  wire _25459 = _13996 ^ _8500;
  wire _25460 = _12373 ^ _21831;
  wire _25461 = _25459 ^ _25460;
  wire _25462 = _16032 ^ _6046;
  wire _25463 = _18511 ^ _19929;
  wire _25464 = _25462 ^ _25463;
  wire _25465 = _25461 ^ _25464;
  wire _25466 = _7306 ^ _2407;
  wire _25467 = _2408 ^ _7312;
  wire _25468 = _25466 ^ _25467;
  wire _25469 = _3172 ^ _8515;
  wire _25470 = uncoded_block[1659] ^ uncoded_block[1664];
  wire _25471 = _3174 ^ _25470;
  wire _25472 = _25469 ^ _25471;
  wire _25473 = _25468 ^ _25472;
  wire _25474 = _25465 ^ _25473;
  wire _25475 = _25458 ^ _25474;
  wire _25476 = uncoded_block[1668] ^ uncoded_block[1671];
  wire _25477 = _7319 ^ _25476;
  wire _25478 = _6700 ^ _11319;
  wire _25479 = _25477 ^ _25478;
  wire _25480 = uncoded_block[1682] ^ uncoded_block[1686];
  wire _25481 = _7325 ^ _25480;
  wire _25482 = _25481 ^ _21391;
  wire _25483 = _25479 ^ _25482;
  wire _25484 = _6711 ^ _8535;
  wire _25485 = _22771 ^ _25484;
  wire _25486 = _848 ^ _851;
  wire _25487 = _22316 ^ _7944;
  wire _25488 = _25486 ^ _25487;
  wire _25489 = _25485 ^ _25488;
  wire _25490 = _25483 ^ _25489;
  wire _25491 = _25490 ^ _10217;
  wire _25492 = _25475 ^ _25491;
  wire _25493 = _25442 ^ _25492;
  wire _25494 = _25308 ^ _25493;
  wire _25495 = _0 ^ _6080;
  wire _25496 = _3993 ^ _9135;
  wire _25497 = _25495 ^ _25496;
  wire _25498 = uncoded_block[17] ^ uncoded_block[21];
  wire _25499 = _18541 ^ _25498;
  wire _25500 = _20453 ^ _2461;
  wire _25501 = _25499 ^ _25500;
  wire _25502 = _25497 ^ _25501;
  wire _25503 = _15080 ^ _15590;
  wire _25504 = _25503 ^ _5434;
  wire _25505 = _886 ^ _888;
  wire _25506 = _7364 ^ _13553;
  wire _25507 = _25505 ^ _25506;
  wire _25508 = _25504 ^ _25507;
  wire _25509 = _25502 ^ _25508;
  wire _25510 = _9705 ^ _11357;
  wire _25511 = _7976 ^ _12438;
  wire _25512 = _25510 ^ _25511;
  wire _25513 = _10246 ^ _17077;
  wire _25514 = _9713 ^ _12442;
  wire _25515 = _25513 ^ _25514;
  wire _25516 = _25512 ^ _25515;
  wire _25517 = uncoded_block[95] ^ uncoded_block[101];
  wire _25518 = _25517 ^ _3250;
  wire _25519 = _1722 ^ _19520;
  wire _25520 = _25518 ^ _25519;
  wire _25521 = uncoded_block[113] ^ uncoded_block[118];
  wire _25522 = _25521 ^ _2501;
  wire _25523 = _4753 ^ _3262;
  wire _25524 = _25522 ^ _25523;
  wire _25525 = _25520 ^ _25524;
  wire _25526 = _25516 ^ _25525;
  wire _25527 = _25509 ^ _25526;
  wire _25528 = _4754 ^ _3263;
  wire _25529 = _6136 ^ _24178;
  wire _25530 = _25528 ^ _25529;
  wire _25531 = _11383 ^ _20488;
  wire _25532 = _21906 ^ _4053;
  wire _25533 = _25531 ^ _25532;
  wire _25534 = _25530 ^ _25533;
  wire _25535 = _2516 ^ _7399;
  wire _25536 = _15123 ^ _1756;
  wire _25537 = _25535 ^ _25536;
  wire _25538 = _940 ^ _17106;
  wire _25539 = _7409 ^ _2531;
  wire _25540 = _25538 ^ _25539;
  wire _25541 = _25537 ^ _25540;
  wire _25542 = _25534 ^ _25541;
  wire _25543 = _10277 ^ _16116;
  wire _25544 = uncoded_block[199] ^ uncoded_block[206];
  wire _25545 = uncoded_block[207] ^ uncoded_block[215];
  wire _25546 = _25544 ^ _25545;
  wire _25547 = _25543 ^ _25546;
  wire _25548 = _17613 ^ _5497;
  wire _25549 = _2545 ^ _7422;
  wire _25550 = _25548 ^ _25549;
  wire _25551 = _25547 ^ _25550;
  wire _25552 = _20994 ^ _9756;
  wire _25553 = _10860 ^ _16626;
  wire _25554 = _25552 ^ _25553;
  wire _25555 = _4803 ^ _2559;
  wire _25556 = _119 ^ _20523;
  wire _25557 = _25555 ^ _25556;
  wire _25558 = _25554 ^ _25557;
  wire _25559 = _25551 ^ _25558;
  wire _25560 = _25542 ^ _25559;
  wire _25561 = _25527 ^ _25560;
  wire _25562 = _985 ^ _128;
  wire _25563 = _5512 ^ _4814;
  wire _25564 = _25562 ^ _25563;
  wire _25565 = _7448 ^ _16144;
  wire _25566 = _11425 ^ _25565;
  wire _25567 = _25564 ^ _25566;
  wire _25568 = _137 ^ _4824;
  wire _25569 = uncoded_block[306] ^ uncoded_block[311];
  wire _25570 = _1000 ^ _25569;
  wire _25571 = _25568 ^ _25570;
  wire _25572 = _16149 ^ _1008;
  wire _25573 = _13625 ^ _1014;
  wire _25574 = _25572 ^ _25573;
  wire _25575 = _25571 ^ _25574;
  wire _25576 = _25567 ^ _25575;
  wire _25577 = uncoded_block[331] ^ uncoded_block[334];
  wire _25578 = _2584 ^ _25577;
  wire _25579 = uncoded_block[335] ^ uncoded_block[345];
  wire _25580 = _25579 ^ _1023;
  wire _25581 = _25578 ^ _25580;
  wire _25582 = _1028 ^ _21497;
  wire _25583 = _5542 ^ _25582;
  wire _25584 = _25581 ^ _25583;
  wire _25585 = _6866 ^ _9250;
  wire _25586 = _25585 ^ _8656;
  wire _25587 = _10895 ^ _9798;
  wire _25588 = _25587 ^ _7477;
  wire _25589 = _25586 ^ _25588;
  wire _25590 = _25584 ^ _25589;
  wire _25591 = _25576 ^ _25590;
  wire _25592 = uncoded_block[383] ^ uncoded_block[389];
  wire _25593 = _25592 ^ _10908;
  wire _25594 = _25593 ^ _23782;
  wire _25595 = _2623 ^ _12545;
  wire _25596 = _25595 ^ _6886;
  wire _25597 = _25594 ^ _25596;
  wire _25598 = _6249 ^ _11477;
  wire _25599 = _1060 ^ _2637;
  wire _25600 = _25598 ^ _25599;
  wire _25601 = uncoded_block[437] ^ uncoded_block[440];
  wire _25602 = _25601 ^ _3408;
  wire _25603 = _9272 ^ _25602;
  wire _25604 = _25600 ^ _25603;
  wire _25605 = _25597 ^ _25604;
  wire _25606 = _1864 ^ _4176;
  wire _25607 = uncoded_block[450] ^ uncoded_block[454];
  wire _25608 = _25607 ^ _213;
  wire _25609 = _25606 ^ _25608;
  wire _25610 = _14697 ^ _21981;
  wire _25611 = _25609 ^ _25610;
  wire _25612 = _6266 ^ _21526;
  wire _25613 = _8110 ^ _8694;
  wire _25614 = _25612 ^ _25613;
  wire _25615 = _7516 ^ _225;
  wire _25616 = _1094 ^ _20592;
  wire _25617 = _25615 ^ _25616;
  wire _25618 = _25614 ^ _25617;
  wire _25619 = _25611 ^ _25618;
  wire _25620 = _25605 ^ _25619;
  wire _25621 = _25591 ^ _25620;
  wire _25622 = _25561 ^ _25621;
  wire _25623 = _6921 ^ _10375;
  wire _25624 = _7531 ^ _15220;
  wire _25625 = _25623 ^ _25624;
  wire _25626 = _4910 ^ _10947;
  wire _25627 = _6289 ^ _1114;
  wire _25628 = _25626 ^ _25627;
  wire _25629 = _25625 ^ _25628;
  wire _25630 = uncoded_block[546] ^ uncoded_block[552];
  wire _25631 = uncoded_block[554] ^ uncoded_block[557];
  wire _25632 = _25630 ^ _25631;
  wire _25633 = _8133 ^ _25632;
  wire _25634 = _23829 ^ _4224;
  wire _25635 = _8140 ^ _25634;
  wire _25636 = _25633 ^ _25635;
  wire _25637 = _25629 ^ _25636;
  wire _25638 = _12057 ^ _1138;
  wire _25639 = _25638 ^ _4231;
  wire _25640 = uncoded_block[596] ^ uncoded_block[599];
  wire _25641 = _25640 ^ _2707;
  wire _25642 = _10406 ^ _25641;
  wire _25643 = _25639 ^ _25642;
  wire _25644 = _2711 ^ _19165;
  wire _25645 = _7563 ^ _13713;
  wire _25646 = _4243 ^ _1946;
  wire _25647 = _25645 ^ _25646;
  wire _25648 = _25644 ^ _25647;
  wire _25649 = _25643 ^ _25648;
  wire _25650 = _25637 ^ _25649;
  wire _25651 = _10979 ^ _6966;
  wire _25652 = _8161 ^ _3501;
  wire _25653 = _25651 ^ _25652;
  wire _25654 = _11543 ^ _4255;
  wire _25655 = _6336 ^ _3505;
  wire _25656 = _25654 ^ _25655;
  wire _25657 = _25653 ^ _25656;
  wire _25658 = _8165 ^ _1960;
  wire _25659 = _19181 ^ _305;
  wire _25660 = _25658 ^ _25659;
  wire _25661 = _309 ^ _9886;
  wire _25662 = _16750 ^ _25661;
  wire _25663 = _25660 ^ _25662;
  wire _25664 = _25657 ^ _25663;
  wire _25665 = _19185 ^ _13731;
  wire _25666 = _25665 ^ _20647;
  wire _25667 = _2750 ^ _6358;
  wire _25668 = _3529 ^ _11562;
  wire _25669 = _25667 ^ _25668;
  wire _25670 = _25666 ^ _25669;
  wire _25671 = _6361 ^ _4996;
  wire _25672 = _2762 ^ _10452;
  wire _25673 = _25671 ^ _25672;
  wire _25674 = _17762 ^ _9369;
  wire _25675 = _5003 ^ _2768;
  wire _25676 = _25674 ^ _25675;
  wire _25677 = _25673 ^ _25676;
  wire _25678 = _25670 ^ _25677;
  wire _25679 = _25664 ^ _25678;
  wire _25680 = _25650 ^ _25679;
  wire _25681 = _7002 ^ _1995;
  wire _25682 = uncoded_block[741] ^ uncoded_block[752];
  wire _25683 = _7005 ^ _25682;
  wire _25684 = _25681 ^ _25683;
  wire _25685 = uncoded_block[754] ^ uncoded_block[758];
  wire _25686 = _25685 ^ _13761;
  wire _25687 = _10470 ^ _11019;
  wire _25688 = _25686 ^ _25687;
  wire _25689 = _25684 ^ _25688;
  wire _25690 = _15799 ^ _2014;
  wire _25691 = uncoded_block[781] ^ uncoded_block[783];
  wire _25692 = _13219 ^ _25691;
  wire _25693 = _25690 ^ _25692;
  wire _25694 = uncoded_block[784] ^ uncoded_block[787];
  wire _25695 = _25694 ^ _5033;
  wire _25696 = uncoded_block[791] ^ uncoded_block[796];
  wire _25697 = _25696 ^ _7628;
  wire _25698 = _25695 ^ _25697;
  wire _25699 = _25693 ^ _25698;
  wire _25700 = _25689 ^ _25699;
  wire _25701 = _3577 ^ _3581;
  wire _25702 = _5041 ^ _11596;
  wire _25703 = _25701 ^ _25702;
  wire _25704 = _5045 ^ _1241;
  wire _25705 = _25704 ^ _14292;
  wire _25706 = _25703 ^ _25705;
  wire _25707 = _7039 ^ _2033;
  wire _25708 = _16293 ^ _7043;
  wire _25709 = _25707 ^ _25708;
  wire _25710 = uncoded_block[841] ^ uncoded_block[846];
  wire _25711 = uncoded_block[849] ^ uncoded_block[851];
  wire _25712 = _25710 ^ _25711;
  wire _25713 = _2046 ^ _23010;
  wire _25714 = _25712 ^ _25713;
  wire _25715 = _25709 ^ _25714;
  wire _25716 = _25706 ^ _25715;
  wire _25717 = _25700 ^ _25716;
  wire _25718 = _17304 ^ _5072;
  wire _25719 = uncoded_block[875] ^ uncoded_block[877];
  wire _25720 = _9953 ^ _25719;
  wire _25721 = _25718 ^ _25720;
  wire _25722 = uncoded_block[878] ^ uncoded_block[886];
  wire _25723 = _25722 ^ _7660;
  wire _25724 = _4354 ^ _3614;
  wire _25725 = _25723 ^ _25724;
  wire _25726 = _25721 ^ _25725;
  wire _25727 = _5085 ^ _8826;
  wire _25728 = _2844 ^ _15345;
  wire _25729 = _25727 ^ _25728;
  wire _25730 = _2070 ^ _12708;
  wire _25731 = uncoded_block[913] ^ uncoded_block[915];
  wire _25732 = _25731 ^ _3631;
  wire _25733 = _25730 ^ _25732;
  wire _25734 = _25729 ^ _25733;
  wire _25735 = _25726 ^ _25734;
  wire _25736 = uncoded_block[933] ^ uncoded_block[937];
  wire _25737 = _4368 ^ _25736;
  wire _25738 = _8269 ^ _2086;
  wire _25739 = _25737 ^ _25738;
  wire _25740 = _5777 ^ _19748;
  wire _25741 = uncoded_block[959] ^ uncoded_block[964];
  wire _25742 = _2090 ^ _25741;
  wire _25743 = _25740 ^ _25742;
  wire _25744 = _25739 ^ _25743;
  wire _25745 = _7682 ^ _468;
  wire _25746 = _8286 ^ _8855;
  wire _25747 = _25745 ^ _25746;
  wire _25748 = _4401 ^ _8293;
  wire _25749 = _1319 ^ _25748;
  wire _25750 = _25747 ^ _25749;
  wire _25751 = _25744 ^ _25750;
  wire _25752 = _25735 ^ _25751;
  wire _25753 = _25717 ^ _25752;
  wire _25754 = _25680 ^ _25753;
  wire _25755 = _25622 ^ _25754;
  wire _25756 = _5798 ^ _7691;
  wire _25757 = _4404 ^ _484;
  wire _25758 = _25756 ^ _25757;
  wire _25759 = uncoded_block[1006] ^ uncoded_block[1011];
  wire _25760 = _25759 ^ _4412;
  wire _25761 = _8871 ^ _9998;
  wire _25762 = _25760 ^ _25761;
  wire _25763 = _25758 ^ _25762;
  wire _25764 = uncoded_block[1034] ^ uncoded_block[1038];
  wire _25765 = _25297 ^ _25764;
  wire _25766 = _6475 ^ _6478;
  wire _25767 = _25765 ^ _25766;
  wire _25768 = uncoded_block[1054] ^ uncoded_block[1058];
  wire _25769 = _2136 ^ _25768;
  wire _25770 = _25301 ^ _25769;
  wire _25771 = _25767 ^ _25770;
  wire _25772 = _25763 ^ _25771;
  wire _25773 = uncoded_block[1068] ^ uncoded_block[1070];
  wire _25774 = uncoded_block[1075] ^ uncoded_block[1079];
  wire _25775 = _25773 ^ _25774;
  wire _25776 = _6484 ^ _25775;
  wire _25777 = _12219 ^ _20753;
  wire _25778 = _25777 ^ _8907;
  wire _25779 = _25776 ^ _25778;
  wire _25780 = _537 ^ _5169;
  wire _25781 = _15405 ^ _8336;
  wire _25782 = _25780 ^ _25781;
  wire _25783 = _550 ^ _23075;
  wire _25784 = _13322 ^ _10587;
  wire _25785 = _25783 ^ _25784;
  wire _25786 = _25782 ^ _25785;
  wire _25787 = _25779 ^ _25786;
  wire _25788 = _25772 ^ _25787;
  wire _25789 = _558 ^ _9494;
  wire _25790 = uncoded_block[1139] ^ uncoded_block[1144];
  wire _25791 = _20266 ^ _25790;
  wire _25792 = _25789 ^ _25791;
  wire _25793 = uncoded_block[1154] ^ uncoded_block[1160];
  wire _25794 = _4468 ^ _25793;
  wire _25795 = _17385 ^ _25794;
  wire _25796 = _25792 ^ _25795;
  wire _25797 = _2958 ^ _21248;
  wire _25798 = _2967 ^ _5872;
  wire _25799 = _25797 ^ _25798;
  wire _25800 = _6519 ^ _2195;
  wire _25801 = _10053 ^ _1420;
  wire _25802 = _25800 ^ _25801;
  wire _25803 = _25799 ^ _25802;
  wire _25804 = _25796 ^ _25803;
  wire _25805 = uncoded_block[1194] ^ uncoded_block[1199];
  wire _25806 = _25805 ^ _6529;
  wire _25807 = _2216 ^ _4496;
  wire _25808 = _25806 ^ _25807;
  wire _25809 = _1432 ^ _3765;
  wire _25810 = _6532 ^ _8377;
  wire _25811 = _25809 ^ _25810;
  wire _25812 = _25808 ^ _25811;
  wire _25813 = _5221 ^ _6536;
  wire _25814 = _20295 ^ _25813;
  wire _25815 = _2995 ^ _6538;
  wire _25816 = uncoded_block[1250] ^ uncoded_block[1255];
  wire _25817 = _2232 ^ _25816;
  wire _25818 = _25815 ^ _25817;
  wire _25819 = _25814 ^ _25818;
  wire _25820 = _25812 ^ _25819;
  wire _25821 = _25804 ^ _25820;
  wire _25822 = _25788 ^ _25821;
  wire _25823 = _13369 ^ _627;
  wire _25824 = _7179 ^ _628;
  wire _25825 = _25823 ^ _25824;
  wire _25826 = uncoded_block[1273] ^ uncoded_block[1276];
  wire _25827 = _25826 ^ _5908;
  wire _25828 = _10077 ^ _639;
  wire _25829 = _25827 ^ _25828;
  wire _25830 = _25825 ^ _25829;
  wire _25831 = uncoded_block[1291] ^ uncoded_block[1299];
  wire _25832 = _25831 ^ _10650;
  wire _25833 = _648 ^ _3808;
  wire _25834 = _25832 ^ _25833;
  wire _25835 = _2261 ^ _18426;
  wire _25836 = _25835 ^ _24492;
  wire _25837 = _25834 ^ _25836;
  wire _25838 = _25830 ^ _25837;
  wire _25839 = _23139 ^ _4550;
  wire _25840 = _3034 ^ _13399;
  wire _25841 = _25839 ^ _25840;
  wire _25842 = _5266 ^ _24040;
  wire _25843 = _5938 ^ _5272;
  wire _25844 = _25842 ^ _25843;
  wire _25845 = _25841 ^ _25844;
  wire _25846 = _673 ^ _3045;
  wire _25847 = _7211 ^ _11226;
  wire _25848 = _25846 ^ _25847;
  wire _25849 = uncoded_block[1373] ^ uncoded_block[1376];
  wire _25850 = _25849 ^ _4564;
  wire _25851 = _10108 ^ _688;
  wire _25852 = _25850 ^ _25851;
  wire _25853 = _25848 ^ _25852;
  wire _25854 = _25845 ^ _25853;
  wire _25855 = _25838 ^ _25854;
  wire _25856 = uncoded_block[1396] ^ uncoded_block[1402];
  wire _25857 = _24511 ^ _25856;
  wire _25858 = _25857 ^ _3848;
  wire _25859 = _5963 ^ _16464;
  wire _25860 = _25858 ^ _25859;
  wire _25861 = _9588 ^ _2308;
  wire _25862 = _25861 ^ _5300;
  wire _25863 = _2313 ^ _14978;
  wire _25864 = _2319 ^ _9033;
  wire _25865 = _25863 ^ _25864;
  wire _25866 = _25862 ^ _25865;
  wire _25867 = _25860 ^ _25866;
  wire _25868 = _16970 ^ _6622;
  wire _25869 = _3088 ^ _8452;
  wire _25870 = _25868 ^ _25869;
  wire _25871 = uncoded_block[1467] ^ uncoded_block[1472];
  wire _25872 = _8455 ^ _25871;
  wire _25873 = _6627 ^ _1558;
  wire _25874 = _25872 ^ _25873;
  wire _25875 = _25870 ^ _25874;
  wire _25876 = _5989 ^ _13451;
  wire _25877 = uncoded_block[1493] ^ uncoded_block[1501];
  wire _25878 = _4610 ^ _25877;
  wire _25879 = _3894 ^ _750;
  wire _25880 = _25878 ^ _25879;
  wire _25881 = _25876 ^ _25880;
  wire _25882 = _25875 ^ _25881;
  wire _25883 = _25867 ^ _25882;
  wire _25884 = _25855 ^ _25883;
  wire _25885 = _25822 ^ _25884;
  wire _25886 = uncoded_block[1526] ^ uncoded_block[1535];
  wire _25887 = _16988 ^ _25886;
  wire _25888 = _7266 ^ _25887;
  wire _25889 = _3906 ^ _8478;
  wire _25890 = _6008 ^ _3912;
  wire _25891 = _25889 ^ _25890;
  wire _25892 = _25888 ^ _25891;
  wire _25893 = _8484 ^ _2372;
  wire _25894 = uncoded_block[1564] ^ uncoded_block[1568];
  wire _25895 = uncoded_block[1569] ^ uncoded_block[1570];
  wire _25896 = _25894 ^ _25895;
  wire _25897 = _25893 ^ _25896;
  wire _25898 = _25450 ^ _782;
  wire _25899 = _784 ^ _25008;
  wire _25900 = _25898 ^ _25899;
  wire _25901 = _25897 ^ _25900;
  wire _25902 = _25892 ^ _25901;
  wire _25903 = _16026 ^ _11847;
  wire _25904 = _25903 ^ _17017;
  wire _25905 = uncoded_block[1614] ^ uncoded_block[1618];
  wire _25906 = uncoded_block[1620] ^ uncoded_block[1624];
  wire _25907 = _25905 ^ _25906;
  wire _25908 = _1628 ^ _25907;
  wire _25909 = _25904 ^ _25908;
  wire _25910 = _1639 ^ _7914;
  wire _25911 = _12948 ^ _25910;
  wire _25912 = _2407 ^ _2412;
  wire _25913 = _12387 ^ _12389;
  wire _25914 = _25912 ^ _25913;
  wire _25915 = _25911 ^ _25914;
  wire _25916 = _25909 ^ _25915;
  wire _25917 = _25902 ^ _25916;
  wire _25918 = _12390 ^ _823;
  wire _25919 = _19939 ^ _3183;
  wire _25920 = _25918 ^ _25919;
  wire _25921 = _17538 ^ _4691;
  wire _25922 = _3965 ^ _13519;
  wire _25923 = _25921 ^ _25922;
  wire _25924 = _25920 ^ _25923;
  wire _25925 = uncoded_block[1699] ^ uncoded_block[1707];
  wire _25926 = _2430 ^ _25925;
  wire _25927 = _20433 ^ _25926;
  wire _25928 = uncoded_block[1714] ^ uncoded_block[1718];
  wire _25929 = _11879 ^ _25928;
  wire _25930 = _25929 ^ _861;
  wire _25931 = _25927 ^ _25930;
  wire _25932 = _25924 ^ _25931;
  wire _25933 = _25917 ^ _25932;
  wire _25934 = _25885 ^ _25933;
  wire _25935 = _25755 ^ _25934;
  wire _25936 = _0 ^ _14038;
  wire _25937 = uncoded_block[14] ^ uncoded_block[20];
  wire _25938 = _19001 ^ _25937;
  wire _25939 = _25936 ^ _25938;
  wire _25940 = _3219 ^ _4001;
  wire _25941 = uncoded_block[28] ^ uncoded_block[33];
  wire _25942 = _25941 ^ _16;
  wire _25943 = _25940 ^ _25942;
  wire _25944 = _25939 ^ _25943;
  wire _25945 = _11894 ^ _7965;
  wire _25946 = _3232 ^ _13547;
  wire _25947 = _25945 ^ _25946;
  wire _25948 = uncoded_block[53] ^ uncoded_block[59];
  wire _25949 = _25948 ^ _2472;
  wire _25950 = uncoded_block[67] ^ uncoded_block[69];
  wire _25951 = _2474 ^ _25950;
  wire _25952 = _25949 ^ _25951;
  wire _25953 = _25947 ^ _25952;
  wire _25954 = _25944 ^ _25953;
  wire _25955 = uncoded_block[79] ^ uncoded_block[81];
  wire _25956 = _19511 ^ _25955;
  wire _25957 = uncoded_block[86] ^ uncoded_block[89];
  wire _25958 = _9161 ^ _25957;
  wire _25959 = _25956 ^ _25958;
  wire _25960 = _4741 ^ _910;
  wire _25961 = _7986 ^ _911;
  wire _25962 = _25960 ^ _25961;
  wire _25963 = _25959 ^ _25962;
  wire _25964 = _19520 ^ _7990;
  wire _25965 = _2495 ^ _6128;
  wire _25966 = _25964 ^ _25965;
  wire _25967 = uncoded_block[120] ^ uncoded_block[124];
  wire _25968 = _25967 ^ _13017;
  wire _25969 = _4754 ^ _16599;
  wire _25970 = _25968 ^ _25969;
  wire _25971 = _25966 ^ _25970;
  wire _25972 = _25963 ^ _25971;
  wire _25973 = _25954 ^ _25972;
  wire _25974 = _6138 ^ _1742;
  wire _25975 = _25974 ^ _1746;
  wire _25976 = uncoded_block[157] ^ uncoded_block[166];
  wire _25977 = _20488 ^ _25976;
  wire _25978 = _1752 ^ _14614;
  wire _25979 = _25977 ^ _25978;
  wire _25980 = _25975 ^ _25979;
  wire _25981 = _11933 ^ _7408;
  wire _25982 = _25981 ^ _8013;
  wire _25983 = uncoded_block[199] ^ uncoded_block[202];
  wire _25984 = _6800 ^ _25983;
  wire _25985 = _1764 ^ _11405;
  wire _25986 = _25984 ^ _25985;
  wire _25987 = _25982 ^ _25986;
  wire _25988 = _25980 ^ _25987;
  wire _25989 = _98 ^ _1767;
  wire _25990 = uncoded_block[222] ^ uncoded_block[228];
  wire _25991 = _17613 ^ _25990;
  wire _25992 = _25989 ^ _25991;
  wire _25993 = uncoded_block[229] ^ uncoded_block[233];
  wire _25994 = _25993 ^ _10289;
  wire _25995 = _21465 ^ _8617;
  wire _25996 = _25994 ^ _25995;
  wire _25997 = _25992 ^ _25996;
  wire _25998 = _23746 ^ _119;
  wire _25999 = _17129 ^ _25998;
  wire _26000 = uncoded_block[264] ^ uncoded_block[267];
  wire _26001 = _6185 ^ _26000;
  wire _26002 = _14642 ^ _14124;
  wire _26003 = _26001 ^ _26002;
  wire _26004 = _25999 ^ _26003;
  wire _26005 = _25997 ^ _26004;
  wire _26006 = _25988 ^ _26005;
  wire _26007 = _25973 ^ _26006;
  wire _26008 = _20527 ^ _11424;
  wire _26009 = _1803 ^ _3327;
  wire _26010 = _26008 ^ _26009;
  wire _26011 = _9226 ^ _994;
  wire _26012 = uncoded_block[298] ^ uncoded_block[301];
  wire _26013 = _4820 ^ _26012;
  wire _26014 = _26011 ^ _26013;
  wire _26015 = _26010 ^ _26014;
  wire _26016 = uncoded_block[307] ^ uncoded_block[313];
  wire _26017 = _14652 ^ _26016;
  wire _26018 = _3340 ^ _11439;
  wire _26019 = _26017 ^ _26018;
  wire _26020 = _1008 ^ _15677;
  wire _26021 = uncoded_block[330] ^ uncoded_block[334];
  wire _26022 = _21947 ^ _26021;
  wire _26023 = _26020 ^ _26022;
  wire _26024 = _26019 ^ _26023;
  wire _26025 = _26015 ^ _26024;
  wire _26026 = uncoded_block[338] ^ uncoded_block[341];
  wire _26027 = _2592 ^ _26026;
  wire _26028 = _6859 ^ _1023;
  wire _26029 = _26027 ^ _26028;
  wire _26030 = _24690 ^ _2603;
  wire _26031 = _26029 ^ _26030;
  wire _26032 = uncoded_block[363] ^ uncoded_block[366];
  wire _26033 = _2606 ^ _26032;
  wire _26034 = _1835 ^ _1838;
  wire _26035 = _26033 ^ _26034;
  wire _26036 = _4853 ^ _4143;
  wire _26037 = _26036 ^ _10337;
  wire _26038 = _26035 ^ _26037;
  wire _26039 = _26031 ^ _26038;
  wire _26040 = _26025 ^ _26039;
  wire _26041 = _6239 ^ _3383;
  wire _26042 = uncoded_block[396] ^ uncoded_block[398];
  wire _26043 = _1847 ^ _26042;
  wire _26044 = _26041 ^ _26043;
  wire _26045 = uncoded_block[407] ^ uncoded_block[410];
  wire _26046 = _26045 ^ _9266;
  wire _26047 = _6885 ^ _26046;
  wire _26048 = _26044 ^ _26047;
  wire _26049 = _5565 ^ _6249;
  wire _26050 = _26049 ^ _4165;
  wire _26051 = _2633 ^ _6894;
  wire _26052 = _6254 ^ _201;
  wire _26053 = _26051 ^ _26052;
  wire _26054 = _26050 ^ _26053;
  wire _26055 = _26048 ^ _26054;
  wire _26056 = _12559 ^ _10356;
  wire _26057 = _8677 ^ _26056;
  wire _26058 = _4177 ^ _1075;
  wire _26059 = _1076 ^ _8681;
  wire _26060 = _26058 ^ _26059;
  wire _26061 = _26057 ^ _26060;
  wire _26062 = _4181 ^ _1874;
  wire _26063 = _12023 ^ _1879;
  wire _26064 = _26062 ^ _26063;
  wire _26065 = _11494 ^ _1085;
  wire _26066 = uncoded_block[481] ^ uncoded_block[489];
  wire _26067 = _26066 ^ _10937;
  wire _26068 = _26065 ^ _26067;
  wire _26069 = _26064 ^ _26068;
  wire _26070 = _26061 ^ _26069;
  wire _26071 = _26055 ^ _26070;
  wire _26072 = _26040 ^ _26071;
  wire _26073 = _26007 ^ _26072;
  wire _26074 = _6279 ^ _1887;
  wire _26075 = _13140 ^ _26074;
  wire _26076 = _7529 ^ _4908;
  wire _26077 = _3439 ^ _1107;
  wire _26078 = _26076 ^ _26077;
  wire _26079 = _26075 ^ _26078;
  wire _26080 = uncoded_block[522] ^ uncoded_block[526];
  wire _26081 = uncoded_block[527] ^ uncoded_block[534];
  wire _26082 = _26080 ^ _26081;
  wire _26083 = _14719 ^ _14198;
  wire _26084 = _26082 ^ _26083;
  wire _26085 = _5628 ^ _8720;
  wire _26086 = _8721 ^ _1123;
  wire _26087 = _26085 ^ _26086;
  wire _26088 = _26084 ^ _26087;
  wire _26089 = _26079 ^ _26088;
  wire _26090 = uncoded_block[558] ^ uncoded_block[563];
  wire _26091 = _26090 ^ _1126;
  wire _26092 = _3468 ^ _17221;
  wire _26093 = _26091 ^ _26092;
  wire _26094 = uncoded_block[573] ^ uncoded_block[579];
  wire _26095 = _26094 ^ _6947;
  wire _26096 = uncoded_block[586] ^ uncoded_block[589];
  wire _26097 = _2696 ^ _26096;
  wire _26098 = _26095 ^ _26097;
  wire _26099 = _26093 ^ _26098;
  wire _26100 = _2700 ^ _15247;
  wire _26101 = _26100 ^ _25193;
  wire _26102 = _15757 ^ _12609;
  wire _26103 = _26102 ^ _17726;
  wire _26104 = _26101 ^ _26103;
  wire _26105 = _26099 ^ _26104;
  wire _26106 = _26089 ^ _26105;
  wire _26107 = _20125 ^ _14224;
  wire _26108 = uncoded_block[631] ^ uncoded_block[635];
  wire _26109 = _5658 ^ _26108;
  wire _26110 = _26107 ^ _26109;
  wire _26111 = _4249 ^ _22479;
  wire _26112 = uncoded_block[646] ^ uncoded_block[649];
  wire _26113 = _4972 ^ _26112;
  wire _26114 = _26111 ^ _26113;
  wire _26115 = _26110 ^ _26114;
  wire _26116 = _303 ^ _23852;
  wire _26117 = uncoded_block[664] ^ uncoded_block[669];
  wire _26118 = _12630 ^ _26117;
  wire _26119 = _26118 ^ _10435;
  wire _26120 = _26116 ^ _26119;
  wire _26121 = _26115 ^ _26120;
  wire _26122 = _3521 ^ _5678;
  wire _26123 = _26122 ^ _22491;
  wire _26124 = _4987 ^ _19195;
  wire _26125 = _11562 ^ _6361;
  wire _26126 = _26124 ^ _26125;
  wire _26127 = _26123 ^ _26126;
  wire _26128 = _3533 ^ _8190;
  wire _26129 = _26128 ^ _20656;
  wire _26130 = _4999 ^ _5690;
  wire _26131 = _9904 ^ _4286;
  wire _26132 = _26130 ^ _26131;
  wire _26133 = _26129 ^ _26132;
  wire _26134 = _26127 ^ _26133;
  wire _26135 = _26121 ^ _26134;
  wire _26136 = _26106 ^ _26135;
  wire _26137 = uncoded_block[731] ^ uncoded_block[739];
  wire _26138 = _26137 ^ _1207;
  wire _26139 = _26138 ^ _22506;
  wire _26140 = _2002 ^ _8779;
  wire _26141 = _3559 ^ _13761;
  wire _26142 = _26140 ^ _26141;
  wire _26143 = _26139 ^ _26142;
  wire _26144 = uncoded_block[764] ^ uncoded_block[772];
  wire _26145 = _26144 ^ _2012;
  wire _26146 = _14278 ^ _13219;
  wire _26147 = _26145 ^ _26146;
  wire _26148 = _18277 ^ _1224;
  wire _26149 = _4311 ^ _4314;
  wire _26150 = _26148 ^ _26149;
  wire _26151 = _26147 ^ _26150;
  wire _26152 = _26143 ^ _26151;
  wire _26153 = _1233 ^ _383;
  wire _26154 = _12126 ^ _3581;
  wire _26155 = _26153 ^ _26154;
  wire _26156 = _11596 ^ _9397;
  wire _26157 = _1242 ^ _23450;
  wire _26158 = _26156 ^ _26157;
  wire _26159 = _26155 ^ _26158;
  wire _26160 = uncoded_block[830] ^ uncoded_block[836];
  wire _26161 = _26160 ^ _14809;
  wire _26162 = _7640 ^ _1257;
  wire _26163 = _26161 ^ _26162;
  wire _26164 = uncoded_block[850] ^ uncoded_block[853];
  wire _26165 = _26164 ^ _15330;
  wire _26166 = _6410 ^ _413;
  wire _26167 = _26165 ^ _26166;
  wire _26168 = _26163 ^ _26167;
  wire _26169 = _26159 ^ _26168;
  wire _26170 = _26152 ^ _26169;
  wire _26171 = uncoded_block[864] ^ uncoded_block[868];
  wire _26172 = _26171 ^ _6415;
  wire _26173 = _13791 ^ _12151;
  wire _26174 = _26172 ^ _26173;
  wire _26175 = _20696 ^ _8820;
  wire _26176 = _13797 ^ _11060;
  wire _26177 = _26175 ^ _26176;
  wire _26178 = _26174 ^ _26177;
  wire _26179 = _4355 ^ _8826;
  wire _26180 = _429 ^ _2065;
  wire _26181 = _26179 ^ _26180;
  wire _26182 = _431 ^ _19252;
  wire _26183 = uncoded_block[921] ^ uncoded_block[927];
  wire _26184 = _21182 ^ _26183;
  wire _26185 = _26182 ^ _26184;
  wire _26186 = _26181 ^ _26185;
  wire _26187 = _26178 ^ _26186;
  wire _26188 = _448 ^ _5101;
  wire _26189 = uncoded_block[938] ^ uncoded_block[945];
  wire _26190 = _26189 ^ _5777;
  wire _26191 = _26188 ^ _26190;
  wire _26192 = _8274 ^ _9437;
  wire _26193 = uncoded_block[962] ^ uncoded_block[967];
  wire _26194 = _4385 ^ _26193;
  wire _26195 = _26192 ^ _26194;
  wire _26196 = _26191 ^ _26195;
  wire _26197 = uncoded_block[968] ^ uncoded_block[972];
  wire _26198 = _26197 ^ _470;
  wire _26199 = _26198 ^ _10535;
  wire _26200 = _13822 ^ _8856;
  wire _26201 = _26200 ^ _24856;
  wire _26202 = _26199 ^ _26201;
  wire _26203 = _26196 ^ _26202;
  wire _26204 = _26187 ^ _26203;
  wire _26205 = _26170 ^ _26204;
  wire _26206 = _26136 ^ _26205;
  wire _26207 = _26073 ^ _26206;
  wire _26208 = uncoded_block[998] ^ uncoded_block[1005];
  wire _26209 = _13277 ^ _26208;
  wire _26210 = _26209 ^ _7099;
  wire _26211 = _5131 ^ _5134;
  wire _26212 = _8872 ^ _3675;
  wire _26213 = _26211 ^ _26212;
  wire _26214 = _26210 ^ _26213;
  wire _26215 = _22595 ^ _512;
  wire _26216 = _514 ^ _23964;
  wire _26217 = _26215 ^ _26216;
  wire _26218 = _15871 ^ _519;
  wire _26219 = _26218 ^ _1365;
  wire _26220 = _26217 ^ _26219;
  wire _26221 = _26214 ^ _26220;
  wire _26222 = _8889 ^ _8892;
  wire _26223 = _2924 ^ _8895;
  wire _26224 = _26222 ^ _26223;
  wire _26225 = uncoded_block[1083] ^ uncoded_block[1089];
  wire _26226 = _26225 ^ _10026;
  wire _26227 = uncoded_block[1101] ^ uncoded_block[1105];
  wire _26228 = _5846 ^ _26227;
  wire _26229 = _26226 ^ _26228;
  wire _26230 = _26224 ^ _26229;
  wire _26231 = _549 ^ _13319;
  wire _26232 = _5175 ^ _8343;
  wire _26233 = _26231 ^ _26232;
  wire _26234 = _561 ^ _6501;
  wire _26235 = _10593 ^ _567;
  wire _26236 = _26234 ^ _26235;
  wire _26237 = _26233 ^ _26236;
  wire _26238 = _26230 ^ _26237;
  wire _26239 = _26221 ^ _26238;
  wire _26240 = uncoded_block[1150] ^ uncoded_block[1154];
  wire _26241 = _568 ^ _26240;
  wire _26242 = _9500 ^ _24442;
  wire _26243 = _26241 ^ _26242;
  wire _26244 = uncoded_block[1163] ^ uncoded_block[1166];
  wire _26245 = _26244 ^ _4476;
  wire _26246 = _26245 ^ _24449;
  wire _26247 = _26243 ^ _26246;
  wire _26248 = _5872 ^ _3742;
  wire _26249 = _26248 ^ _4487;
  wire _26250 = uncoded_block[1192] ^ uncoded_block[1197];
  wire _26251 = _2971 ^ _26250;
  wire _26252 = _26251 ^ _24457;
  wire _26253 = _26249 ^ _26252;
  wire _26254 = _26247 ^ _26253;
  wire _26255 = _23544 ^ _18395;
  wire _26256 = uncoded_block[1224] ^ uncoded_block[1228];
  wire _26257 = _4498 ^ _26256;
  wire _26258 = _26255 ^ _26257;
  wire _26259 = _2995 ^ _2997;
  wire _26260 = _21729 ^ _26259;
  wire _26261 = _26258 ^ _26260;
  wire _26262 = _2998 ^ _2235;
  wire _26263 = _7780 ^ _8970;
  wire _26264 = _26262 ^ _26263;
  wire _26265 = _628 ^ _2247;
  wire _26266 = _13371 ^ _26265;
  wire _26267 = _26264 ^ _26266;
  wire _26268 = _26261 ^ _26267;
  wire _26269 = _26254 ^ _26268;
  wire _26270 = _26239 ^ _26269;
  wire _26271 = uncoded_block[1282] ^ uncoded_block[1287];
  wire _26272 = _631 ^ _26271;
  wire _26273 = _26272 ^ _16927;
  wire _26274 = uncoded_block[1294] ^ uncoded_block[1298];
  wire _26275 = _26274 ^ _16424;
  wire _26276 = uncoded_block[1308] ^ uncoded_block[1312];
  wire _26277 = _26276 ^ _21748;
  wire _26278 = _26275 ^ _26277;
  wire _26279 = _26273 ^ _26278;
  wire _26280 = _7805 ^ _3814;
  wire _26281 = _26280 ^ _3033;
  wire _26282 = _4553 ^ _5937;
  wire _26283 = _662 ^ _26282;
  wire _26284 = _26281 ^ _26283;
  wire _26285 = _26279 ^ _26284;
  wire _26286 = _14447 ^ _7211;
  wire _26287 = _24501 ^ _26286;
  wire _26288 = _684 ^ _2289;
  wire _26289 = _5284 ^ _3059;
  wire _26290 = _26288 ^ _26289;
  wire _26291 = _26287 ^ _26290;
  wire _26292 = _25399 ^ _1513;
  wire _26293 = _26292 ^ _12873;
  wire _26294 = _6600 ^ _1519;
  wire _26295 = _16954 ^ _8436;
  wire _26296 = _26294 ^ _26295;
  wire _26297 = _26293 ^ _26296;
  wire _26298 = _26291 ^ _26297;
  wire _26299 = _26285 ^ _26298;
  wire _26300 = _4580 ^ _20347;
  wire _26301 = uncoded_block[1417] ^ uncoded_block[1421];
  wire _26302 = _8438 ^ _26301;
  wire _26303 = _26300 ^ _26302;
  wire _26304 = _9588 ^ _17963;
  wire _26305 = _5968 ^ _16962;
  wire _26306 = _26304 ^ _26305;
  wire _26307 = _26303 ^ _26306;
  wire _26308 = _15982 ^ _5970;
  wire _26309 = uncoded_block[1448] ^ uncoded_block[1450];
  wire _26310 = _26309 ^ _11247;
  wire _26311 = _26308 ^ _26310;
  wire _26312 = _723 ^ _8452;
  wire _26313 = _10699 ^ _1551;
  wire _26314 = _26312 ^ _26313;
  wire _26315 = _26311 ^ _26314;
  wire _26316 = _26307 ^ _26315;
  wire _26317 = _1556 ^ _7251;
  wire _26318 = _26317 ^ _24536;
  wire _26319 = _26318 ^ _7261;
  wire _26320 = _24539 ^ _7875;
  wire _26321 = uncoded_block[1513] ^ uncoded_block[1518];
  wire _26322 = _26321 ^ _22723;
  wire _26323 = _26320 ^ _26322;
  wire _26324 = _17499 ^ _5344;
  wire _26325 = _3905 ^ _4632;
  wire _26326 = _26324 ^ _26325;
  wire _26327 = _26323 ^ _26326;
  wire _26328 = _26319 ^ _26327;
  wire _26329 = _26316 ^ _26328;
  wire _26330 = _26299 ^ _26329;
  wire _26331 = _26270 ^ _26330;
  wire _26332 = _6009 ^ _8483;
  wire _26333 = _7277 ^ _769;
  wire _26334 = _22731 ^ _13991;
  wire _26335 = _26333 ^ _26334;
  wire _26336 = _26332 ^ _26335;
  wire _26337 = uncoded_block[1568] ^ uncoded_block[1573];
  wire _26338 = _26337 ^ _6663;
  wire _26339 = _11838 ^ _10172;
  wire _26340 = _26338 ^ _26339;
  wire _26341 = uncoded_block[1590] ^ uncoded_block[1596];
  wire _26342 = _26341 ^ _3934;
  wire _26343 = uncoded_block[1603] ^ uncoded_block[1607];
  wire _26344 = _26343 ^ _3154;
  wire _26345 = _26342 ^ _26344;
  wire _26346 = _26340 ^ _26345;
  wire _26347 = _26336 ^ _26346;
  wire _26348 = _804 ^ _6684;
  wire _26349 = _24114 ^ _26348;
  wire _26350 = _16529 ^ _12949;
  wire _26351 = _2408 ^ _2412;
  wire _26352 = _26350 ^ _26351;
  wire _26353 = _26349 ^ _26352;
  wire _26354 = uncoded_block[1659] ^ uncoded_block[1663];
  wire _26355 = _3174 ^ _26354;
  wire _26356 = uncoded_block[1664] ^ uncoded_block[1668];
  wire _26357 = _26356 ^ _8521;
  wire _26358 = _26355 ^ _26357;
  wire _26359 = uncoded_block[1677] ^ uncoded_block[1683];
  wire _26360 = _26359 ^ _14543;
  wire _26361 = _17037 ^ _26360;
  wire _26362 = _26358 ^ _26361;
  wire _26363 = _26353 ^ _26362;
  wire _26364 = _26347 ^ _26363;
  wire _26365 = uncoded_block[1691] ^ uncoded_block[1695];
  wire _26366 = _10205 ^ _26365;
  wire _26367 = _5409 ^ _3973;
  wire _26368 = _26366 ^ _26367;
  wire _26369 = uncoded_block[1712] ^ uncoded_block[1716];
  wire _26370 = _1672 ^ _26369;
  wire _26371 = _24138 ^ _26370;
  wire _26372 = _26368 ^ _26371;
  wire _26373 = _2443 ^ _12976;
  wire _26374 = _26373 ^ uncoded_block[1722];
  wire _26375 = _26372 ^ _26374;
  wire _26376 = _26364 ^ _26375;
  wire _26377 = _26331 ^ _26376;
  wire _26378 = _26207 ^ _26377;
  wire _26379 = _18057 ^ _14560;
  wire _26380 = _24148 ^ _26379;
  wire _26381 = uncoded_block[17] ^ uncoded_block[23];
  wire _26382 = _26381 ^ _9694;
  wire _26383 = _21412 ^ _875;
  wire _26384 = _26382 ^ _26383;
  wire _26385 = _26380 ^ _26384;
  wire _26386 = _16 ^ _8549;
  wire _26387 = _7965 ^ _15594;
  wire _26388 = _26386 ^ _26387;
  wire _26389 = _19505 ^ _21419;
  wire _26390 = _26388 ^ _26389;
  wire _26391 = _26385 ^ _26390;
  wire _26392 = _7365 ^ _1706;
  wire _26393 = uncoded_block[70] ^ uncoded_block[73];
  wire _26394 = _35 ^ _26393;
  wire _26395 = _26392 ^ _26394;
  wire _26396 = _4020 ^ _2481;
  wire _26397 = _26396 ^ _4736;
  wire _26398 = _26395 ^ _26397;
  wire _26399 = _14586 ^ _18077;
  wire _26400 = _8566 ^ _21888;
  wire _26401 = _26399 ^ _26400;
  wire _26402 = _15097 ^ _19025;
  wire _26403 = _911 ^ _19520;
  wire _26404 = _26402 ^ _26403;
  wire _26405 = _26401 ^ _26404;
  wire _26406 = _26398 ^ _26405;
  wire _26407 = _26391 ^ _26406;
  wire _26408 = _3253 ^ _9721;
  wire _26409 = _10821 ^ _57;
  wire _26410 = _26408 ^ _26409;
  wire _26411 = _4754 ^ _9177;
  wire _26412 = _4760 ^ _1744;
  wire _26413 = _26411 ^ _26412;
  wire _26414 = _26410 ^ _26413;
  wire _26415 = uncoded_block[151] ^ uncoded_block[155];
  wire _26416 = _26415 ^ _73;
  wire _26417 = _6785 ^ _11928;
  wire _26418 = _26416 ^ _26417;
  wire _26419 = uncoded_block[172] ^ uncoded_block[181];
  wire _26420 = _26419 ^ _13583;
  wire _26421 = _20493 ^ _26420;
  wire _26422 = _26418 ^ _26421;
  wire _26423 = _26414 ^ _26422;
  wire _26424 = _1759 ^ _18111;
  wire _26425 = _3283 ^ _8018;
  wire _26426 = _26424 ^ _26425;
  wire _26427 = _8021 ^ _5489;
  wire _26428 = _26427 ^ _16617;
  wire _26429 = _26426 ^ _26428;
  wire _26430 = _6169 ^ _967;
  wire _26431 = _106 ^ _26430;
  wire _26432 = _10289 ^ _7425;
  wire _26433 = _4797 ^ _8616;
  wire _26434 = _26432 ^ _26433;
  wire _26435 = _26431 ^ _26434;
  wire _26436 = _26429 ^ _26435;
  wire _26437 = _26423 ^ _26436;
  wire _26438 = _26407 ^ _26437;
  wire _26439 = _13053 ^ _15656;
  wire _26440 = _11955 ^ _26439;
  wire _26441 = uncoded_block[257] ^ uncoded_block[261];
  wire _26442 = _26441 ^ _4096;
  wire _26443 = _6188 ^ _7440;
  wire _26444 = _26442 ^ _26443;
  wire _26445 = _26440 ^ _26444;
  wire _26446 = _7441 ^ _5512;
  wire _26447 = uncoded_block[279] ^ uncoded_block[282];
  wire _26448 = _5513 ^ _26447;
  wire _26449 = _26446 ^ _26448;
  wire _26450 = _19072 ^ _9226;
  wire _26451 = _16144 ^ _2577;
  wire _26452 = _26450 ^ _26451;
  wire _26453 = _26449 ^ _26452;
  wire _26454 = _26445 ^ _26453;
  wire _26455 = _22400 ^ _1004;
  wire _26456 = _15671 ^ _11439;
  wire _26457 = _4832 ^ _11441;
  wire _26458 = _26456 ^ _26457;
  wire _26459 = _26455 ^ _26458;
  wire _26460 = _4123 ^ _1014;
  wire _26461 = uncoded_block[331] ^ uncoded_block[335];
  wire _26462 = _26461 ^ _7463;
  wire _26463 = _26460 ^ _26462;
  wire _26464 = _9242 ^ _2595;
  wire _26465 = _7465 ^ _4132;
  wire _26466 = _26464 ^ _26465;
  wire _26467 = _26463 ^ _26466;
  wire _26468 = _26459 ^ _26467;
  wire _26469 = _26454 ^ _26468;
  wire _26470 = uncoded_block[355] ^ uncoded_block[360];
  wire _26471 = _26470 ^ _21030;
  wire _26472 = _26471 ^ _13636;
  wire _26473 = _6873 ^ _20056;
  wire _26474 = _13101 ^ _19599;
  wire _26475 = _26473 ^ _26474;
  wire _26476 = _26472 ^ _26475;
  wire _26477 = _3381 ^ _3383;
  wire _26478 = uncoded_block[398] ^ uncoded_block[400];
  wire _26479 = _3384 ^ _26478;
  wire _26480 = _26477 ^ _26479;
  wire _26481 = uncoded_block[406] ^ uncoded_block[411];
  wire _26482 = _4156 ^ _26481;
  wire _26483 = _1054 ^ _8092;
  wire _26484 = _26482 ^ _26483;
  wire _26485 = _26480 ^ _26484;
  wire _26486 = _26476 ^ _26485;
  wire _26487 = _6249 ^ _194;
  wire _26488 = _11479 ^ _198;
  wire _26489 = _26487 ^ _26488;
  wire _26490 = _2638 ^ _4169;
  wire _26491 = uncoded_block[446] ^ uncoded_block[453];
  wire _26492 = _1863 ^ _26491;
  wire _26493 = _26490 ^ _26492;
  wire _26494 = _26489 ^ _26493;
  wire _26495 = uncoded_block[456] ^ uncoded_block[458];
  wire _26496 = _2650 ^ _26495;
  wire _26497 = _13662 ^ _8683;
  wire _26498 = _26496 ^ _26497;
  wire _26499 = _13665 ^ _4188;
  wire _26500 = uncoded_block[480] ^ uncoded_block[484];
  wire _26501 = _5592 ^ _26500;
  wire _26502 = _26499 ^ _26501;
  wire _26503 = _26498 ^ _26502;
  wire _26504 = _26494 ^ _26503;
  wire _26505 = _26486 ^ _26504;
  wire _26506 = _26469 ^ _26505;
  wire _26507 = _26438 ^ _26506;
  wire _26508 = _8116 ^ _22443;
  wire _26509 = _5608 ^ _5612;
  wire _26510 = _26508 ^ _26509;
  wire _26511 = _13676 ^ _4910;
  wire _26512 = _3444 ^ _4210;
  wire _26513 = _26511 ^ _26512;
  wire _26514 = uncoded_block[526] ^ uncoded_block[530];
  wire _26515 = _26514 ^ _18208;
  wire _26516 = _243 ^ _6293;
  wire _26517 = _26515 ^ _26516;
  wire _26518 = _26513 ^ _26517;
  wire _26519 = _26510 ^ _26518;
  wire _26520 = _16715 ^ _2687;
  wire _26521 = _5630 ^ _8724;
  wire _26522 = _26520 ^ _26521;
  wire _26523 = _8139 ^ _9319;
  wire _26524 = _9320 ^ _6309;
  wire _26525 = _26523 ^ _26524;
  wire _26526 = _26522 ^ _26525;
  wire _26527 = _17221 ^ _1133;
  wire _26528 = uncoded_block[582] ^ uncoded_block[588];
  wire _26529 = _26528 ^ _1141;
  wire _26530 = _26527 ^ _26529;
  wire _26531 = _2700 ^ _21565;
  wire _26532 = uncoded_block[601] ^ uncoded_block[605];
  wire _26533 = _4953 ^ _26532;
  wire _26534 = _26531 ^ _26533;
  wire _26535 = _26530 ^ _26534;
  wire _26536 = _26526 ^ _26535;
  wire _26537 = _26519 ^ _26536;
  wire _26538 = _4240 ^ _13176;
  wire _26539 = _7564 ^ _7568;
  wire _26540 = _26538 ^ _26539;
  wire _26541 = _7570 ^ _17238;
  wire _26542 = _22950 ^ _7577;
  wire _26543 = _26541 ^ _26542;
  wire _26544 = _26540 ^ _26543;
  wire _26545 = uncoded_block[637] ^ uncoded_block[639];
  wire _26546 = _26545 ^ _6336;
  wire _26547 = _3505 ^ _14234;
  wire _26548 = _26546 ^ _26547;
  wire _26549 = uncoded_block[656] ^ uncoded_block[658];
  wire _26550 = _26549 ^ _1173;
  wire _26551 = _4976 ^ _26550;
  wire _26552 = _26548 ^ _26551;
  wire _26553 = _26544 ^ _26552;
  wire _26554 = _4265 ^ _8761;
  wire _26555 = _12636 ^ _15281;
  wire _26556 = _26554 ^ _26555;
  wire _26557 = uncoded_block[687] ^ uncoded_block[690];
  wire _26558 = uncoded_block[691] ^ uncoded_block[700];
  wire _26559 = _26557 ^ _26558;
  wire _26560 = _4990 ^ _10447;
  wire _26561 = _26559 ^ _26560;
  wire _26562 = _26556 ^ _26561;
  wire _26563 = _336 ^ _4996;
  wire _26564 = _2762 ^ _12647;
  wire _26565 = _26563 ^ _26564;
  wire _26566 = uncoded_block[727] ^ uncoded_block[733];
  wire _26567 = _1987 ^ _26566;
  wire _26568 = _17763 ^ _26567;
  wire _26569 = _26565 ^ _26568;
  wire _26570 = _26562 ^ _26569;
  wire _26571 = _26553 ^ _26570;
  wire _26572 = _26537 ^ _26571;
  wire _26573 = _1203 ^ _1206;
  wire _26574 = _26573 ^ _24330;
  wire _26575 = _5702 ^ _8778;
  wire _26576 = _7013 ^ _15305;
  wire _26577 = _26575 ^ _26576;
  wire _26578 = _26574 ^ _26577;
  wire _26579 = uncoded_block[758] ^ uncoded_block[761];
  wire _26580 = _26579 ^ _18740;
  wire _26581 = _11018 ^ _12114;
  wire _26582 = _26580 ^ _26581;
  wire _26583 = _20165 ^ _13219;
  wire _26584 = _26583 ^ _18747;
  wire _26585 = _26582 ^ _26584;
  wire _26586 = _26578 ^ _26585;
  wire _26587 = _5033 ^ _4314;
  wire _26588 = uncoded_block[794] ^ uncoded_block[798];
  wire _26589 = uncoded_block[801] ^ uncoded_block[803];
  wire _26590 = _26588 ^ _26589;
  wire _26591 = _26587 ^ _26590;
  wire _26592 = _389 ^ _5041;
  wire _26593 = _5042 ^ _2808;
  wire _26594 = _26592 ^ _26593;
  wire _26595 = _26591 ^ _26594;
  wire _26596 = _22525 ^ _14290;
  wire _26597 = _1247 ^ _7039;
  wire _26598 = _26596 ^ _26597;
  wire _26599 = _400 ^ _16801;
  wire _26600 = _4337 ^ _2815;
  wire _26601 = _26599 ^ _26600;
  wire _26602 = _26598 ^ _26601;
  wire _26603 = _26595 ^ _26602;
  wire _26604 = _26586 ^ _26603;
  wire _26605 = _5060 ^ _2821;
  wire _26606 = _8812 ^ _23010;
  wire _26607 = _26605 ^ _26606;
  wire _26608 = _413 ^ _7650;
  wire _26609 = _1266 ^ _5072;
  wire _26610 = _26608 ^ _26609;
  wire _26611 = _26607 ^ _26610;
  wire _26612 = _1269 ^ _417;
  wire _26613 = _7060 ^ _2836;
  wire _26614 = _26612 ^ _26613;
  wire _26615 = _9416 ^ _2061;
  wire _26616 = _3614 ^ _5758;
  wire _26617 = _26615 ^ _26616;
  wire _26618 = _26614 ^ _26617;
  wire _26619 = _26611 ^ _26618;
  wire _26620 = _6424 ^ _1280;
  wire _26621 = _5761 ^ _3629;
  wire _26622 = _26620 ^ _26621;
  wire _26623 = uncoded_block[924] ^ uncoded_block[928];
  wire _26624 = _26623 ^ _8835;
  wire _26625 = _3633 ^ _26624;
  wire _26626 = _26622 ^ _26625;
  wire _26627 = _8262 ^ _5101;
  wire _26628 = uncoded_block[938] ^ uncoded_block[942];
  wire _26629 = _26628 ^ _1302;
  wire _26630 = _26627 ^ _26629;
  wire _26631 = _460 ^ _5779;
  wire _26632 = _10525 ^ _5107;
  wire _26633 = _26631 ^ _26632;
  wire _26634 = _26630 ^ _26633;
  wire _26635 = _26626 ^ _26634;
  wire _26636 = _26619 ^ _26635;
  wire _26637 = _26604 ^ _26636;
  wire _26638 = _26572 ^ _26637;
  wire _26639 = _26507 ^ _26638;
  wire _26640 = _14845 ^ _7092;
  wire _26641 = _8853 ^ _3659;
  wire _26642 = uncoded_block[986] ^ uncoded_block[992];
  wire _26643 = _26642 ^ _7097;
  wire _26644 = _26641 ^ _26643;
  wire _26645 = _26640 ^ _26644;
  wire _26646 = uncoded_block[1007] ^ uncoded_block[1011];
  wire _26647 = _26646 ^ _9996;
  wire _26648 = _25757 ^ _26647;
  wire _26649 = _2893 ^ _5135;
  wire _26650 = _26649 ^ _8302;
  wire _26651 = _26648 ^ _26650;
  wire _26652 = _26645 ^ _26651;
  wire _26653 = uncoded_block[1031] ^ uncoded_block[1036];
  wire _26654 = _2898 ^ _26653;
  wire _26655 = _26654 ^ _2131;
  wire _26656 = _3681 ^ _10564;
  wire _26657 = _12764 ^ _13849;
  wire _26658 = _26656 ^ _26657;
  wire _26659 = _26655 ^ _26658;
  wire _26660 = _3685 ^ _9475;
  wire _26661 = uncoded_block[1071] ^ uncoded_block[1074];
  wire _26662 = _26661 ^ _8895;
  wire _26663 = _26660 ^ _26662;
  wire _26664 = uncoded_block[1079] ^ uncoded_block[1086];
  wire _26665 = _26664 ^ _2149;
  wire _26666 = _26665 ^ _23509;
  wire _26667 = _26663 ^ _26666;
  wire _26668 = _26659 ^ _26667;
  wire _26669 = _26652 ^ _26668;
  wire _26670 = _11140 ^ _10581;
  wire _26671 = uncoded_block[1110] ^ uncoded_block[1115];
  wire _26672 = _14372 ^ _26671;
  wire _26673 = _13322 ^ _2942;
  wire _26674 = _26672 ^ _26673;
  wire _26675 = _26670 ^ _26674;
  wire _26676 = _5854 ^ _2945;
  wire _26677 = _18834 ^ _3721;
  wire _26678 = _26676 ^ _26677;
  wire _26679 = uncoded_block[1143] ^ uncoded_block[1150];
  wire _26680 = _26679 ^ _8937;
  wire _26681 = _26680 ^ _11712;
  wire _26682 = _26678 ^ _26681;
  wire _26683 = _26675 ^ _26682;
  wire _26684 = _6511 ^ _4476;
  wire _26685 = _5870 ^ _3739;
  wire _26686 = _26684 ^ _26685;
  wire _26687 = _589 ^ _2195;
  wire _26688 = _5200 ^ _9508;
  wire _26689 = _26687 ^ _26688;
  wire _26690 = _26686 ^ _26689;
  wire _26691 = _5203 ^ _2203;
  wire _26692 = _26691 ^ _2208;
  wire _26693 = _16399 ^ _5209;
  wire _26694 = uncoded_block[1211] ^ uncoded_block[1212];
  wire _26695 = _26694 ^ _605;
  wire _26696 = _26693 ^ _26695;
  wire _26697 = _26692 ^ _26696;
  wire _26698 = _26690 ^ _26697;
  wire _26699 = _26683 ^ _26698;
  wire _26700 = _26669 ^ _26699;
  wire _26701 = _606 ^ _608;
  wire _26702 = _1435 ^ _612;
  wire _26703 = _26701 ^ _26702;
  wire _26704 = uncoded_block[1228] ^ uncoded_block[1233];
  wire _26705 = _26704 ^ _2989;
  wire _26706 = _2230 ^ _10627;
  wire _26707 = _26705 ^ _26706;
  wire _26708 = _26703 ^ _26707;
  wire _26709 = uncoded_block[1252] ^ uncoded_block[1256];
  wire _26710 = _621 ^ _26709;
  wire _26711 = _25815 ^ _26710;
  wire _26712 = uncoded_block[1260] ^ uncoded_block[1263];
  wire _26713 = _7780 ^ _26712;
  wire _26714 = _9532 ^ _2245;
  wire _26715 = _26713 ^ _26714;
  wire _26716 = _26711 ^ _26715;
  wire _26717 = _26708 ^ _26716;
  wire _26718 = uncoded_block[1272] ^ uncoded_block[1274];
  wire _26719 = _26718 ^ _7792;
  wire _26720 = _3793 ^ _4525;
  wire _26721 = _26719 ^ _26720;
  wire _26722 = _6560 ^ _4529;
  wire _26723 = _26722 ^ _11755;
  wire _26724 = _26721 ^ _26723;
  wire _26725 = _645 ^ _14939;
  wire _26726 = uncoded_block[1314] ^ uncoded_block[1318];
  wire _26727 = _13917 ^ _26726;
  wire _26728 = _26725 ^ _26727;
  wire _26729 = uncoded_block[1324] ^ uncoded_block[1329];
  wire _26730 = _654 ^ _26729;
  wire _26731 = _8413 ^ _9563;
  wire _26732 = _26730 ^ _26731;
  wire _26733 = _26728 ^ _26732;
  wire _26734 = _26724 ^ _26733;
  wire _26735 = _26717 ^ _26734;
  wire _26736 = uncoded_block[1339] ^ uncoded_block[1344];
  wire _26737 = _26736 ^ _1501;
  wire _26738 = _5269 ^ _672;
  wire _26739 = _26737 ^ _26738;
  wire _26740 = _2283 ^ _10101;
  wire _26741 = _6589 ^ _26740;
  wire _26742 = _26739 ^ _26741;
  wire _26743 = uncoded_block[1377] ^ uncoded_block[1380];
  wire _26744 = _11226 ^ _26743;
  wire _26745 = _687 ^ _5950;
  wire _26746 = _26744 ^ _26745;
  wire _26747 = uncoded_block[1397] ^ uncoded_block[1400];
  wire _26748 = _6597 ^ _26747;
  wire _26749 = uncoded_block[1401] ^ uncoded_block[1404];
  wire _26750 = _26749 ^ _3847;
  wire _26751 = _26748 ^ _26750;
  wire _26752 = _26746 ^ _26751;
  wire _26753 = _26742 ^ _26752;
  wire _26754 = uncoded_block[1416] ^ uncoded_block[1419];
  wire _26755 = _3069 ^ _26754;
  wire _26756 = _9586 ^ _26755;
  wire _26757 = _16463 ^ _3074;
  wire _26758 = _2308 ^ _9591;
  wire _26759 = _26757 ^ _26758;
  wire _26760 = _26756 ^ _26759;
  wire _26761 = uncoded_block[1435] ^ uncoded_block[1439];
  wire _26762 = _26761 ^ _4590;
  wire _26763 = uncoded_block[1447] ^ uncoded_block[1450];
  wire _26764 = _5970 ^ _26763;
  wire _26765 = _26762 ^ _26764;
  wire _26766 = _9037 ^ _8455;
  wire _26767 = _22250 ^ _26766;
  wire _26768 = _26765 ^ _26767;
  wire _26769 = _26760 ^ _26768;
  wire _26770 = _26753 ^ _26769;
  wire _26771 = _26735 ^ _26770;
  wire _26772 = _26700 ^ _26771;
  wire _26773 = uncoded_block[1469] ^ uncoded_block[1474];
  wire _26774 = _5314 ^ _26773;
  wire _26775 = _25423 ^ _4607;
  wire _26776 = _26774 ^ _26775;
  wire _26777 = _5988 ^ _17980;
  wire _26778 = _3103 ^ _9614;
  wire _26779 = _26777 ^ _26778;
  wire _26780 = _26776 ^ _26779;
  wire _26781 = _743 ^ _6635;
  wire _26782 = _7259 ^ _24539;
  wire _26783 = _26781 ^ _26782;
  wire _26784 = uncoded_block[1524] ^ uncoded_block[1529];
  wire _26785 = _26784 ^ _6647;
  wire _26786 = _9056 ^ _26785;
  wire _26787 = _26783 ^ _26786;
  wire _26788 = _26780 ^ _26787;
  wire _26789 = _12914 ^ _6648;
  wire _26790 = _1587 ^ _5350;
  wire _26791 = _26789 ^ _26790;
  wire _26792 = uncoded_block[1545] ^ uncoded_block[1549];
  wire _26793 = _26792 ^ _767;
  wire _26794 = uncoded_block[1560] ^ uncoded_block[1562];
  wire _26795 = _770 ^ _26794;
  wire _26796 = _26793 ^ _26795;
  wire _26797 = _26791 ^ _26796;
  wire _26798 = _5361 ^ _11833;
  wire _26799 = _5363 ^ _4647;
  wire _26800 = _26798 ^ _26799;
  wire _26801 = uncoded_block[1577] ^ uncoded_block[1581];
  wire _26802 = _4648 ^ _26801;
  wire _26803 = _26802 ^ _7899;
  wire _26804 = _26800 ^ _26803;
  wire _26805 = _26797 ^ _26804;
  wire _26806 = _26788 ^ _26805;
  wire _26807 = _3146 ^ _6673;
  wire _26808 = uncoded_block[1597] ^ uncoded_block[1601];
  wire _26809 = _26808 ^ _3153;
  wire _26810 = _26807 ^ _26809;
  wire _26811 = _11303 ^ _1632;
  wire _26812 = uncoded_block[1617] ^ uncoded_block[1623];
  wire _26813 = _26812 ^ _6046;
  wire _26814 = _26811 ^ _26813;
  wire _26815 = _26810 ^ _26814;
  wire _26816 = _3161 ^ _7914;
  wire _26817 = _9659 ^ _7308;
  wire _26818 = _26816 ^ _26817;
  wire _26819 = _6689 ^ _18516;
  wire _26820 = _1649 ^ _3172;
  wire _26821 = _26819 ^ _26820;
  wire _26822 = _26818 ^ _26821;
  wire _26823 = _26815 ^ _26822;
  wire _26824 = _18030 ^ _12957;
  wire _26825 = _26824 ^ _18036;
  wire _26826 = _3962 ^ _833;
  wire _26827 = _11320 ^ _26826;
  wire _26828 = _26825 ^ _26827;
  wire _26829 = _3965 ^ _7935;
  wire _26830 = _3968 ^ _3972;
  wire _26831 = _26829 ^ _26830;
  wire _26832 = uncoded_block[1701] ^ uncoded_block[1704];
  wire _26833 = _11327 ^ _26832;
  wire _26834 = _8536 ^ _851;
  wire _26835 = _26833 ^ _26834;
  wire _26836 = _26831 ^ _26835;
  wire _26837 = _26828 ^ _26836;
  wire _26838 = _26823 ^ _26837;
  wire _26839 = _26806 ^ _26838;
  wire _26840 = _22316 ^ _1677;
  wire _26841 = _26840 ^ uncoded_block[1721];
  wire _26842 = _26839 ^ _26841;
  wire _26843 = _26772 ^ _26842;
  wire _26844 = _26639 ^ _26843;
  wire _26845 = _19001 ^ _3217;
  wire _26846 = _25936 ^ _26845;
  wire _26847 = _6095 ^ _19501;
  wire _26848 = _7354 ^ _26847;
  wire _26849 = _26846 ^ _26848;
  wire _26850 = uncoded_block[43] ^ uncoded_block[48];
  wire _26851 = _4008 ^ _26850;
  wire _26852 = _26851 ^ _10236;
  wire _26853 = _7364 ^ _2474;
  wire _26854 = _25950 ^ _19511;
  wire _26855 = _26853 ^ _26854;
  wire _26856 = _26852 ^ _26855;
  wire _26857 = _26849 ^ _26856;
  wire _26858 = _25955 ^ _6754;
  wire _26859 = _26858 ^ _25960;
  wire _26860 = _25961 ^ _25964;
  wire _26861 = _26859 ^ _26860;
  wire _26862 = _25965 ^ _25968;
  wire _26863 = _4754 ^ _20963;
  wire _26864 = _3265 ^ _6138;
  wire _26865 = _26863 ^ _26864;
  wire _26866 = _26862 ^ _26865;
  wire _26867 = _26861 ^ _26866;
  wire _26868 = _26857 ^ _26867;
  wire _26869 = _1742 ^ _3268;
  wire _26870 = _3269 ^ _1748;
  wire _26871 = _26869 ^ _26870;
  wire _26872 = _11390 ^ _2521;
  wire _26873 = _20979 ^ _13034;
  wire _26874 = _26872 ^ _26873;
  wire _26875 = _26871 ^ _26874;
  wire _26876 = _6798 ^ _6800;
  wire _26877 = _15132 ^ _26876;
  wire _26878 = _4779 ^ _14101;
  wire _26879 = _955 ^ _2540;
  wire _26880 = _26878 ^ _26879;
  wire _26881 = _26877 ^ _26880;
  wire _26882 = _26875 ^ _26881;
  wire _26883 = _3296 ^ _3298;
  wire _26884 = _24657 ^ _16125;
  wire _26885 = _26883 ^ _26884;
  wire _26886 = uncoded_block[236] ^ uncoded_block[244];
  wire _26887 = _24660 ^ _26886;
  wire _26888 = _8617 ^ _7434;
  wire _26889 = _26887 ^ _26888;
  wire _26890 = _26885 ^ _26889;
  wire _26891 = _11419 ^ _23746;
  wire _26892 = _119 ^ _6185;
  wire _26893 = _26891 ^ _26892;
  wire _26894 = _20523 ^ _128;
  wire _26895 = uncoded_block[274] ^ uncoded_block[278];
  wire _26896 = _26895 ^ _7446;
  wire _26897 = _26894 ^ _26896;
  wire _26898 = _26893 ^ _26897;
  wire _26899 = _26890 ^ _26898;
  wire _26900 = _26882 ^ _26899;
  wire _26901 = _26868 ^ _26900;
  wire _26902 = _8632 ^ _992;
  wire _26903 = _10876 ^ _8633;
  wire _26904 = _26902 ^ _26903;
  wire _26905 = uncoded_block[304] ^ uncoded_block[313];
  wire _26906 = _26905 ^ _3340;
  wire _26907 = _13616 ^ _26906;
  wire _26908 = _26904 ^ _26907;
  wire _26909 = _13624 ^ _1818;
  wire _26910 = _4123 ^ _26021;
  wire _26911 = _26909 ^ _26910;
  wire _26912 = _26911 ^ _26029;
  wire _26913 = _26908 ^ _26912;
  wire _26914 = _5541 ^ _19092;
  wire _26915 = _6221 ^ _2606;
  wire _26916 = _26914 ^ _26915;
  wire _26917 = _7470 ^ _1835;
  wire _26918 = _1838 ^ _4853;
  wire _26919 = _26917 ^ _26918;
  wire _26920 = _26916 ^ _26919;
  wire _26921 = _4143 ^ _3377;
  wire _26922 = _13102 ^ _12541;
  wire _26923 = _26921 ^ _26922;
  wire _26924 = _4152 ^ _3384;
  wire _26925 = uncoded_block[401] ^ uncoded_block[404];
  wire _26926 = _26478 ^ _26925;
  wire _26927 = _26924 ^ _26926;
  wire _26928 = _26923 ^ _26927;
  wire _26929 = _26920 ^ _26928;
  wire _26930 = _26913 ^ _26929;
  wire _26931 = _191 ^ _1055;
  wire _26932 = _14680 ^ _26931;
  wire _26933 = _11476 ^ _4163;
  wire _26934 = _4164 ^ _2633;
  wire _26935 = _26933 ^ _26934;
  wire _26936 = _26932 ^ _26935;
  wire _26937 = _13115 ^ _13117;
  wire _26938 = _26937 ^ _8677;
  wire _26939 = _26056 ^ _26058;
  wire _26940 = _26938 ^ _26939;
  wire _26941 = _26936 ^ _26940;
  wire _26942 = _4181 ^ _11491;
  wire _26943 = _26059 ^ _26942;
  wire _26944 = uncoded_block[470] ^ uncoded_block[473];
  wire _26945 = _9283 ^ _26944;
  wire _26946 = _11494 ^ _24723;
  wire _26947 = _26945 ^ _26946;
  wire _26948 = _26943 ^ _26947;
  wire _26949 = _5593 ^ _4194;
  wire _26950 = _10937 ^ _13139;
  wire _26951 = _26949 ^ _26950;
  wire _26952 = _4905 ^ _3434;
  wire _26953 = _2668 ^ _12034;
  wire _26954 = _26952 ^ _26953;
  wire _26955 = _26951 ^ _26954;
  wire _26956 = _26948 ^ _26955;
  wire _26957 = _26941 ^ _26956;
  wire _26958 = _26930 ^ _26957;
  wire _26959 = _26901 ^ _26958;
  wire _26960 = _231 ^ _9295;
  wire _26961 = _10945 ^ _3444;
  wire _26962 = _26960 ^ _26961;
  wire _26963 = _3445 ^ _20099;
  wire _26964 = _26081 ^ _6932;
  wire _26965 = _26963 ^ _26964;
  wire _26966 = _26962 ^ _26965;
  wire _26967 = _4217 ^ _5628;
  wire _26968 = _26967 ^ _8722;
  wire _26969 = _1123 ^ _26090;
  wire _26970 = _1126 ^ _4223;
  wire _26971 = _26969 ^ _26970;
  wire _26972 = _26968 ^ _26971;
  wire _26973 = _26966 ^ _26972;
  wire _26974 = _4224 ^ _11526;
  wire _26975 = _6947 ^ _2696;
  wire _26976 = _26974 ^ _26975;
  wire _26977 = _26096 ^ _2700;
  wire _26978 = _6316 ^ _6952;
  wire _26979 = _26977 ^ _26978;
  wire _26980 = _26976 ^ _26979;
  wire _26981 = _3486 ^ _15757;
  wire _26982 = _12609 ^ _1149;
  wire _26983 = _26981 ^ _26982;
  wire _26984 = _20125 ^ _5658;
  wire _26985 = _26108 ^ _4249;
  wire _26986 = _26984 ^ _26985;
  wire _26987 = _26983 ^ _26986;
  wire _26988 = _26980 ^ _26987;
  wire _26989 = _26973 ^ _26988;
  wire _26990 = _4255 ^ _2727;
  wire _26991 = _26990 ^ _26113;
  wire _26992 = _26991 ^ _26116;
  wire _26993 = _1177 ^ _19185;
  wire _26994 = _26118 ^ _26993;
  wire _26995 = uncoded_block[679] ^ uncoded_block[683];
  wire _26996 = _8177 ^ _26995;
  wire _26997 = _15281 ^ _1974;
  wire _26998 = _26996 ^ _26997;
  wire _26999 = _26994 ^ _26998;
  wire _27000 = _26992 ^ _26999;
  wire _27001 = _26563 ^ _16766;
  wire _27002 = _26126 ^ _27001;
  wire _27003 = _17762 ^ _8198;
  wire _27004 = _3544 ^ _4286;
  wire _27005 = _27003 ^ _27004;
  wire _27006 = _23870 ^ _3550;
  wire _27007 = _2775 ^ _2777;
  wire _27008 = _27006 ^ _27007;
  wire _27009 = _27005 ^ _27008;
  wire _27010 = _27002 ^ _27009;
  wire _27011 = _27000 ^ _27010;
  wire _27012 = _26989 ^ _27011;
  wire _27013 = _8779 ^ _3559;
  wire _27014 = _8781 ^ _1217;
  wire _27015 = _27013 ^ _27014;
  wire _27016 = _1221 ^ _5711;
  wire _27017 = uncoded_block[776] ^ uncoded_block[779];
  wire _27018 = _27017 ^ _3568;
  wire _27019 = _27016 ^ _27018;
  wire _27020 = _27015 ^ _27019;
  wire _27021 = _371 ^ _5032;
  wire _27022 = _1225 ^ _11024;
  wire _27023 = _27021 ^ _27022;
  wire _27024 = _7029 ^ _26589;
  wire _27025 = _3581 ^ _11596;
  wire _27026 = _27024 ^ _27025;
  wire _27027 = _27023 ^ _27026;
  wire _27028 = _27020 ^ _27027;
  wire _27029 = _9397 ^ _1242;
  wire _27030 = _5051 ^ _398;
  wire _27031 = _27029 ^ _27030;
  wire _27032 = _401 ^ _14809;
  wire _27033 = _27032 ^ _26162;
  wire _27034 = _27031 ^ _27033;
  wire _27035 = _14814 ^ _8237;
  wire _27036 = _15330 ^ _6410;
  wire _27037 = _27035 ^ _27036;
  wire _27038 = _413 ^ _26171;
  wire _27039 = _27038 ^ _13792;
  wire _27040 = _27037 ^ _27039;
  wire _27041 = _27034 ^ _27040;
  wire _27042 = _27028 ^ _27041;
  wire _27043 = _25719 ^ _2835;
  wire _27044 = _2836 ^ _423;
  wire _27045 = _27043 ^ _27044;
  wire _27046 = uncoded_block[887] ^ uncoded_block[890];
  wire _27047 = _27046 ^ _5083;
  wire _27048 = uncoded_block[895] ^ uncoded_block[899];
  wire _27049 = _27048 ^ _429;
  wire _27050 = _27047 ^ _27049;
  wire _27051 = _27045 ^ _27050;
  wire _27052 = _2065 ^ _431;
  wire _27053 = _19252 ^ _17820;
  wire _27054 = _27052 ^ _27053;
  wire _27055 = _448 ^ _1299;
  wire _27056 = _452 ^ _455;
  wire _27057 = _27055 ^ _27056;
  wire _27058 = _27054 ^ _27057;
  wire _27059 = _27051 ^ _27058;
  wire _27060 = _5777 ^ _8274;
  wire _27061 = _461 ^ _2090;
  wire _27062 = _27060 ^ _27061;
  wire _27063 = _4385 ^ _3653;
  wire _27064 = _2093 ^ _1315;
  wire _27065 = _27063 ^ _27064;
  wire _27066 = _27062 ^ _27065;
  wire _27067 = _5790 ^ _6451;
  wire _27068 = _11093 ^ _27067;
  wire _27069 = _23940 ^ _13278;
  wire _27070 = _27068 ^ _27069;
  wire _27071 = _27066 ^ _27070;
  wire _27072 = _27059 ^ _27071;
  wire _27073 = _27042 ^ _27072;
  wire _27074 = _27012 ^ _27073;
  wire _27075 = _26959 ^ _27074;
  wire _27076 = _5798 ^ _2114;
  wire _27077 = uncoded_block[1007] ^ uncoded_block[1010];
  wire _27078 = _27077 ^ _8296;
  wire _27079 = _27076 ^ _27078;
  wire _27080 = _7703 ^ _5137;
  wire _27081 = uncoded_block[1025] ^ uncoded_block[1029];
  wire _27082 = _27081 ^ _2907;
  wire _27083 = _27080 ^ _27082;
  wire _27084 = _27079 ^ _27083;
  wire _27085 = uncoded_block[1036] ^ uncoded_block[1042];
  wire _27086 = _27085 ^ _2130;
  wire _27087 = _8309 ^ _15871;
  wire _27088 = _27086 ^ _27087;
  wire _27089 = uncoded_block[1058] ^ uncoded_block[1066];
  wire _27090 = _519 ^ _27089;
  wire _27091 = _5828 ^ _21685;
  wire _27092 = _27090 ^ _27091;
  wire _27093 = _27088 ^ _27092;
  wire _27094 = _27084 ^ _27093;
  wire _27095 = _15883 ^ _12222;
  wire _27096 = _2935 ^ _26227;
  wire _27097 = _27095 ^ _27096;
  wire _27098 = _8915 ^ _2165;
  wire _27099 = _5175 ^ _23981;
  wire _27100 = _27098 ^ _27099;
  wire _27101 = _27097 ^ _27100;
  wire _27102 = _15896 ^ _8929;
  wire _27103 = _27102 ^ _569;
  wire _27104 = _26240 ^ _9500;
  wire _27105 = uncoded_block[1158] ^ uncoded_block[1163];
  wire _27106 = _27105 ^ _5193;
  wire _27107 = _27104 ^ _27106;
  wire _27108 = _27103 ^ _27107;
  wire _27109 = _27101 ^ _27108;
  wire _27110 = _27094 ^ _27109;
  wire _27111 = uncoded_block[1171] ^ uncoded_block[1176];
  wire _27112 = _11160 ^ _27111;
  wire _27113 = uncoded_block[1180] ^ uncoded_block[1184];
  wire _27114 = _4481 ^ _27113;
  wire _27115 = _27112 ^ _27114;
  wire _27116 = uncoded_block[1185] ^ uncoded_block[1187];
  wire _27117 = _27116 ^ _3747;
  wire _27118 = _3749 ^ _1421;
  wire _27119 = _27117 ^ _27118;
  wire _27120 = _27115 ^ _27119;
  wire _27121 = _2206 ^ _2974;
  wire _27122 = _2216 ^ _1427;
  wire _27123 = _27121 ^ _27122;
  wire _27124 = _4498 ^ _10061;
  wire _27125 = _11180 ^ _3771;
  wire _27126 = _27124 ^ _27125;
  wire _27127 = _27123 ^ _27126;
  wire _27128 = _27120 ^ _27127;
  wire _27129 = uncoded_block[1241] ^ uncoded_block[1243];
  wire _27130 = _16915 ^ _27129;
  wire _27131 = _13365 ^ _2232;
  wire _27132 = _27130 ^ _27131;
  wire _27133 = _27132 ^ _26264;
  wire _27134 = _628 ^ _7792;
  wire _27135 = _13371 ^ _27134;
  wire _27136 = _3793 ^ _23123;
  wire _27137 = _4526 ^ _641;
  wire _27138 = _27136 ^ _27137;
  wire _27139 = _27135 ^ _27138;
  wire _27140 = _27133 ^ _27139;
  wire _27141 = _27128 ^ _27140;
  wire _27142 = _27110 ^ _27141;
  wire _27143 = _10646 ^ _12843;
  wire _27144 = _2254 ^ _26276;
  wire _27145 = _27143 ^ _27144;
  wire _27146 = _1483 ^ _5926;
  wire _27147 = _27146 ^ _4544;
  wire _27148 = _27145 ^ _27147;
  wire _27149 = _656 ^ _1490;
  wire _27150 = _27149 ^ _19849;
  wire _27151 = uncoded_block[1340] ^ uncoded_block[1345];
  wire _27152 = _3822 ^ _27151;
  wire _27153 = _18434 ^ _18436;
  wire _27154 = _27152 ^ _27153;
  wire _27155 = _27150 ^ _27154;
  wire _27156 = _27148 ^ _27155;
  wire _27157 = uncoded_block[1360] ^ uncoded_block[1363];
  wire _27158 = _12857 ^ _27157;
  wire _27159 = _27158 ^ _12306;
  wire _27160 = uncoded_block[1377] ^ uncoded_block[1382];
  wire _27161 = _27160 ^ _10108;
  wire _27162 = _27161 ^ _18898;
  wire _27163 = _27159 ^ _27162;
  wire _27164 = _21774 ^ _5955;
  wire _27165 = _27164 ^ _4579;
  wire _27166 = _10113 ^ _4580;
  wire _27167 = _13422 ^ _2306;
  wire _27168 = _27166 ^ _27167;
  wire _27169 = _27165 ^ _27168;
  wire _27170 = _27163 ^ _27169;
  wire _27171 = _27156 ^ _27170;
  wire _27172 = _10684 ^ _1531;
  wire _27173 = _7843 ^ _27172;
  wire _27174 = _16962 ^ _15982;
  wire _27175 = uncoded_block[1441] ^ uncoded_block[1445];
  wire _27176 = _27175 ^ _26309;
  wire _27177 = _27174 ^ _27176;
  wire _27178 = _27173 ^ _27177;
  wire _27179 = _11247 ^ _723;
  wire _27180 = _8452 ^ _8455;
  wire _27181 = _27179 ^ _27180;
  wire _27182 = uncoded_block[1472] ^ uncoded_block[1478];
  wire _27183 = _22254 ^ _27182;
  wire _27184 = uncoded_block[1484] ^ uncoded_block[1487];
  wire _27185 = _27184 ^ _740;
  wire _27186 = _27183 ^ _27185;
  wire _27187 = _27181 ^ _27186;
  wire _27188 = _27178 ^ _27187;
  wire _27189 = _24536 ^ _7257;
  wire _27190 = _7260 ^ _26320;
  wire _27191 = _27189 ^ _27190;
  wire _27192 = _26321 ^ _1579;
  wire _27193 = _755 ^ _1582;
  wire _27194 = _27192 ^ _27193;
  wire _27195 = _9633 ^ _6009;
  wire _27196 = _27194 ^ _27195;
  wire _27197 = _27191 ^ _27196;
  wire _27198 = _27188 ^ _27197;
  wire _27199 = _27171 ^ _27198;
  wire _27200 = _27142 ^ _27199;
  wire _27201 = _8483 ^ _16997;
  wire _27202 = uncoded_block[1563] ^ uncoded_block[1568];
  wire _27203 = _18941 ^ _27202;
  wire _27204 = _14506 ^ _16513;
  wire _27205 = _27203 ^ _27204;
  wire _27206 = _27201 ^ _27205;
  wire _27207 = _10172 ^ _26341;
  wire _27208 = _3934 ^ _10742;
  wire _27209 = _27207 ^ _27208;
  wire _27210 = _3154 ^ _7908;
  wire _27211 = _6679 ^ _16032;
  wire _27212 = _27210 ^ _27211;
  wire _27213 = _27209 ^ _27212;
  wire _27214 = _27206 ^ _27213;
  wire _27215 = uncoded_block[1618] ^ uncoded_block[1621];
  wire _27216 = _27215 ^ _16529;
  wire _27217 = _12949 ^ _17527;
  wire _27218 = _27216 ^ _27217;
  wire _27219 = _1649 ^ _9106;
  wire _27220 = _27219 ^ _4681;
  wire _27221 = _27218 ^ _27220;
  wire _27222 = _1654 ^ _25476;
  wire _27223 = _6700 ^ _830;
  wire _27224 = _27222 ^ _27223;
  wire _27225 = _12398 ^ _13517;
  wire _27226 = _27225 ^ _16547;
  wire _27227 = _27224 ^ _27226;
  wire _27228 = _27221 ^ _27227;
  wire _27229 = _27214 ^ _27228;
  wire _27230 = _26365 ^ _5409;
  wire _27231 = _3973 ^ _24137;
  wire _27232 = _27230 ^ _27231;
  wire _27233 = _8535 ^ _1672;
  wire _27234 = _26369 ^ _2443;
  wire _27235 = _27233 ^ _27234;
  wire _27236 = _27232 ^ _27235;
  wire _27237 = _27236 ^ _12977;
  wire _27238 = _27229 ^ _27237;
  wire _27239 = _27200 ^ _27238;
  wire _27240 = _27075 ^ _27239;
  wire _27241 = uncoded_block[2] ^ uncoded_block[6];
  wire _27242 = _3209 ^ _27241;
  wire _27243 = _1684 ^ _14560;
  wire _27244 = _27242 ^ _27243;
  wire _27245 = uncoded_block[19] ^ uncoded_block[25];
  wire _27246 = _1687 ^ _27245;
  wire _27247 = _7959 ^ _5429;
  wire _27248 = _27246 ^ _27247;
  wire _27249 = _27244 ^ _27248;
  wire _27250 = _20941 ^ _12425;
  wire _27251 = _26847 ^ _27250;
  wire _27252 = uncoded_block[49] ^ uncoded_block[59];
  wire _27253 = _7359 ^ _27252;
  wire _27254 = _13553 ^ _10806;
  wire _27255 = _27253 ^ _27254;
  wire _27256 = _27251 ^ _27255;
  wire _27257 = _27249 ^ _27256;
  wire _27258 = _4020 ^ _901;
  wire _27259 = _898 ^ _27258;
  wire _27260 = _17077 ^ _6755;
  wire _27261 = _21885 ^ _27260;
  wire _27262 = _27259 ^ _27261;
  wire _27263 = _8566 ^ _6115;
  wire _27264 = _1719 ^ _15097;
  wire _27265 = _27263 ^ _27264;
  wire _27266 = _15101 ^ _14595;
  wire _27267 = _2491 ^ _6126;
  wire _27268 = _27266 ^ _27267;
  wire _27269 = _27265 ^ _27268;
  wire _27270 = _27262 ^ _27269;
  wire _27271 = _27257 ^ _27270;
  wire _27272 = _23269 ^ _7386;
  wire _27273 = _8576 ^ _27272;
  wire _27274 = uncoded_block[133] ^ uncoded_block[137];
  wire _27275 = uncoded_block[139] ^ uncoded_block[144];
  wire _27276 = _27274 ^ _27275;
  wire _27277 = _12458 ^ _27276;
  wire _27278 = _27273 ^ _27277;
  wire _27279 = _8000 ^ _9186;
  wire _27280 = _4049 ^ _4053;
  wire _27281 = _27279 ^ _27280;
  wire _27282 = _81 ^ _15126;
  wire _27283 = _18578 ^ _27282;
  wire _27284 = _27281 ^ _27283;
  wire _27285 = _27278 ^ _27284;
  wire _27286 = _2525 ^ _17106;
  wire _27287 = _18111 ^ _18113;
  wire _27288 = _27286 ^ _27287;
  wire _27289 = uncoded_block[193] ^ uncoded_block[197];
  wire _27290 = _27289 ^ _9745;
  wire _27291 = _14099 ^ _1764;
  wire _27292 = _27290 ^ _27291;
  wire _27293 = _27288 ^ _27292;
  wire _27294 = _8600 ^ _955;
  wire _27295 = uncoded_block[214] ^ uncoded_block[216];
  wire _27296 = _19549 ^ _27295;
  wire _27297 = _27294 ^ _27296;
  wire _27298 = _960 ^ _5492;
  wire _27299 = _109 ^ _1774;
  wire _27300 = _27298 ^ _27299;
  wire _27301 = _27297 ^ _27300;
  wire _27302 = _27293 ^ _27301;
  wire _27303 = _27285 ^ _27302;
  wire _27304 = _27271 ^ _27303;
  wire _27305 = uncoded_block[231] ^ uncoded_block[237];
  wire _27306 = _27305 ^ _10860;
  wire _27307 = _27306 ^ _6827;
  wire _27308 = _11420 ^ _26442;
  wire _27309 = _27307 ^ _27308;
  wire _27310 = _21007 ^ _4813;
  wire _27311 = _10303 ^ _1796;
  wire _27312 = _27310 ^ _27311;
  wire _27313 = _4819 ^ _8636;
  wire _27314 = _23757 ^ _27313;
  wire _27315 = _27312 ^ _27314;
  wire _27316 = _27309 ^ _27315;
  wire _27317 = _142 ^ _4114;
  wire _27318 = _27317 ^ _20042;
  wire _27319 = _20539 ^ _1008;
  wire _27320 = uncoded_block[323] ^ uncoded_block[329];
  wire _27321 = _3346 ^ _27320;
  wire _27322 = _27319 ^ _27321;
  wire _27323 = _27318 ^ _27322;
  wire _27324 = _4126 ^ _1018;
  wire _27325 = _27324 ^ _13088;
  wire _27326 = uncoded_block[352] ^ uncoded_block[356];
  wire _27327 = _1023 ^ _27326;
  wire _27328 = uncoded_block[362] ^ uncoded_block[366];
  wire _27329 = _27328 ^ _1835;
  wire _27330 = _27327 ^ _27329;
  wire _27331 = _27325 ^ _27330;
  wire _27332 = _27323 ^ _27331;
  wire _27333 = _27316 ^ _27332;
  wire _27334 = uncoded_block[373] ^ uncoded_block[377];
  wire _27335 = _27334 ^ _6876;
  wire _27336 = _9796 ^ _27335;
  wire _27337 = _5552 ^ _3381;
  wire _27338 = _14678 ^ _25141;
  wire _27339 = _27337 ^ _27338;
  wire _27340 = _27336 ^ _27339;
  wire _27341 = uncoded_block[407] ^ uncoded_block[411];
  wire _27342 = _27341 ^ _2630;
  wire _27343 = _27342 ^ _9268;
  wire _27344 = uncoded_block[422] ^ uncoded_block[426];
  wire _27345 = _27344 ^ _9816;
  wire _27346 = _1063 ^ _9271;
  wire _27347 = _27345 ^ _27346;
  wire _27348 = _27343 ^ _27347;
  wire _27349 = _27340 ^ _27348;
  wire _27350 = uncoded_block[435] ^ uncoded_block[439];
  wire _27351 = _27350 ^ _206;
  wire _27352 = _4177 ^ _14173;
  wire _27353 = _27351 ^ _27352;
  wire _27354 = uncoded_block[459] ^ uncoded_block[463];
  wire _27355 = _27354 ^ _21523;
  wire _27356 = _221 ^ _5590;
  wire _27357 = _27355 ^ _27356;
  wire _27358 = _27353 ^ _27357;
  wire _27359 = _1090 ^ _17198;
  wire _27360 = _17195 ^ _27359;
  wire _27361 = uncoded_block[503] ^ uncoded_block[506];
  wire _27362 = _27361 ^ _5611;
  wire _27363 = _6280 ^ _27362;
  wire _27364 = _27360 ^ _27363;
  wire _27365 = _27358 ^ _27364;
  wire _27366 = _27349 ^ _27365;
  wire _27367 = _27333 ^ _27366;
  wire _27368 = _27304 ^ _27367;
  wire _27369 = uncoded_block[509] ^ uncoded_block[512];
  wire _27370 = _27369 ^ _10945;
  wire _27371 = _20598 ^ _237;
  wire _27372 = _27370 ^ _27371;
  wire _27373 = uncoded_block[527] ^ uncoded_block[532];
  wire _27374 = _4921 ^ _27373;
  wire _27375 = uncoded_block[534] ^ uncoded_block[537];
  wire _27376 = uncoded_block[539] ^ uncoded_block[544];
  wire _27377 = _27375 ^ _27376;
  wire _27378 = _27374 ^ _27377;
  wire _27379 = _27372 ^ _27378;
  wire _27380 = _1912 ^ _5630;
  wire _27381 = _1123 ^ _24284;
  wire _27382 = _27380 ^ _27381;
  wire _27383 = _24289 ^ _270;
  wire _27384 = _1131 ^ _27383;
  wire _27385 = _27382 ^ _27384;
  wire _27386 = _27379 ^ _27385;
  wire _27387 = _20618 ^ _15247;
  wire _27388 = _27387 ^ _2708;
  wire _27389 = _9870 ^ _12609;
  wire _27390 = uncoded_block[618] ^ uncoded_block[623];
  wire _27391 = _5652 ^ _27390;
  wire _27392 = _27389 ^ _27391;
  wire _27393 = _27388 ^ _27392;
  wire _27394 = _1154 ^ _12620;
  wire _27395 = uncoded_block[633] ^ uncoded_block[640];
  wire _27396 = _27395 ^ _294;
  wire _27397 = _27394 ^ _27396;
  wire _27398 = uncoded_block[645] ^ uncoded_block[650];
  wire _27399 = _27398 ^ _302;
  wire _27400 = _3508 ^ _2739;
  wire _27401 = _27399 ^ _27400;
  wire _27402 = _27397 ^ _27401;
  wire _27403 = _27393 ^ _27402;
  wire _27404 = _27386 ^ _27403;
  wire _27405 = _4978 ^ _309;
  wire _27406 = _1174 ^ _17745;
  wire _27407 = _27405 ^ _27406;
  wire _27408 = uncoded_block[677] ^ uncoded_block[681];
  wire _27409 = _10434 ^ _27408;
  wire _27410 = _2750 ^ _325;
  wire _27411 = _27409 ^ _27410;
  wire _27412 = _27407 ^ _27411;
  wire _27413 = uncoded_block[695] ^ uncoded_block[701];
  wire _27414 = _6985 ^ _27413;
  wire _27415 = _24320 ^ _11004;
  wire _27416 = _27414 ^ _27415;
  wire _27417 = _6999 ^ _8200;
  wire _27418 = _9370 ^ _27417;
  wire _27419 = _27416 ^ _27418;
  wire _27420 = _27412 ^ _27419;
  wire _27421 = _8201 ^ _1995;
  wire _27422 = _27421 ^ _21135;
  wire _27423 = _11576 ^ _10464;
  wire _27424 = _1210 ^ _2003;
  wire _27425 = _27423 ^ _27424;
  wire _27426 = _27422 ^ _27425;
  wire _27427 = uncoded_block[763] ^ uncoded_block[767];
  wire _27428 = _27427 ^ _9917;
  wire _27429 = _14269 ^ _27428;
  wire _27430 = _15799 ^ _6386;
  wire _27431 = _16786 ^ _19709;
  wire _27432 = _27430 ^ _27431;
  wire _27433 = _27429 ^ _27432;
  wire _27434 = _27426 ^ _27433;
  wire _27435 = _27420 ^ _27434;
  wire _27436 = _27404 ^ _27435;
  wire _27437 = _5723 ^ _8223;
  wire _27438 = _8224 ^ _8793;
  wire _27439 = _27437 ^ _27438;
  wire _27440 = _5041 ^ _10483;
  wire _27441 = uncoded_block[815] ^ uncoded_block[824];
  wire _27442 = _10485 ^ _27441;
  wire _27443 = _27440 ^ _27442;
  wire _27444 = _27439 ^ _27443;
  wire _27445 = _23896 ^ _4331;
  wire _27446 = _4336 ^ _9938;
  wire _27447 = _27445 ^ _27446;
  wire _27448 = _13238 ^ _26164;
  wire _27449 = _5059 ^ _27448;
  wire _27450 = _27447 ^ _27449;
  wire _27451 = _27444 ^ _27450;
  wire _27452 = uncoded_block[865] ^ uncoded_block[868];
  wire _27453 = _27452 ^ _4346;
  wire _27454 = _23459 ^ _27453;
  wire _27455 = _11620 ^ _2835;
  wire _27456 = _5079 ^ _14821;
  wire _27457 = _27455 ^ _27456;
  wire _27458 = _27454 ^ _27457;
  wire _27459 = _7660 ^ _4354;
  wire _27460 = _18307 ^ _428;
  wire _27461 = _27459 ^ _27460;
  wire _27462 = _2843 ^ _1280;
  wire _27463 = uncoded_block[911] ^ uncoded_block[915];
  wire _27464 = _1284 ^ _27463;
  wire _27465 = _27462 ^ _27464;
  wire _27466 = _27461 ^ _27465;
  wire _27467 = _27458 ^ _27466;
  wire _27468 = _27451 ^ _27467;
  wire _27469 = _2852 ^ _18775;
  wire _27470 = _11634 ^ _4371;
  wire _27471 = _27469 ^ _27470;
  wire _27472 = _5101 ^ _7080;
  wire _27473 = _453 ^ _13263;
  wire _27474 = _27472 ^ _27473;
  wire _27475 = _27471 ^ _27474;
  wire _27476 = uncoded_block[946] ^ uncoded_block[951];
  wire _27477 = _27476 ^ _5779;
  wire _27478 = uncoded_block[957] ^ uncoded_block[961];
  wire _27479 = _2869 ^ _27478;
  wire _27480 = _27477 ^ _27479;
  wire _27481 = _19268 ^ _11092;
  wire _27482 = _7089 ^ _27481;
  wire _27483 = _27480 ^ _27482;
  wire _27484 = _27475 ^ _27483;
  wire _27485 = _476 ^ _12186;
  wire _27486 = _15369 ^ _1323;
  wire _27487 = _27485 ^ _27486;
  wire _27488 = _6453 ^ _11101;
  wire _27489 = _27488 ^ _18335;
  wire _27490 = _27487 ^ _27489;
  wire _27491 = _20730 ^ _486;
  wire _27492 = _487 ^ _492;
  wire _27493 = _27491 ^ _27492;
  wire _27494 = uncoded_block[1023] ^ uncoded_block[1026];
  wire _27495 = _7108 ^ _27494;
  wire _27496 = uncoded_block[1027] ^ uncoded_block[1032];
  wire _27497 = _27496 ^ _501;
  wire _27498 = _27495 ^ _27497;
  wire _27499 = _27493 ^ _27498;
  wire _27500 = _27490 ^ _27499;
  wire _27501 = _27484 ^ _27500;
  wire _27502 = _27468 ^ _27501;
  wire _27503 = _27436 ^ _27502;
  wire _27504 = _27368 ^ _27503;
  wire _27505 = uncoded_block[1036] ^ uncoded_block[1040];
  wire _27506 = _27505 ^ _512;
  wire _27507 = uncoded_block[1046] ^ uncoded_block[1056];
  wire _27508 = _27507 ^ _7117;
  wire _27509 = _27506 ^ _27508;
  wire _27510 = _13849 ^ _8889;
  wire _27511 = _12217 ^ _2146;
  wire _27512 = _27510 ^ _27511;
  wire _27513 = _27509 ^ _27512;
  wire _27514 = _8895 ^ _11126;
  wire _27515 = uncoded_block[1083] ^ uncoded_block[1090];
  wire _27516 = _27515 ^ _22610;
  wire _27517 = _27514 ^ _27516;
  wire _27518 = _3698 ^ _12224;
  wire _27519 = uncoded_block[1103] ^ uncoded_block[1106];
  wire _27520 = _27519 ^ _7132;
  wire _27521 = _27518 ^ _27520;
  wire _27522 = _27517 ^ _27521;
  wire _27523 = _27513 ^ _27522;
  wire _27524 = _3714 ^ _2942;
  wire _27525 = _23520 ^ _27524;
  wire _27526 = uncoded_block[1131] ^ uncoded_block[1135];
  wire _27527 = _23523 ^ _27526;
  wire _27528 = uncoded_block[1138] ^ uncoded_block[1142];
  wire _27529 = _27528 ^ _2180;
  wire _27530 = _27527 ^ _27529;
  wire _27531 = _27525 ^ _27530;
  wire _27532 = uncoded_block[1149] ^ uncoded_block[1151];
  wire _27533 = _27532 ^ _4468;
  wire _27534 = uncoded_block[1156] ^ uncoded_block[1162];
  wire _27535 = _27534 ^ _15907;
  wire _27536 = _27533 ^ _27535;
  wire _27537 = uncoded_block[1169] ^ uncoded_block[1172];
  wire _27538 = _27537 ^ _3739;
  wire _27539 = uncoded_block[1178] ^ uncoded_block[1180];
  wire _27540 = _17396 ^ _27539;
  wire _27541 = _27538 ^ _27540;
  wire _27542 = _27536 ^ _27541;
  wire _27543 = _27531 ^ _27542;
  wire _27544 = _27523 ^ _27543;
  wire _27545 = uncoded_block[1181] ^ uncoded_block[1186];
  wire _27546 = _27545 ^ _2201;
  wire _27547 = _3749 ^ _24910;
  wire _27548 = _27546 ^ _27547;
  wire _27549 = uncoded_block[1198] ^ uncoded_block[1201];
  wire _27550 = _22179 ^ _27549;
  wire _27551 = _6529 ^ _2979;
  wire _27552 = _27550 ^ _27551;
  wire _27553 = _27548 ^ _27552;
  wire _27554 = _18395 ^ _2219;
  wire _27555 = _606 ^ _4502;
  wire _27556 = _27554 ^ _27555;
  wire _27557 = _26702 ^ _14411;
  wire _27558 = _27556 ^ _27557;
  wire _27559 = _27553 ^ _27558;
  wire _27560 = _5219 ^ _2230;
  wire _27561 = uncoded_block[1243] ^ uncoded_block[1251];
  wire _27562 = _10627 ^ _27561;
  wire _27563 = _27560 ^ _27562;
  wire _27564 = uncoded_block[1255] ^ uncoded_block[1264];
  wire _27565 = _27564 ^ _24927;
  wire _27566 = _27565 ^ _10637;
  wire _27567 = _27563 ^ _27566;
  wire _27568 = _6557 ^ _5243;
  wire _27569 = _24482 ^ _25377;
  wire _27570 = _27568 ^ _27569;
  wire _27571 = _3805 ^ _648;
  wire _27572 = _26275 ^ _27571;
  wire _27573 = _27570 ^ _27572;
  wire _27574 = _27567 ^ _27573;
  wire _27575 = _27559 ^ _27574;
  wire _27576 = _27544 ^ _27575;
  wire _27577 = _6572 ^ _14430;
  wire _27578 = _3811 ^ _3028;
  wire _27579 = _27577 ^ _27578;
  wire _27580 = _5931 ^ _3034;
  wire _27581 = _658 ^ _27580;
  wire _27582 = _27579 ^ _27581;
  wire _27583 = uncoded_block[1347] ^ uncoded_block[1357];
  wire _27584 = _27583 ^ _7821;
  wire _27585 = _9004 ^ _27584;
  wire _27586 = _22224 ^ _22229;
  wire _27587 = _1505 ^ _27586;
  wire _27588 = _27585 ^ _27587;
  wire _27589 = _27582 ^ _27588;
  wire _27590 = uncoded_block[1384] ^ uncoded_block[1388];
  wire _27591 = _687 ^ _27590;
  wire _27592 = _4569 ^ _7834;
  wire _27593 = _27591 ^ _27592;
  wire _27594 = _9585 ^ _5961;
  wire _27595 = _20838 ^ _27594;
  wire _27596 = _27593 ^ _27595;
  wire _27597 = _17461 ^ _13422;
  wire _27598 = _705 ^ _16463;
  wire _27599 = _27597 ^ _27598;
  wire _27600 = _15494 ^ _15498;
  wire _27601 = _10690 ^ _2318;
  wire _27602 = _27600 ^ _27601;
  wire _27603 = _27599 ^ _27602;
  wire _27604 = _27596 ^ _27603;
  wire _27605 = _27589 ^ _27604;
  wire _27606 = _4590 ^ _5970;
  wire _27607 = _27606 ^ _13436;
  wire _27608 = _20852 ^ _13437;
  wire _27609 = _3870 ^ _8455;
  wire _27610 = _27608 ^ _27609;
  wire _27611 = _27607 ^ _27610;
  wire _27612 = _1548 ^ _25871;
  wire _27613 = _27612 ^ _17978;
  wire _27614 = _3884 ^ _21799;
  wire _27615 = _7251 ^ _4610;
  wire _27616 = _27614 ^ _27615;
  wire _27617 = _27613 ^ _27616;
  wire _27618 = _27611 ^ _27617;
  wire _27619 = _7257 ^ _14486;
  wire _27620 = _7262 ^ _11266;
  wire _27621 = uncoded_block[1517] ^ uncoded_block[1519];
  wire _27622 = _9621 ^ _27621;
  wire _27623 = _27620 ^ _27622;
  wire _27624 = _27619 ^ _27623;
  wire _27625 = _2359 ^ _6002;
  wire _27626 = uncoded_block[1539] ^ uncoded_block[1544];
  wire _27627 = _15009 ^ _27626;
  wire _27628 = _27625 ^ _27627;
  wire _27629 = _1593 ^ _13472;
  wire _27630 = _7885 ^ _22731;
  wire _27631 = _27629 ^ _27630;
  wire _27632 = _27628 ^ _27631;
  wire _27633 = _27624 ^ _27632;
  wire _27634 = _27618 ^ _27633;
  wire _27635 = _27605 ^ _27634;
  wire _27636 = _27576 ^ _27635;
  wire _27637 = _6016 ^ _23640;
  wire _27638 = _5363 ^ _6028;
  wire _27639 = _27637 ^ _27638;
  wire _27640 = _784 ^ _1612;
  wire _27641 = uncoded_block[1590] ^ uncoded_block[1594];
  wire _27642 = _2386 ^ _27641;
  wire _27643 = _27640 ^ _27642;
  wire _27644 = _27639 ^ _27643;
  wire _27645 = _11295 ^ _6039;
  wire _27646 = uncoded_block[1604] ^ uncoded_block[1609];
  wire _27647 = _27646 ^ _1633;
  wire _27648 = _27645 ^ _27647;
  wire _27649 = uncoded_block[1621] ^ uncoded_block[1628];
  wire _27650 = _27649 ^ _4667;
  wire _27651 = uncoded_block[1641] ^ uncoded_block[1643];
  wire _27652 = _5392 ^ _27651;
  wire _27653 = _27650 ^ _27652;
  wire _27654 = _27648 ^ _27653;
  wire _27655 = _27644 ^ _27654;
  wire _27656 = _17529 ^ _6696;
  wire _27657 = _18517 ^ _27656;
  wire _27658 = _4680 ^ _3179;
  wire _27659 = _7322 ^ _830;
  wire _27660 = _27658 ^ _27659;
  wire _27661 = _27657 ^ _27660;
  wire _27662 = _1662 ^ _10766;
  wire _27663 = _6061 ^ _24130;
  wire _27664 = _27662 ^ _27663;
  wire _27665 = _837 ^ _839;
  wire _27666 = _27665 ^ _22771;
  wire _27667 = _27664 ^ _27666;
  wire _27668 = _27661 ^ _27667;
  wire _27669 = _27655 ^ _27668;
  wire _27670 = _25037 ^ _20920;
  wire _27671 = uncoded_block[1708] ^ uncoded_block[1710];
  wire _27672 = _27671 ^ _7337;
  wire _27673 = _27670 ^ _27672;
  wire _27674 = _7944 ^ _3988;
  wire _27675 = _27674 ^ uncoded_block[1721];
  wire _27676 = _27673 ^ _27675;
  wire _27677 = _27669 ^ _27676;
  wire _27678 = _27636 ^ _27677;
  wire _27679 = _27504 ^ _27678;
  wire _27680 = _26846 ^ _25943;
  wire _27681 = _25945 ^ _3234;
  wire _27682 = _4014 ^ _7364;
  wire _27683 = _27682 ^ _25951;
  wire _27684 = _27681 ^ _27683;
  wire _27685 = _27680 ^ _27684;
  wire _27686 = _6754 ^ _6757;
  wire _27687 = _25956 ^ _27686;
  wire _27688 = _7375 ^ _49;
  wire _27689 = _27688 ^ _2492;
  wire _27690 = _27687 ^ _27689;
  wire _27691 = _54 ^ _2498;
  wire _27692 = _10817 ^ _27691;
  wire _27693 = _7386 ^ _923;
  wire _27694 = _1735 ^ _4043;
  wire _27695 = _27693 ^ _27694;
  wire _27696 = _27692 ^ _27695;
  wire _27697 = _27690 ^ _27696;
  wire _27698 = _27685 ^ _27697;
  wire _27699 = _7392 ^ _21901;
  wire _27700 = _27699 ^ _20489;
  wire _27701 = uncoded_block[157] ^ uncoded_block[167];
  wire _27702 = _27701 ^ _1752;
  wire _27703 = _14614 ^ _11933;
  wire _27704 = _27702 ^ _27703;
  wire _27705 = _27700 ^ _27704;
  wire _27706 = _7408 ^ _945;
  wire _27707 = _27706 ^ _15636;
  wire _27708 = _27707 ^ _26880;
  wire _27709 = _27705 ^ _27708;
  wire _27710 = _4791 ^ _967;
  wire _27711 = _26883 ^ _27710;
  wire _27712 = _10289 ^ _21465;
  wire _27713 = _27712 ^ _26888;
  wire _27714 = _27711 ^ _27713;
  wire _27715 = _20523 ^ _14642;
  wire _27716 = uncoded_block[278] ^ uncoded_block[282];
  wire _27717 = _14124 ^ _27716;
  wire _27718 = _27715 ^ _27717;
  wire _27719 = _26893 ^ _27718;
  wire _27720 = _27714 ^ _27719;
  wire _27721 = _27709 ^ _27720;
  wire _27722 = _27698 ^ _27721;
  wire _27723 = _26009 ^ _26011;
  wire _27724 = _26013 ^ _26017;
  wire _27725 = _27723 ^ _27724;
  wire _27726 = _3340 ^ _13624;
  wire _27727 = _1818 ^ _4123;
  wire _27728 = _27726 ^ _27727;
  wire _27729 = _9782 ^ _1017;
  wire _27730 = _7463 ^ _1021;
  wire _27731 = _27729 ^ _27730;
  wire _27732 = _27728 ^ _27731;
  wire _27733 = _27725 ^ _27732;
  wire _27734 = _7465 ^ _3359;
  wire _27735 = _14662 ^ _2601;
  wire _27736 = _27734 ^ _27735;
  wire _27737 = _2602 ^ _2606;
  wire _27738 = _17163 ^ _17165;
  wire _27739 = _27737 ^ _27738;
  wire _27740 = _27736 ^ _27739;
  wire _27741 = _4140 ^ _10898;
  wire _27742 = _13101 ^ _11999;
  wire _27743 = _27741 ^ _27742;
  wire _27744 = _27743 ^ _26044;
  wire _27745 = _27740 ^ _27744;
  wire _27746 = _27733 ^ _27745;
  wire _27747 = _4867 ^ _191;
  wire _27748 = _6885 ^ _27747;
  wire _27749 = _1055 ^ _193;
  wire _27750 = _27749 ^ _14161;
  wire _27751 = _27748 ^ _27750;
  wire _27752 = uncoded_block[425] ^ uncoded_block[429];
  wire _27753 = _8671 ^ _27752;
  wire _27754 = _6254 ^ _16187;
  wire _27755 = _27753 ^ _27754;
  wire _27756 = uncoded_block[447] ^ uncoded_block[451];
  wire _27757 = _9275 ^ _27756;
  wire _27758 = _207 ^ _27757;
  wire _27759 = _27755 ^ _27758;
  wire _27760 = _27751 ^ _27759;
  wire _27761 = _2645 ^ _2650;
  wire _27762 = _27761 ^ _18185;
  wire _27763 = _13662 ^ _1874;
  wire _27764 = _27763 ^ _26063;
  wire _27765 = _27762 ^ _27764;
  wire _27766 = uncoded_block[481] ^ uncoded_block[487];
  wire _27767 = _27766 ^ _17198;
  wire _27768 = _26065 ^ _27767;
  wire _27769 = uncoded_block[494] ^ uncoded_block[496];
  wire _27770 = _27769 ^ _5604;
  wire _27771 = _228 ^ _19135;
  wire _27772 = _27770 ^ _27771;
  wire _27773 = _27768 ^ _27772;
  wire _27774 = _27765 ^ _27773;
  wire _27775 = _27760 ^ _27774;
  wire _27776 = _27746 ^ _27775;
  wire _27777 = _27722 ^ _27776;
  wire _27778 = _17203 ^ _4909;
  wire _27779 = _1900 ^ _1905;
  wire _27780 = _1899 ^ _27779;
  wire _27781 = _27778 ^ _27780;
  wire _27782 = uncoded_block[540] ^ uncoded_block[546];
  wire _27783 = _14197 ^ _27782;
  wire _27784 = _12592 ^ _3459;
  wire _27785 = _27783 ^ _27784;
  wire _27786 = _1925 ^ _1927;
  wire _27787 = _8138 ^ _27786;
  wire _27788 = _27785 ^ _27787;
  wire _27789 = _27781 ^ _27788;
  wire _27790 = _17221 ^ _26094;
  wire _27791 = _27790 ^ _26975;
  wire _27792 = _27791 ^ _26979;
  wire _27793 = _3486 ^ _1941;
  wire _27794 = _6323 ^ _15758;
  wire _27795 = _27793 ^ _27794;
  wire _27796 = _13713 ^ _20125;
  wire _27797 = uncoded_block[622] ^ uncoded_block[628];
  wire _27798 = _27797 ^ _1953;
  wire _27799 = _27796 ^ _27798;
  wire _27800 = _27795 ^ _27799;
  wire _27801 = _27792 ^ _27800;
  wire _27802 = _27789 ^ _27801;
  wire _27803 = _5661 ^ _1161;
  wire _27804 = _27803 ^ _12077;
  wire _27805 = _1960 ^ _19181;
  wire _27806 = _26547 ^ _27805;
  wire _27807 = _27804 ^ _27806;
  wire _27808 = _308 ^ _311;
  wire _27809 = _11548 ^ _27808;
  wire _27810 = _16752 ^ _10434;
  wire _27811 = _27810 ^ _26122;
  wire _27812 = _27809 ^ _27811;
  wire _27813 = _27807 ^ _27812;
  wire _27814 = _22491 ^ _26124;
  wire _27815 = _26125 ^ _26563;
  wire _27816 = _27814 ^ _27815;
  wire _27817 = _16766 ^ _19693;
  wire _27818 = uncoded_block[729] ^ uncoded_block[739];
  wire _27819 = _6999 ^ _27818;
  wire _27820 = _1207 ^ _5702;
  wire _27821 = _27819 ^ _27820;
  wire _27822 = _27817 ^ _27821;
  wire _27823 = _27816 ^ _27822;
  wire _27824 = _27813 ^ _27823;
  wire _27825 = _27802 ^ _27824;
  wire _27826 = _356 ^ _4295;
  wire _27827 = uncoded_block[755] ^ uncoded_block[759];
  wire _27828 = _27827 ^ _9914;
  wire _27829 = _27826 ^ _27828;
  wire _27830 = _1217 ^ _1221;
  wire _27831 = _3562 ^ _368;
  wire _27832 = _27830 ^ _27831;
  wire _27833 = _27829 ^ _27832;
  wire _27834 = _3568 ^ _371;
  wire _27835 = _5032 ^ _1225;
  wire _27836 = _27834 ^ _27835;
  wire _27837 = _11024 ^ _7628;
  wire _27838 = _385 ^ _1235;
  wire _27839 = _27837 ^ _27838;
  wire _27840 = _27836 ^ _27839;
  wire _27841 = _27833 ^ _27840;
  wire _27842 = _14287 ^ _2806;
  wire _27843 = uncoded_block[820] ^ uncoded_block[822];
  wire _27844 = _22525 ^ _27843;
  wire _27845 = _27842 ^ _27844;
  wire _27846 = uncoded_block[830] ^ uncoded_block[835];
  wire _27847 = _23450 ^ _27846;
  wire _27848 = _12138 ^ _5057;
  wire _27849 = _27847 ^ _27848;
  wire _27850 = _27845 ^ _27849;
  wire _27851 = _14812 ^ _11610;
  wire _27852 = _12146 ^ _15330;
  wire _27853 = _27851 ^ _27852;
  wire _27854 = _26166 ^ _26172;
  wire _27855 = _27853 ^ _27854;
  wire _27856 = _27850 ^ _27855;
  wire _27857 = _27841 ^ _27856;
  wire _27858 = _13791 ^ _25719;
  wire _27859 = _27858 ^ _2837;
  wire _27860 = _423 ^ _27046;
  wire _27861 = _5083 ^ _27048;
  wire _27862 = _27860 ^ _27861;
  wire _27863 = _27859 ^ _27862;
  wire _27864 = _26180 ^ _26182;
  wire _27865 = _26184 ^ _27055;
  wire _27866 = _27864 ^ _27865;
  wire _27867 = _27863 ^ _27866;
  wire _27868 = _27056 ^ _27060;
  wire _27869 = _27061 ^ _26194;
  wire _27870 = _27868 ^ _27869;
  wire _27871 = _27870 ^ _26202;
  wire _27872 = _27867 ^ _27871;
  wire _27873 = _27857 ^ _27872;
  wire _27874 = _27825 ^ _27873;
  wire _27875 = _27777 ^ _27874;
  wire _27876 = _13277 ^ _5798;
  wire _27877 = _2114 ^ _27077;
  wire _27878 = _27876 ^ _27877;
  wire _27879 = _8296 ^ _7703;
  wire _27880 = _1334 ^ _27081;
  wire _27881 = _27879 ^ _27880;
  wire _27882 = _27878 ^ _27881;
  wire _27883 = _2907 ^ _27085;
  wire _27884 = _27883 ^ _14866;
  wire _27885 = _1363 ^ _2921;
  wire _27886 = _26218 ^ _27885;
  wire _27887 = _27884 ^ _27886;
  wire _27888 = _27882 ^ _27887;
  wire _27889 = _8895 ^ _26225;
  wire _27890 = _27091 ^ _27889;
  wire _27891 = _19790 ^ _13320;
  wire _27892 = _27890 ^ _27891;
  wire _27893 = _27099 ^ _27102;
  wire _27894 = _4462 ^ _5859;
  wire _27895 = _26679 ^ _3727;
  wire _27896 = _27894 ^ _27895;
  wire _27897 = _27893 ^ _27896;
  wire _27898 = _27892 ^ _27897;
  wire _27899 = _27888 ^ _27898;
  wire _27900 = _5190 ^ _26244;
  wire _27901 = _27900 ^ _25340;
  wire _27902 = uncoded_block[1173] ^ uncoded_block[1176];
  wire _27903 = _27902 ^ _4481;
  wire _27904 = _27113 ^ _27116;
  wire _27905 = _27903 ^ _27904;
  wire _27906 = _27901 ^ _27905;
  wire _27907 = _3747 ^ _3749;
  wire _27908 = _1421 ^ _17400;
  wire _27909 = _27907 ^ _27908;
  wire _27910 = _24456 ^ _23544;
  wire _27911 = uncoded_block[1211] ^ uncoded_block[1215];
  wire _27912 = uncoded_block[1217] ^ uncoded_block[1224];
  wire _27913 = _27911 ^ _27912;
  wire _27914 = _27910 ^ _27913;
  wire _27915 = _27909 ^ _27914;
  wire _27916 = _27906 ^ _27915;
  wire _27917 = _27125 ^ _27130;
  wire _27918 = _27131 ^ _26262;
  wire _27919 = _27917 ^ _27918;
  wire _27920 = _26263 ^ _13371;
  wire _27921 = _27134 ^ _27136;
  wire _27922 = _27920 ^ _27921;
  wire _27923 = _27919 ^ _27922;
  wire _27924 = _27916 ^ _27923;
  wire _27925 = _27899 ^ _27924;
  wire _27926 = _18866 ^ _3800;
  wire _27927 = _27926 ^ _27143;
  wire _27928 = _27144 ^ _27146;
  wire _27929 = _27927 ^ _27928;
  wire _27930 = _4544 ^ _27149;
  wire _27931 = _19849 ^ _27152;
  wire _27932 = _27930 ^ _27931;
  wire _27933 = _27929 ^ _27932;
  wire _27934 = _27153 ^ _27158;
  wire _27935 = _27934 ^ _26290;
  wire _27936 = _27935 ^ _26297;
  wire _27937 = _27933 ^ _27936;
  wire _27938 = _4580 ^ _13422;
  wire _27939 = _2306 ^ _7842;
  wire _27940 = _27938 ^ _27939;
  wire _27941 = _1527 ^ _10684;
  wire _27942 = _1531 ^ _16962;
  wire _27943 = _27941 ^ _27942;
  wire _27944 = _27940 ^ _27943;
  wire _27945 = _8455 ^ _22254;
  wire _27946 = _26312 ^ _27945;
  wire _27947 = _26311 ^ _27946;
  wire _27948 = _27944 ^ _27947;
  wire _27949 = _27182 ^ _11807;
  wire _27950 = _27949 ^ _27615;
  wire _27951 = _12896 ^ _743;
  wire _27952 = _6634 ^ _7258;
  wire _27953 = _27951 ^ _27952;
  wire _27954 = _27950 ^ _27953;
  wire _27955 = _26782 ^ _9054;
  wire _27956 = _1582 ^ _9631;
  wire _27957 = _756 ^ _27956;
  wire _27958 = _27955 ^ _27957;
  wire _27959 = _27954 ^ _27958;
  wire _27960 = _27948 ^ _27959;
  wire _27961 = _27937 ^ _27960;
  wire _27962 = _27925 ^ _27961;
  wire _27963 = _5347 ^ _6651;
  wire _27964 = _27963 ^ _16500;
  wire _27965 = _13473 ^ _16997;
  wire _27966 = _27964 ^ _27965;
  wire _27967 = _2386 ^ _12934;
  wire _27968 = uncoded_block[1600] ^ uncoded_block[1605];
  wire _27969 = _13486 ^ _27968;
  wire _27970 = _27967 ^ _27969;
  wire _27971 = _27205 ^ _27970;
  wire _27972 = _27966 ^ _27971;
  wire _27973 = _2396 ^ _3937;
  wire _27974 = _1632 ^ _16032;
  wire _27975 = _27973 ^ _27974;
  wire _27976 = _27975 ^ _27218;
  wire _27977 = uncoded_block[1652] ^ uncoded_block[1657];
  wire _27978 = _1649 ^ _27977;
  wire _27979 = _1653 ^ _12960;
  wire _27980 = _27978 ^ _27979;
  wire _27981 = _26357 ^ _17037;
  wire _27982 = _27980 ^ _27981;
  wire _27983 = _27976 ^ _27982;
  wire _27984 = _27972 ^ _27983;
  wire _27985 = _13519 ^ _26365;
  wire _27986 = _26360 ^ _27985;
  wire _27987 = _26367 ^ _24138;
  wire _27988 = _27986 ^ _27987;
  wire _27989 = _26370 ^ _26373;
  wire _27990 = _27989 ^ uncoded_block[1722];
  wire _27991 = _27988 ^ _27990;
  wire _27992 = _27984 ^ _27991;
  wire _27993 = _27962 ^ _27992;
  wire _27994 = _27875 ^ _27993;
  wire _27995 = _3209 ^ _24147;
  wire _27996 = _6083 ^ _15075;
  wire _27997 = _27995 ^ _27996;
  wire _27998 = uncoded_block[20] ^ uncoded_block[24];
  wire _27999 = _5423 ^ _27998;
  wire _28000 = uncoded_block[26] ^ uncoded_block[32];
  wire _28001 = _28000 ^ _18548;
  wire _28002 = _27999 ^ _28001;
  wire _28003 = _27997 ^ _28002;
  wire _28004 = _18 ^ _15591;
  wire _28005 = _8554 ^ _1699;
  wire _28006 = _28004 ^ _28005;
  wire _28007 = _8556 ^ _7364;
  wire _28008 = uncoded_block[66] ^ uncoded_block[70];
  wire _28009 = _10806 ^ _28008;
  wire _28010 = _28007 ^ _28009;
  wire _28011 = _28006 ^ _28010;
  wire _28012 = _28003 ^ _28011;
  wire _28013 = _22805 ^ _25957;
  wire _28014 = _19017 ^ _28013;
  wire _28015 = _12442 ^ _46;
  wire _28016 = _3249 ^ _15101;
  wire _28017 = _28015 ^ _28016;
  wire _28018 = _28014 ^ _28017;
  wire _28019 = _6120 ^ _20957;
  wire _28020 = _28019 ^ _916;
  wire _28021 = uncoded_block[119] ^ uncoded_block[125];
  wire _28022 = uncoded_block[127] ^ uncoded_block[132];
  wire _28023 = _28021 ^ _28022;
  wire _28024 = _28023 ^ _11917;
  wire _28025 = _28020 ^ _28024;
  wire _28026 = _28018 ^ _28025;
  wire _28027 = _28012 ^ _28026;
  wire _28028 = _64 ^ _4761;
  wire _28029 = _70 ^ _24642;
  wire _28030 = _28028 ^ _28029;
  wire _28031 = _12463 ^ _8589;
  wire _28032 = _21907 ^ _28031;
  wire _28033 = _28030 ^ _28032;
  wire _28034 = _11390 ^ _81;
  wire _28035 = _19539 ^ _14092;
  wire _28036 = _28034 ^ _28035;
  wire _28037 = uncoded_block[181] ^ uncoded_block[184];
  wire _28038 = _28037 ^ _3284;
  wire _28039 = _11402 ^ _6805;
  wire _28040 = _28038 ^ _28039;
  wire _28041 = _28036 ^ _28040;
  wire _28042 = _28033 ^ _28041;
  wire _28043 = uncoded_block[205] ^ uncoded_block[208];
  wire _28044 = _12479 ^ _28043;
  wire _28045 = _28044 ^ _14104;
  wire _28046 = uncoded_block[217] ^ uncoded_block[220];
  wire _28047 = _3296 ^ _28046;
  wire _28048 = _28047 ^ _10858;
  wire _28049 = _28045 ^ _28048;
  wire _28050 = _6821 ^ _967;
  wire _28051 = _968 ^ _7423;
  wire _28052 = _28050 ^ _28051;
  wire _28053 = _15144 ^ _116;
  wire _28054 = _13609 ^ _6831;
  wire _28055 = _28053 ^ _28054;
  wire _28056 = _28052 ^ _28055;
  wire _28057 = _28049 ^ _28056;
  wire _28058 = _28042 ^ _28057;
  wire _28059 = _28027 ^ _28058;
  wire _28060 = _985 ^ _3320;
  wire _28061 = _28060 ^ _6195;
  wire _28062 = _988 ^ _991;
  wire _28063 = _28062 ^ _20037;
  wire _28064 = _28061 ^ _28063;
  wire _28065 = uncoded_block[295] ^ uncoded_block[302];
  wire _28066 = _995 ^ _28065;
  wire _28067 = uncoded_block[305] ^ uncoded_block[308];
  wire _28068 = _4826 ^ _28067;
  wire _28069 = _28066 ^ _28068;
  wire _28070 = _3337 ^ _15670;
  wire _28071 = _28070 ^ _147;
  wire _28072 = _28069 ^ _28071;
  wire _28073 = _28064 ^ _28072;
  wire _28074 = _149 ^ _6850;
  wire _28075 = _8642 ^ _4837;
  wire _28076 = _28074 ^ _28075;
  wire _28077 = _4126 ^ _3353;
  wire _28078 = _11450 ^ _18621;
  wire _28079 = _28077 ^ _28078;
  wire _28080 = _28076 ^ _28079;
  wire _28081 = _17651 ^ _2602;
  wire _28082 = _6864 ^ _6866;
  wire _28083 = _28081 ^ _28082;
  wire _28084 = _168 ^ _17165;
  wire _28085 = _6873 ^ _4853;
  wire _28086 = _28084 ^ _28085;
  wire _28087 = _28083 ^ _28086;
  wire _28088 = _28080 ^ _28087;
  wire _28089 = _28073 ^ _28088;
  wire _28090 = uncoded_block[381] ^ uncoded_block[385];
  wire _28091 = uncoded_block[386] ^ uncoded_block[388];
  wire _28092 = _28090 ^ _28091;
  wire _28093 = _18629 ^ _28092;
  wire _28094 = _26042 ^ _26925;
  wire _28095 = _17667 ^ _28094;
  wire _28096 = _28093 ^ _28095;
  wire _28097 = _1051 ^ _191;
  wire _28098 = uncoded_block[420] ^ uncoded_block[423];
  wire _28099 = _28098 ^ _8672;
  wire _28100 = _28097 ^ _28099;
  wire _28101 = uncoded_block[427] ^ uncoded_block[430];
  wire _28102 = _28101 ^ _6254;
  wire _28103 = uncoded_block[437] ^ uncoded_block[441];
  wire _28104 = _6255 ^ _28103;
  wire _28105 = _28102 ^ _28104;
  wire _28106 = _28100 ^ _28105;
  wire _28107 = _28096 ^ _28106;
  wire _28108 = uncoded_block[450] ^ uncoded_block[456];
  wire _28109 = _28108 ^ _1873;
  wire _28110 = _6899 ^ _28109;
  wire _28111 = _1874 ^ _1082;
  wire _28112 = _28111 ^ _5591;
  wire _28113 = _28110 ^ _28112;
  wire _28114 = _19128 ^ _21528;
  wire _28115 = _28114 ^ _7519;
  wire _28116 = _13140 ^ _24267;
  wire _28117 = _28115 ^ _28116;
  wire _28118 = _28113 ^ _28117;
  wire _28119 = _28107 ^ _28118;
  wire _28120 = _28089 ^ _28119;
  wire _28121 = _28059 ^ _28120;
  wire _28122 = uncoded_block[511] ^ uncoded_block[517];
  wire _28123 = _3437 ^ _28122;
  wire _28124 = _9841 ^ _1108;
  wire _28125 = _28123 ^ _28124;
  wire _28126 = _20602 ^ _4925;
  wire _28127 = _10384 ^ _1114;
  wire _28128 = _28126 ^ _28127;
  wire _28129 = _28125 ^ _28128;
  wire _28130 = uncoded_block[544] ^ uncoded_block[551];
  wire _28131 = _14197 ^ _28130;
  wire _28132 = uncoded_block[555] ^ uncoded_block[559];
  wire _28133 = uncoded_block[560] ^ uncoded_block[567];
  wire _28134 = _28132 ^ _28133;
  wire _28135 = _28131 ^ _28134;
  wire _28136 = uncoded_block[575] ^ uncoded_block[578];
  wire _28137 = _28136 ^ _5641;
  wire _28138 = _28137 ^ _15246;
  wire _28139 = _28135 ^ _28138;
  wire _28140 = _28129 ^ _28139;
  wire _28141 = _23835 ^ _8149;
  wire _28142 = _4953 ^ _3489;
  wire _28143 = _28141 ^ _28142;
  wire _28144 = _9870 ^ _17232;
  wire _28145 = _28144 ^ _12612;
  wire _28146 = _28143 ^ _28145;
  wire _28147 = uncoded_block[617] ^ uncoded_block[621];
  wire _28148 = _28147 ^ _10979;
  wire _28149 = _1156 ^ _22950;
  wire _28150 = _28148 ^ _28149;
  wire _28151 = _4255 ^ _6338;
  wire _28152 = _25203 ^ _28151;
  wire _28153 = _28150 ^ _28152;
  wire _28154 = _28146 ^ _28153;
  wire _28155 = _28140 ^ _28154;
  wire _28156 = uncoded_block[656] ^ uncoded_block[661];
  wire _28157 = _13187 ^ _28156;
  wire _28158 = uncoded_block[667] ^ uncoded_block[671];
  wire _28159 = _21113 ^ _28158;
  wire _28160 = _28157 ^ _28159;
  wire _28161 = _8760 ^ _1968;
  wire _28162 = _1971 ^ _9891;
  wire _28163 = _28161 ^ _28162;
  wire _28164 = _28160 ^ _28163;
  wire _28165 = _6357 ^ _4272;
  wire _28166 = _28165 ^ _18720;
  wire _28167 = _14255 ^ _8190;
  wire _28168 = _15780 ^ _28167;
  wire _28169 = _28166 ^ _28168;
  wire _28170 = _28164 ^ _28169;
  wire _28171 = _3536 ^ _1194;
  wire _28172 = _8193 ^ _9369;
  wire _28173 = _28171 ^ _28172;
  wire _28174 = _344 ^ _7002;
  wire _28175 = _28174 ^ _26573;
  wire _28176 = _28173 ^ _28175;
  wire _28177 = _23870 ^ _5699;
  wire _28178 = _5704 ^ _24331;
  wire _28179 = _28177 ^ _28178;
  wire _28180 = _7015 ^ _18740;
  wire _28181 = _4301 ^ _10470;
  wire _28182 = _28180 ^ _28181;
  wire _28183 = _28179 ^ _28182;
  wire _28184 = _28176 ^ _28183;
  wire _28185 = _28170 ^ _28184;
  wire _28186 = _28155 ^ _28185;
  wire _28187 = _1218 ^ _1221;
  wire _28188 = _28187 ^ _26146;
  wire _28189 = _12673 ^ _6388;
  wire _28190 = _3574 ^ _11591;
  wire _28191 = _28189 ^ _28190;
  wire _28192 = _28188 ^ _28191;
  wire _28193 = _7029 ^ _3577;
  wire _28194 = _16791 ^ _5042;
  wire _28195 = _28193 ^ _28194;
  wire _28196 = _2026 ^ _1241;
  wire _28197 = uncoded_block[819] ^ uncoded_block[822];
  wire _28198 = _28197 ^ _23896;
  wire _28199 = _28196 ^ _28198;
  wire _28200 = _28195 ^ _28199;
  wire _28201 = _28192 ^ _28200;
  wire _28202 = _12686 ^ _9938;
  wire _28203 = _5057 ^ _2043;
  wire _28204 = _28202 ^ _28203;
  wire _28205 = _11614 ^ _5069;
  wire _28206 = _5065 ^ _28205;
  wire _28207 = _28204 ^ _28206;
  wire _28208 = _22540 ^ _5072;
  wire _28209 = _416 ^ _11620;
  wire _28210 = _28208 ^ _28209;
  wire _28211 = _18770 ^ _15342;
  wire _28212 = _12704 ^ _19735;
  wire _28213 = _28211 ^ _28212;
  wire _28214 = _28210 ^ _28213;
  wire _28215 = _28207 ^ _28214;
  wire _28216 = _28201 ^ _28215;
  wire _28217 = uncoded_block[900] ^ uncoded_block[905];
  wire _28218 = _1278 ^ _28217;
  wire _28219 = _6428 ^ _7665;
  wire _28220 = _28218 ^ _28219;
  wire _28221 = _16315 ^ _4371;
  wire _28222 = _22555 ^ _28221;
  wire _28223 = _28220 ^ _28222;
  wire _28224 = uncoded_block[934] ^ uncoded_block[941];
  wire _28225 = _5773 ^ _28224;
  wire _28226 = _12171 ^ _8271;
  wire _28227 = _28225 ^ _28226;
  wire _28228 = _9975 ^ _12175;
  wire _28229 = _12726 ^ _4385;
  wire _28230 = _28228 ^ _28229;
  wire _28231 = _28227 ^ _28230;
  wire _28232 = _28223 ^ _28231;
  wire _28233 = uncoded_block[974] ^ uncoded_block[977];
  wire _28234 = _10531 ^ _28233;
  wire _28235 = _2100 ^ _7093;
  wire _28236 = _28234 ^ _28235;
  wire _28237 = _8856 ^ _8859;
  wire _28238 = _19275 ^ _13277;
  wire _28239 = _28237 ^ _28238;
  wire _28240 = _28236 ^ _28239;
  wire _28241 = uncoded_block[998] ^ uncoded_block[1000];
  wire _28242 = _28241 ^ _2112;
  wire _28243 = _4405 ^ _2890;
  wire _28244 = _28242 ^ _28243;
  wire _28245 = _8871 ^ _5137;
  wire _28246 = uncoded_block[1024] ^ uncoded_block[1030];
  wire _28247 = _28246 ^ _11668;
  wire _28248 = _28245 ^ _28247;
  wire _28249 = _28244 ^ _28248;
  wire _28250 = _28240 ^ _28249;
  wire _28251 = _28232 ^ _28250;
  wire _28252 = _28216 ^ _28251;
  wire _28253 = _28186 ^ _28252;
  wire _28254 = _28121 ^ _28253;
  wire _28255 = _2908 ^ _11677;
  wire _28256 = uncoded_block[1048] ^ uncoded_block[1051];
  wire _28257 = _28256 ^ _1359;
  wire _28258 = _28255 ^ _28257;
  wire _28259 = _1360 ^ _521;
  wire _28260 = uncoded_block[1064] ^ uncoded_block[1070];
  wire _28261 = _522 ^ _28260;
  wire _28262 = _28259 ^ _28261;
  wire _28263 = _28258 ^ _28262;
  wire _28264 = _5834 ^ _11687;
  wire _28265 = _8323 ^ _28264;
  wire _28266 = uncoded_block[1093] ^ uncoded_block[1098];
  wire _28267 = _13857 ^ _28266;
  wire _28268 = _11142 ^ _8914;
  wire _28269 = _28267 ^ _28268;
  wire _28270 = _28265 ^ _28269;
  wire _28271 = _28263 ^ _28270;
  wire _28272 = _13319 ^ _7133;
  wire _28273 = _3713 ^ _5853;
  wire _28274 = _28272 ^ _28273;
  wire _28275 = _12789 ^ _15894;
  wire _28276 = _4460 ^ _10591;
  wire _28277 = _28275 ^ _28276;
  wire _28278 = _28274 ^ _28277;
  wire _28279 = _10593 ^ _20269;
  wire _28280 = _28279 ^ _7142;
  wire _28281 = _17882 ^ _5190;
  wire _28282 = _1404 ^ _8356;
  wire _28283 = _28281 ^ _28282;
  wire _28284 = _28280 ^ _28283;
  wire _28285 = _28278 ^ _28284;
  wire _28286 = _28271 ^ _28285;
  wire _28287 = _8362 ^ _5195;
  wire _28288 = _4477 ^ _28287;
  wire _28289 = uncoded_block[1179] ^ uncoded_block[1184];
  wire _28290 = _28289 ^ _2200;
  wire _28291 = _6522 ^ _24910;
  wire _28292 = _28290 ^ _28291;
  wire _28293 = _28288 ^ _28292;
  wire _28294 = _22179 ^ _7160;
  wire _28295 = _7162 ^ _2209;
  wire _28296 = _28294 ^ _28295;
  wire _28297 = _2210 ^ _2216;
  wire _28298 = _26694 ^ _12813;
  wire _28299 = _28297 ^ _28298;
  wire _28300 = _28296 ^ _28299;
  wire _28301 = _28293 ^ _28300;
  wire _28302 = _3763 ^ _3765;
  wire _28303 = _13355 ^ _11177;
  wire _28304 = _28302 ^ _28303;
  wire _28305 = _10067 ^ _4509;
  wire _28306 = _22643 ^ _28305;
  wire _28307 = _28304 ^ _28306;
  wire _28308 = _11734 ^ _7778;
  wire _28309 = _28308 ^ _20799;
  wire _28310 = _20801 ^ _3784;
  wire _28311 = _1459 ^ _16419;
  wire _28312 = _28310 ^ _28311;
  wire _28313 = _28309 ^ _28312;
  wire _28314 = _28307 ^ _28313;
  wire _28315 = _28301 ^ _28314;
  wire _28316 = _28286 ^ _28315;
  wire _28317 = uncoded_block[1284] ^ uncoded_block[1286];
  wire _28318 = _10638 ^ _28317;
  wire _28319 = _6561 ^ _1469;
  wire _28320 = _28318 ^ _28319;
  wire _28321 = uncoded_block[1296] ^ uncoded_block[1302];
  wire _28322 = _28321 ^ _3805;
  wire _28323 = _1479 ^ _8992;
  wire _28324 = _28322 ^ _28323;
  wire _28325 = _28320 ^ _28324;
  wire _28326 = uncoded_block[1314] ^ uncoded_block[1319];
  wire _28327 = _28326 ^ _5254;
  wire _28328 = _19377 ^ _3822;
  wire _28329 = _28327 ^ _28328;
  wire _28330 = _9564 ^ _10659;
  wire _28331 = _3042 ^ _5272;
  wire _28332 = _28330 ^ _28331;
  wire _28333 = _28329 ^ _28332;
  wire _28334 = _28325 ^ _28333;
  wire _28335 = uncoded_block[1358] ^ uncoded_block[1362];
  wire _28336 = _28335 ^ _2283;
  wire _28337 = _3052 ^ _8423;
  wire _28338 = _28336 ^ _28337;
  wire _28339 = _7824 ^ _3059;
  wire _28340 = uncoded_block[1391] ^ uncoded_block[1396];
  wire _28341 = _688 ^ _28340;
  wire _28342 = _28339 ^ _28341;
  wire _28343 = _28338 ^ _28342;
  wire _28344 = uncoded_block[1406] ^ uncoded_block[1410];
  wire _28345 = _26749 ^ _28344;
  wire _28346 = _21316 ^ _28345;
  wire _28347 = _5962 ^ _5964;
  wire _28348 = _28347 ^ _20351;
  wire _28349 = _28346 ^ _28348;
  wire _28350 = _28343 ^ _28349;
  wire _28351 = _28334 ^ _28350;
  wire _28352 = _22242 ^ _2318;
  wire _28353 = _20352 ^ _28352;
  wire _28354 = uncoded_block[1441] ^ uncoded_block[1443];
  wire _28355 = _28354 ^ _9033;
  wire _28356 = _3865 ^ _1544;
  wire _28357 = _28355 ^ _28356;
  wire _28358 = _28353 ^ _28357;
  wire _28359 = _5309 ^ _724;
  wire _28360 = _8455 ^ _727;
  wire _28361 = _28359 ^ _28360;
  wire _28362 = _20367 ^ _25423;
  wire _28363 = uncoded_block[1485] ^ uncoded_block[1490];
  wire _28364 = _11807 ^ _28363;
  wire _28365 = _28362 ^ _28364;
  wire _28366 = _28361 ^ _28365;
  wire _28367 = _28358 ^ _28366;
  wire _28368 = _5329 ^ _7864;
  wire _28369 = _28368 ^ _7867;
  wire _28370 = _3894 ^ _24539;
  wire _28371 = _1575 ^ _9621;
  wire _28372 = _28370 ^ _28371;
  wire _28373 = _28369 ^ _28372;
  wire _28374 = _9058 ^ _23194;
  wire _28375 = uncoded_block[1531] ^ uncoded_block[1536];
  wire _28376 = _8474 ^ _28375;
  wire _28377 = _28374 ^ _28376;
  wire _28378 = uncoded_block[1553] ^ uncoded_block[1556];
  wire _28379 = _26792 ^ _28378;
  wire _28380 = _6652 ^ _28379;
  wire _28381 = _28377 ^ _28380;
  wire _28382 = _28373 ^ _28381;
  wire _28383 = _28367 ^ _28382;
  wire _28384 = _28351 ^ _28383;
  wire _28385 = _28316 ^ _28384;
  wire _28386 = uncoded_block[1559] ^ uncoded_block[1563];
  wire _28387 = _11281 ^ _28386;
  wire _28388 = uncoded_block[1566] ^ uncoded_block[1569];
  wire _28389 = _2376 ^ _28388;
  wire _28390 = _28387 ^ _28389;
  wire _28391 = _4645 ^ _10163;
  wire _28392 = _784 ^ _15537;
  wire _28393 = _28391 ^ _28392;
  wire _28394 = _28390 ^ _28393;
  wire _28395 = _15031 ^ _4653;
  wire _28396 = _11292 ^ _11295;
  wire _28397 = _28395 ^ _28396;
  wire _28398 = _11847 ^ _9088;
  wire _28399 = _28398 ^ _16030;
  wire _28400 = _28397 ^ _28399;
  wire _28401 = _28394 ^ _28400;
  wire _28402 = _1632 ^ _24115;
  wire _28403 = _28402 ^ _8508;
  wire _28404 = _14525 ^ _5388;
  wire _28405 = _7914 ^ _11858;
  wire _28406 = _28404 ^ _28405;
  wire _28407 = _28403 ^ _28406;
  wire _28408 = _1649 ^ _4677;
  wire _28409 = _817 ^ _28408;
  wire _28410 = uncoded_block[1656] ^ uncoded_block[1659];
  wire _28411 = _4678 ^ _28410;
  wire _28412 = _28411 ^ _19467;
  wire _28413 = _28409 ^ _28412;
  wire _28414 = _28407 ^ _28413;
  wire _28415 = _28401 ^ _28414;
  wire _28416 = _1656 ^ _5401;
  wire _28417 = _9113 ^ _4693;
  wire _28418 = _28416 ^ _28417;
  wire _28419 = _24130 ^ _837;
  wire _28420 = _28419 ^ _21393;
  wire _28421 = _28418 ^ _28420;
  wire _28422 = _9677 ^ _22772;
  wire _28423 = _20920 ^ _15063;
  wire _28424 = _28422 ^ _28423;
  wire _28425 = uncoded_block[1715] ^ uncoded_block[1721];
  wire _28426 = _12407 ^ _28425;
  wire _28427 = _28426 ^ uncoded_block[1722];
  wire _28428 = _28424 ^ _28427;
  wire _28429 = _28421 ^ _28428;
  wire _28430 = _28415 ^ _28429;
  wire _28431 = _28385 ^ _28430;
  wire _28432 = _28254 ^ _28431;
  wire _28433 = _25948 ^ _31;
  wire _28434 = _8559 ^ _6745;
  wire _28435 = _28433 ^ _28434;
  wire _28436 = _25947 ^ _28435;
  wire _28437 = _27680 ^ _28436;
  wire _28438 = uncoded_block[81] ^ uncoded_block[83];
  wire _28439 = _6109 ^ _28438;
  wire _28440 = _25957 ^ _4741;
  wire _28441 = _28439 ^ _28440;
  wire _28442 = _910 ^ _7986;
  wire _28443 = _28442 ^ _26403;
  wire _28444 = _28441 ^ _28443;
  wire _28445 = _7990 ^ _2495;
  wire _28446 = _6128 ^ _25967;
  wire _28447 = _28445 ^ _28446;
  wire _28448 = _13017 ^ _4754;
  wire _28449 = uncoded_block[132] ^ uncoded_block[139];
  wire _28450 = _28449 ^ _4043;
  wire _28451 = _28448 ^ _28450;
  wire _28452 = _28447 ^ _28451;
  wire _28453 = _28444 ^ _28452;
  wire _28454 = _28437 ^ _28453;
  wire _28455 = _26890 ^ _27719;
  wire _28456 = _27709 ^ _28455;
  wire _28457 = _28454 ^ _28456;
  wire _28458 = _14652 ^ _145;
  wire _28459 = _26013 ^ _28458;
  wire _28460 = _27723 ^ _28459;
  wire _28461 = _146 ^ _1008;
  wire _28462 = _15677 ^ _21947;
  wire _28463 = _28461 ^ _28462;
  wire _28464 = _26021 ^ _2592;
  wire _28465 = _26026 ^ _6859;
  wire _28466 = _28464 ^ _28465;
  wire _28467 = _28463 ^ _28466;
  wire _28468 = _28460 ^ _28467;
  wire _28469 = _19092 ^ _6221;
  wire _28470 = _18155 ^ _28469;
  wire _28471 = _2606 ^ _17163;
  wire _28472 = _17165 ^ _4140;
  wire _28473 = _28471 ^ _28472;
  wire _28474 = _28470 ^ _28473;
  wire _28475 = _10898 ^ _13101;
  wire _28476 = _11999 ^ _6239;
  wire _28477 = _28475 ^ _28476;
  wire _28478 = _26042 ^ _181;
  wire _28479 = _17667 ^ _28478;
  wire _28480 = _28477 ^ _28479;
  wire _28481 = _28474 ^ _28480;
  wire _28482 = _28468 ^ _28481;
  wire _28483 = _2629 ^ _9266;
  wire _28484 = _25147 ^ _28483;
  wire _28485 = _28484 ^ _26050;
  wire _28486 = _2633 ^ _13115;
  wire _28487 = _13117 ^ _1863;
  wire _28488 = _28486 ^ _28487;
  wire _28489 = _5578 ^ _12559;
  wire _28490 = _28489 ^ _10357;
  wire _28491 = _28488 ^ _28490;
  wire _28492 = _28485 ^ _28491;
  wire _28493 = _11491 ^ _9283;
  wire _28494 = _3418 ^ _1083;
  wire _28495 = _28493 ^ _28494;
  wire _28496 = _10361 ^ _28495;
  wire _28497 = _2658 ^ _27767;
  wire _28498 = _28497 ^ _27772;
  wire _28499 = _28496 ^ _28498;
  wire _28500 = _28492 ^ _28499;
  wire _28501 = _28482 ^ _28500;
  wire _28502 = _28457 ^ _28501;
  wire _28503 = uncoded_block[515] ^ uncoded_block[520];
  wire _28504 = _28503 ^ _3445;
  wire _28505 = _20099 ^ _26081;
  wire _28506 = _28504 ^ _28505;
  wire _28507 = _27778 ^ _28506;
  wire _28508 = _6932 ^ _4217;
  wire _28509 = _28508 ^ _26085;
  wire _28510 = _26086 ^ _26091;
  wire _28511 = _28509 ^ _28510;
  wire _28512 = _28507 ^ _28511;
  wire _28513 = _15747 ^ _4946;
  wire _28514 = _4225 ^ _28513;
  wire _28515 = _8733 ^ _13705;
  wire _28516 = _1938 ^ _15247;
  wire _28517 = _28515 ^ _28516;
  wire _28518 = _28514 ^ _28517;
  wire _28519 = uncoded_block[599] ^ uncoded_block[604];
  wire _28520 = _2706 ^ _28519;
  wire _28521 = _28520 ^ _27794;
  wire _28522 = _8745 ^ _3495;
  wire _28523 = _28522 ^ _26109;
  wire _28524 = _28521 ^ _28523;
  wire _28525 = _28518 ^ _28524;
  wire _28526 = _28512 ^ _28525;
  wire _28527 = _4249 ^ _4255;
  wire _28528 = _2727 ^ _4972;
  wire _28529 = _28527 ^ _28528;
  wire _28530 = _26112 ^ _301;
  wire _28531 = _302 ^ _14755;
  wire _28532 = _28530 ^ _28531;
  wire _28533 = _28529 ^ _28532;
  wire _28534 = _4261 ^ _12630;
  wire _28535 = _26117 ^ _1177;
  wire _28536 = _28534 ^ _28535;
  wire _28537 = _26995 ^ _15281;
  wire _28538 = _24312 ^ _28537;
  wire _28539 = _28536 ^ _28538;
  wire _28540 = _28533 ^ _28539;
  wire _28541 = _1974 ^ _4987;
  wire _28542 = _19195 ^ _11562;
  wire _28543 = _28541 ^ _28542;
  wire _28544 = _6361 ^ _336;
  wire _28545 = _4996 ^ _2762;
  wire _28546 = _28544 ^ _28545;
  wire _28547 = _28543 ^ _28546;
  wire _28548 = _6374 ^ _6999;
  wire _28549 = _26130 ^ _28548;
  wire _28550 = _27818 ^ _1207;
  wire _28551 = _28550 ^ _22506;
  wire _28552 = _28549 ^ _28551;
  wire _28553 = _28547 ^ _28552;
  wire _28554 = _28540 ^ _28553;
  wire _28555 = _28526 ^ _28554;
  wire _28556 = _4295 ^ _27827;
  wire _28557 = _28556 ^ _18270;
  wire _28558 = _28557 ^ _26147;
  wire _28559 = uncoded_block[795] ^ uncoded_block[799];
  wire _28560 = _28559 ^ _385;
  wire _28561 = _1235 ^ _14287;
  wire _28562 = _28560 ^ _28561;
  wire _28563 = _26150 ^ _28562;
  wire _28564 = _28558 ^ _28563;
  wire _28565 = _2806 ^ _22525;
  wire _28566 = _27843 ^ _23450;
  wire _28567 = _28565 ^ _28566;
  wire _28568 = _27846 ^ _12138;
  wire _28569 = _5057 ^ _14812;
  wire _28570 = _28568 ^ _28569;
  wire _28571 = _28567 ^ _28570;
  wire _28572 = _11610 ^ _12146;
  wire _28573 = _2046 ^ _20692;
  wire _28574 = _28572 ^ _28573;
  wire _28575 = _9950 ^ _14306;
  wire _28576 = _28574 ^ _28575;
  wire _28577 = _28571 ^ _28576;
  wire _28578 = _28564 ^ _28577;
  wire _28579 = _417 ^ _16815;
  wire _28580 = _28579 ^ _26175;
  wire _28581 = _4355 ^ _2843;
  wire _28582 = _26176 ^ _28581;
  wire _28583 = _28580 ^ _28582;
  wire _28584 = _10508 ^ _8254;
  wire _28585 = _11067 ^ _7665;
  wire _28586 = _28584 ^ _28585;
  wire _28587 = _17820 ^ _448;
  wire _28588 = _1299 ^ _452;
  wire _28589 = _28587 ^ _28588;
  wire _28590 = _28586 ^ _28589;
  wire _28591 = _28583 ^ _28590;
  wire _28592 = _8274 ^ _461;
  wire _28593 = _24385 ^ _28592;
  wire _28594 = _2090 ^ _4385;
  wire _28595 = _26193 ^ _26197;
  wire _28596 = _28594 ^ _28595;
  wire _28597 = _28593 ^ _28596;
  wire _28598 = _470 ^ _5789;
  wire _28599 = _2100 ^ _13822;
  wire _28600 = _28598 ^ _28599;
  wire _28601 = _8856 ^ _16338;
  wire _28602 = _28601 ^ _19276;
  wire _28603 = _28600 ^ _28602;
  wire _28604 = _28597 ^ _28603;
  wire _28605 = _28591 ^ _28604;
  wire _28606 = _28578 ^ _28605;
  wire _28607 = _28555 ^ _28606;
  wire _28608 = _28502 ^ _28607;
  wire _28609 = _11101 ^ _9991;
  wire _28610 = _28609 ^ _7099;
  wire _28611 = _5131 ^ _12750;
  wire _28612 = _5137 ^ _27081;
  wire _28613 = _28611 ^ _28612;
  wire _28614 = _28610 ^ _28613;
  wire _28615 = uncoded_block[1058] ^ uncoded_block[1065];
  wire _28616 = _28615 ^ _8889;
  wire _28617 = _26218 ^ _28616;
  wire _28618 = _27884 ^ _28617;
  wire _28619 = _28614 ^ _28618;
  wire _28620 = _8892 ^ _5832;
  wire _28621 = _28620 ^ _26226;
  wire _28622 = _545 ^ _13318;
  wire _28623 = _13319 ^ _5175;
  wire _28624 = _28622 ^ _28623;
  wire _28625 = _28621 ^ _28624;
  wire _28626 = _23981 ^ _15896;
  wire _28627 = _8929 ^ _567;
  wire _28628 = _28626 ^ _28627;
  wire _28629 = _9500 ^ _27105;
  wire _28630 = _26241 ^ _28629;
  wire _28631 = _28628 ^ _28630;
  wire _28632 = _28625 ^ _28631;
  wire _28633 = _28619 ^ _28632;
  wire _28634 = _8362 ^ _5872;
  wire _28635 = _17888 ^ _28634;
  wire _28636 = _3742 ^ _4486;
  wire _28637 = _2200 ^ _2971;
  wire _28638 = _28636 ^ _28637;
  wire _28639 = _28635 ^ _28638;
  wire _28640 = _13347 ^ _7160;
  wire _28641 = _8370 ^ _24456;
  wire _28642 = _28640 ^ _28641;
  wire _28643 = _23544 ^ _27911;
  wire _28644 = _27912 ^ _11180;
  wire _28645 = _28643 ^ _28644;
  wire _28646 = _28642 ^ _28645;
  wire _28647 = _28639 ^ _28646;
  wire _28648 = _3771 ^ _16915;
  wire _28649 = _27129 ^ _13365;
  wire _28650 = _28648 ^ _28649;
  wire _28651 = _2232 ^ _2998;
  wire _28652 = _2235 ^ _7780;
  wire _28653 = _28651 ^ _28652;
  wire _28654 = _28650 ^ _28653;
  wire _28655 = _8970 ^ _4516;
  wire _28656 = _2239 ^ _628;
  wire _28657 = _28655 ^ _28656;
  wire _28658 = _23123 ^ _18866;
  wire _28659 = _19364 ^ _28658;
  wire _28660 = _28657 ^ _28659;
  wire _28661 = _28654 ^ _28660;
  wire _28662 = _28647 ^ _28661;
  wire _28663 = _28633 ^ _28662;
  wire _28664 = _8399 ^ _26274;
  wire _28665 = uncoded_block[1303] ^ uncoded_block[1308];
  wire _28666 = _16424 ^ _28665;
  wire _28667 = _28664 ^ _28666;
  wire _28668 = _14430 ^ _21748;
  wire _28669 = _28668 ^ _26280;
  wire _28670 = _28667 ^ _28669;
  wire _28671 = _8411 ^ _11764;
  wire _28672 = _2268 ^ _660;
  wire _28673 = _28671 ^ _28672;
  wire _28674 = _661 ^ _4553;
  wire _28675 = _5937 ^ _3042;
  wire _28676 = _28674 ^ _28675;
  wire _28677 = _28673 ^ _28676;
  wire _28678 = _28670 ^ _28677;
  wire _28679 = uncoded_block[1356] ^ uncoded_block[1360];
  wire _28680 = _5272 ^ _28679;
  wire _28681 = uncoded_block[1363] ^ uncoded_block[1372];
  wire _28682 = _28681 ^ _9572;
  wire _28683 = _28680 ^ _28682;
  wire _28684 = _12305 ^ _27160;
  wire _28685 = _10108 ^ _3838;
  wire _28686 = _28684 ^ _28685;
  wire _28687 = _28683 ^ _28686;
  wire _28688 = _13412 ^ _21774;
  wire _28689 = _5955 ^ _3841;
  wire _28690 = _28688 ^ _28689;
  wire _28691 = _4578 ^ _10113;
  wire _28692 = _28691 ^ _5963;
  wire _28693 = _28690 ^ _28692;
  wire _28694 = _28687 ^ _28693;
  wire _28695 = _28678 ^ _28694;
  wire _28696 = _26302 ^ _26304;
  wire _28697 = _5968 ^ _9591;
  wire _28698 = _2314 ^ _8449;
  wire _28699 = _28697 ^ _28698;
  wire _28700 = _28696 ^ _28699;
  wire _28701 = _26310 ^ _26312;
  wire _28702 = _27945 ^ _27949;
  wire _28703 = _28701 ^ _28702;
  wire _28704 = _28700 ^ _28703;
  wire _28705 = _2349 ^ _25426;
  wire _28706 = _28705 ^ _24079;
  wire _28707 = _2352 ^ _747;
  wire _28708 = _28707 ^ _11265;
  wire _28709 = _28706 ^ _28708;
  wire _28710 = _15002 ^ _7875;
  wire _28711 = _28710 ^ _27192;
  wire _28712 = _27193 ^ _9633;
  wire _28713 = _28711 ^ _28712;
  wire _28714 = _28709 ^ _28713;
  wire _28715 = _28704 ^ _28714;
  wire _28716 = _28695 ^ _28715;
  wire _28717 = _28663 ^ _28716;
  wire _28718 = _16997 ^ _27203;
  wire _28719 = _26332 ^ _28718;
  wire _28720 = _27204 ^ _27207;
  wire _28721 = _27208 ^ _27210;
  wire _28722 = _28720 ^ _28721;
  wire _28723 = _28719 ^ _28722;
  wire _28724 = uncoded_block[1621] ^ uncoded_block[1632];
  wire _28725 = _28724 ^ _7306;
  wire _28726 = _12944 ^ _28725;
  wire _28727 = uncoded_block[1639] ^ uncoded_block[1642];
  wire _28728 = _28727 ^ _2412;
  wire _28729 = _12387 ^ _3174;
  wire _28730 = _28728 ^ _28729;
  wire _28731 = _28726 ^ _28730;
  wire _28732 = _4680 ^ _1654;
  wire _28733 = _25476 ^ _6700;
  wire _28734 = _28732 ^ _28733;
  wire _28735 = _830 ^ _12398;
  wire _28736 = _28735 ^ _22307;
  wire _28737 = _28734 ^ _28736;
  wire _28738 = _28731 ^ _28737;
  wire _28739 = _28723 ^ _28738;
  wire _28740 = _27985 ^ _26367;
  wire _28741 = _28740 ^ _26371;
  wire _28742 = _28741 ^ _26374;
  wire _28743 = _28739 ^ _28742;
  wire _28744 = _28717 ^ _28743;
  wire _28745 = _28608 ^ _28744;
  wire _28746 = _19959 ^ _6083;
  wire _28747 = _2 ^ _28746;
  wire _28748 = _3216 ^ _9692;
  wire _28749 = _3217 ^ _9139;
  wire _28750 = _28748 ^ _28749;
  wire _28751 = _28747 ^ _28750;
  wire _28752 = uncoded_block[26] ^ uncoded_block[31];
  wire _28753 = uncoded_block[32] ^ uncoded_block[36];
  wire _28754 = _28752 ^ _28753;
  wire _28755 = _10796 ^ _23;
  wire _28756 = _28754 ^ _28755;
  wire _28757 = uncoded_block[54] ^ uncoded_block[59];
  wire _28758 = _4014 ^ _28757;
  wire _28759 = _18068 ^ _28758;
  wire _28760 = _28756 ^ _28759;
  wire _28761 = _28751 ^ _28760;
  wire _28762 = _2472 ^ _2474;
  wire _28763 = _12435 ^ _7367;
  wire _28764 = _28762 ^ _28763;
  wire _28765 = uncoded_block[78] ^ uncoded_block[80];
  wire _28766 = _5442 ^ _28765;
  wire _28767 = uncoded_block[82] ^ uncoded_block[90];
  wire _28768 = _28767 ^ _907;
  wire _28769 = _28766 ^ _28768;
  wire _28770 = _28764 ^ _28769;
  wire _28771 = _1719 ^ _4028;
  wire _28772 = _17584 ^ _6123;
  wire _28773 = _28771 ^ _28772;
  wire _28774 = _6763 ^ _2497;
  wire _28775 = _1729 ^ _20961;
  wire _28776 = _28774 ^ _28775;
  wire _28777 = _28773 ^ _28776;
  wire _28778 = _28770 ^ _28777;
  wire _28779 = _28761 ^ _28778;
  wire _28780 = _1733 ^ _15112;
  wire _28781 = uncoded_block[140] ^ uncoded_block[147];
  wire _28782 = _9729 ^ _28781;
  wire _28783 = _28780 ^ _28782;
  wire _28784 = _14082 ^ _26415;
  wire _28785 = _73 ^ _20975;
  wire _28786 = _28784 ^ _28785;
  wire _28787 = _28783 ^ _28786;
  wire _28788 = uncoded_block[164] ^ uncoded_block[169];
  wire _28789 = _28788 ^ _15123;
  wire _28790 = _940 ^ _1757;
  wire _28791 = _28789 ^ _28790;
  wire _28792 = _4067 ^ _17112;
  wire _28793 = _27706 ^ _28792;
  wire _28794 = _28791 ^ _28793;
  wire _28795 = _28787 ^ _28794;
  wire _28796 = uncoded_block[202] ^ uncoded_block[209];
  wire _28797 = uncoded_block[211] ^ uncoded_block[216];
  wire _28798 = _28796 ^ _28797;
  wire _28799 = _14105 ^ _5497;
  wire _28800 = _28798 ^ _28799;
  wire _28801 = _23300 ^ _6824;
  wire _28802 = _25101 ^ _28801;
  wire _28803 = _28800 ^ _28802;
  wire _28804 = _10860 ^ _4799;
  wire _28805 = uncoded_block[250] ^ uncoded_block[255];
  wire _28806 = _28805 ^ _13055;
  wire _28807 = _28804 ^ _28806;
  wire _28808 = _6185 ^ _977;
  wire _28809 = _11421 ^ _128;
  wire _28810 = _28808 ^ _28809;
  wire _28811 = _28807 ^ _28810;
  wire _28812 = _28803 ^ _28811;
  wire _28813 = _28795 ^ _28812;
  wire _28814 = _28779 ^ _28813;
  wire _28815 = _4813 ^ _10303;
  wire _28816 = _28815 ^ _5516;
  wire _28817 = uncoded_block[290] ^ uncoded_block[294];
  wire _28818 = _28817 ^ _1806;
  wire _28819 = _13066 ^ _28818;
  wire _28820 = _28816 ^ _28819;
  wire _28821 = _1811 ^ _8056;
  wire _28822 = _17642 ^ _4118;
  wire _28823 = _28821 ^ _28822;
  wire _28824 = _6209 ^ _1014;
  wire _28825 = _2586 ^ _1821;
  wire _28826 = _28824 ^ _28825;
  wire _28827 = _28823 ^ _28826;
  wire _28828 = _28820 ^ _28827;
  wire _28829 = _1017 ^ _4840;
  wire _28830 = _11450 ^ _159;
  wire _28831 = _28829 ^ _28830;
  wire _28832 = _5541 ^ _1028;
  wire _28833 = _28832 ^ _3363;
  wire _28834 = _28831 ^ _28833;
  wire _28835 = _12530 ^ _5548;
  wire _28836 = _13093 ^ _4140;
  wire _28837 = _28835 ^ _28836;
  wire _28838 = uncoded_block[374] ^ uncoded_block[377];
  wire _28839 = _28838 ^ _2612;
  wire _28840 = _4149 ^ _176;
  wire _28841 = _28839 ^ _28840;
  wire _28842 = _28837 ^ _28841;
  wire _28843 = _28834 ^ _28842;
  wire _28844 = _28828 ^ _28843;
  wire _28845 = uncoded_block[395] ^ uncoded_block[399];
  wire _28846 = _28845 ^ _5559;
  wire _28847 = _28846 ^ _5562;
  wire _28848 = _8091 ^ _4871;
  wire _28849 = _18175 ^ _4164;
  wire _28850 = _28848 ^ _28849;
  wire _28851 = _28847 ^ _28850;
  wire _28852 = _2638 ^ _9271;
  wire _28853 = _199 ^ _28852;
  wire _28854 = _4169 ^ _21049;
  wire _28855 = _206 ^ _1866;
  wire _28856 = _28854 ^ _28855;
  wire _28857 = _28853 ^ _28856;
  wire _28858 = _28851 ^ _28857;
  wire _28859 = _3415 ^ _21057;
  wire _28860 = _17186 ^ _28859;
  wire _28861 = uncoded_block[464] ^ uncoded_block[469];
  wire _28862 = _28861 ^ _3418;
  wire _28863 = _4188 ^ _2657;
  wire _28864 = _28862 ^ _28863;
  wire _28865 = _28860 ^ _28864;
  wire _28866 = uncoded_block[478] ^ uncoded_block[483];
  wire _28867 = _28866 ^ _4897;
  wire _28868 = _224 ^ _8115;
  wire _28869 = _28867 ^ _28868;
  wire _28870 = _4905 ^ _6279;
  wire _28871 = _18193 ^ _28870;
  wire _28872 = _28869 ^ _28871;
  wire _28873 = _28865 ^ _28872;
  wire _28874 = _28858 ^ _28873;
  wire _28875 = _28844 ^ _28874;
  wire _28876 = _28814 ^ _28875;
  wire _28877 = uncoded_block[514] ^ uncoded_block[523];
  wire _28878 = _9295 ^ _28877;
  wire _28879 = uncoded_block[529] ^ uncoded_block[533];
  wire _28880 = _28879 ^ _1905;
  wire _28881 = _28878 ^ _28880;
  wire _28882 = uncoded_block[541] ^ uncoded_block[544];
  wire _28883 = _4217 ^ _28882;
  wire _28884 = _28883 ^ _15235;
  wire _28885 = _28881 ^ _28884;
  wire _28886 = _247 ^ _4937;
  wire _28887 = uncoded_block[566] ^ uncoded_block[571];
  wire _28888 = _10395 ^ _28887;
  wire _28889 = _28886 ^ _28888;
  wire _28890 = _6945 ^ _265;
  wire _28891 = uncoded_block[584] ^ uncoded_block[588];
  wire _28892 = _28891 ^ _4234;
  wire _28893 = _28890 ^ _28892;
  wire _28894 = _28889 ^ _28893;
  wire _28895 = _28885 ^ _28894;
  wire _28896 = uncoded_block[598] ^ uncoded_block[602];
  wire _28897 = _6952 ^ _28896;
  wire _28898 = _8152 ^ _6323;
  wire _28899 = _28897 ^ _28898;
  wire _28900 = _6957 ^ _5652;
  wire _28901 = uncoded_block[625] ^ uncoded_block[630];
  wire _28902 = _16238 ^ _28901;
  wire _28903 = _28900 ^ _28902;
  wire _28904 = _28899 ^ _28903;
  wire _28905 = uncoded_block[632] ^ uncoded_block[637];
  wire _28906 = _28905 ^ _4255;
  wire _28907 = _28906 ^ _28528;
  wire _28908 = uncoded_block[651] ^ uncoded_block[653];
  wire _28909 = _8165 ^ _28908;
  wire _28910 = _12629 ^ _3513;
  wire _28911 = _28909 ^ _28910;
  wire _28912 = _28907 ^ _28911;
  wire _28913 = _28904 ^ _28912;
  wire _28914 = _28895 ^ _28913;
  wire _28915 = uncoded_block[665] ^ uncoded_block[670];
  wire _28916 = _14238 ^ _28915;
  wire _28917 = _12087 ^ _6352;
  wire _28918 = _28916 ^ _28917;
  wire _28919 = _2750 ^ _26557;
  wire _28920 = _2755 ^ _18719;
  wire _28921 = _28919 ^ _28920;
  wire _28922 = _28918 ^ _28921;
  wire _28923 = _11564 ^ _19688;
  wire _28924 = _15286 ^ _28923;
  wire _28925 = _340 ^ _22049;
  wire _28926 = _28171 ^ _28925;
  wire _28927 = _28924 ^ _28926;
  wire _28928 = _28922 ^ _28927;
  wire _28929 = _11006 ^ _1203;
  wire _28930 = uncoded_block[742] ^ uncoded_block[748];
  wire _28931 = _1206 ^ _28930;
  wire _28932 = _28929 ^ _28931;
  wire _28933 = uncoded_block[764] ^ uncoded_block[767];
  wire _28934 = _2781 ^ _28933;
  wire _28935 = _2779 ^ _28934;
  wire _28936 = _28932 ^ _28935;
  wire _28937 = _1218 ^ _12114;
  wire _28938 = uncoded_block[778] ^ uncoded_block[784];
  wire _28939 = _2792 ^ _28938;
  wire _28940 = _28937 ^ _28939;
  wire _28941 = _8215 ^ _1225;
  wire _28942 = _5035 ^ _5039;
  wire _28943 = _28941 ^ _28942;
  wire _28944 = _28940 ^ _28943;
  wire _28945 = _28936 ^ _28944;
  wire _28946 = _28928 ^ _28945;
  wire _28947 = _28914 ^ _28946;
  wire _28948 = _15814 ^ _15318;
  wire _28949 = _11030 ^ _1241;
  wire _28950 = _28948 ^ _28949;
  wire _28951 = _2029 ^ _14291;
  wire _28952 = _7039 ^ _11042;
  wire _28953 = _28951 ^ _28952;
  wire _28954 = _28950 ^ _28953;
  wire _28955 = uncoded_block[842] ^ uncoded_block[850];
  wire _28956 = _28955 ^ _8237;
  wire _28957 = _28956 ^ _27036;
  wire _28958 = _5072 ^ _9412;
  wire _28959 = _1267 ^ _28958;
  wire _28960 = _28957 ^ _28959;
  wire _28961 = _28954 ^ _28960;
  wire _28962 = uncoded_block[887] ^ uncoded_block[891];
  wire _28963 = _28962 ^ _3614;
  wire _28964 = _27044 ^ _28963;
  wire _28965 = uncoded_block[900] ^ uncoded_block[902];
  wire _28966 = _14829 ^ _28965;
  wire _28967 = _4360 ^ _2070;
  wire _28968 = _28966 ^ _28967;
  wire _28969 = _28964 ^ _28968;
  wire _28970 = _7665 ^ _5092;
  wire _28971 = _28970 ^ _3633;
  wire _28972 = _1295 ^ _4371;
  wire _28973 = _28972 ^ _20212;
  wire _28974 = _28971 ^ _28973;
  wire _28975 = _28969 ^ _28974;
  wire _28976 = _28961 ^ _28975;
  wire _28977 = _21191 ^ _14329;
  wire _28978 = _18783 ^ _28977;
  wire _28979 = _1308 ^ _5108;
  wire _28980 = uncoded_block[976] ^ uncoded_block[980];
  wire _28981 = _11649 ^ _28980;
  wire _28982 = _28979 ^ _28981;
  wire _28983 = _28978 ^ _28982;
  wire _28984 = uncoded_block[982] ^ uncoded_block[989];
  wire _28985 = uncoded_block[994] ^ uncoded_block[998];
  wire _28986 = _28984 ^ _28985;
  wire _28987 = _9449 ^ _6459;
  wire _28988 = _28986 ^ _28987;
  wire _28989 = uncoded_block[1015] ^ uncoded_block[1019];
  wire _28990 = _2117 ^ _28989;
  wire _28991 = _2120 ^ _4415;
  wire _28992 = _28990 ^ _28991;
  wire _28993 = _28988 ^ _28992;
  wire _28994 = _28983 ^ _28993;
  wire _28995 = uncoded_block[1033] ^ uncoded_block[1038];
  wire _28996 = _28995 ^ _15387;
  wire _28997 = _10007 ^ _28996;
  wire _28998 = _14866 ^ _19296;
  wire _28999 = _28997 ^ _28998;
  wire _29000 = _9465 ^ _10566;
  wire _29001 = _5825 ^ _14357;
  wire _29002 = _29000 ^ _29001;
  wire _29003 = _5831 ^ _8895;
  wire _29004 = _11123 ^ _29003;
  wire _29005 = _29002 ^ _29004;
  wire _29006 = _28999 ^ _29005;
  wire _29007 = _28994 ^ _29006;
  wire _29008 = _28976 ^ _29007;
  wire _29009 = _28947 ^ _29008;
  wire _29010 = _28876 ^ _29009;
  wire _29011 = _11126 ^ _2928;
  wire _29012 = _3696 ^ _8906;
  wire _29013 = _29011 ^ _29012;
  wire _29014 = uncoded_block[1092] ^ uncoded_block[1095];
  wire _29015 = _29014 ^ _5843;
  wire _29016 = _13316 ^ _3707;
  wire _29017 = _29015 ^ _29016;
  wire _29018 = _29013 ^ _29017;
  wire _29019 = _7133 ^ _8339;
  wire _29020 = _4452 ^ _29019;
  wire _29021 = _15894 ^ _23981;
  wire _29022 = _4456 ^ _29021;
  wire _29023 = _29020 ^ _29022;
  wire _29024 = _29018 ^ _29023;
  wire _29025 = _8346 ^ _2179;
  wire _29026 = _3724 ^ _6505;
  wire _29027 = _29025 ^ _29026;
  wire _29028 = uncoded_block[1158] ^ uncoded_block[1160];
  wire _29029 = _6507 ^ _29028;
  wire _29030 = _1407 ^ _15907;
  wire _29031 = _29029 ^ _29030;
  wire _29032 = _29027 ^ _29031;
  wire _29033 = _1408 ^ _17392;
  wire _29034 = _585 ^ _2193;
  wire _29035 = _29033 ^ _29034;
  wire _29036 = _8944 ^ _12808;
  wire _29037 = _29036 ^ _25349;
  wire _29038 = _29035 ^ _29037;
  wire _29039 = _29032 ^ _29038;
  wire _29040 = _29024 ^ _29039;
  wire _29041 = _14398 ^ _11721;
  wire _29042 = _2207 ^ _1425;
  wire _29043 = _29041 ^ _29042;
  wire _29044 = _26694 ^ _1432;
  wire _29045 = uncoded_block[1221] ^ uncoded_block[1225];
  wire _29046 = uncoded_block[1227] ^ uncoded_block[1230];
  wire _29047 = _29045 ^ _29046;
  wire _29048 = _29044 ^ _29047;
  wire _29049 = _29043 ^ _29048;
  wire _29050 = uncoded_block[1235] ^ uncoded_block[1240];
  wire _29051 = _5219 ^ _29050;
  wire _29052 = _16408 ^ _6538;
  wire _29053 = _29051 ^ _29052;
  wire _29054 = _24471 ^ _3784;
  wire _29055 = _16917 ^ _29054;
  wire _29056 = _29053 ^ _29055;
  wire _29057 = _29049 ^ _29056;
  wire _29058 = _6550 ^ _23559;
  wire _29059 = _29058 ^ _7793;
  wire _29060 = _12834 ^ _638;
  wire _29061 = _5243 ^ _4529;
  wire _29062 = _29060 ^ _29061;
  wire _29063 = _29059 ^ _29062;
  wire _29064 = _3801 ^ _4531;
  wire _29065 = uncoded_block[1302] ^ uncoded_block[1308];
  wire _29066 = _18870 ^ _29065;
  wire _29067 = _29064 ^ _29066;
  wire _29068 = uncoded_block[1309] ^ uncoded_block[1316];
  wire _29069 = _29068 ^ _21293;
  wire _29070 = _2265 ^ _3032;
  wire _29071 = _29069 ^ _29070;
  wire _29072 = _29067 ^ _29071;
  wire _29073 = _29063 ^ _29072;
  wire _29074 = _29057 ^ _29073;
  wire _29075 = _29040 ^ _29074;
  wire _29076 = _5261 ^ _11215;
  wire _29077 = _23140 ^ _29076;
  wire _29078 = _14442 ^ _3042;
  wire _29079 = _14956 ^ _12300;
  wire _29080 = _29078 ^ _29079;
  wire _29081 = _29077 ^ _29080;
  wire _29082 = _11776 ^ _8423;
  wire _29083 = uncoded_block[1380] ^ uncoded_block[1384];
  wire _29084 = _20334 ^ _29083;
  wire _29085 = _29082 ^ _29084;
  wire _29086 = _12311 ^ _12867;
  wire _29087 = _29086 ^ _4570;
  wire _29088 = _29085 ^ _29087;
  wire _29089 = _29081 ^ _29088;
  wire _29090 = uncoded_block[1398] ^ uncoded_block[1402];
  wire _29091 = _3065 ^ _29090;
  wire _29092 = _3846 ^ _15489;
  wire _29093 = _29091 ^ _29092;
  wire _29094 = _8438 ^ _6607;
  wire _29095 = uncoded_block[1421] ^ uncoded_block[1426];
  wire _29096 = _29095 ^ _9590;
  wire _29097 = _29094 ^ _29096;
  wire _29098 = _29093 ^ _29097;
  wire _29099 = _22242 ^ _13432;
  wire _29100 = _6613 ^ _3084;
  wire _29101 = _29099 ^ _29100;
  wire _29102 = _3868 ^ _724;
  wire _29103 = _4595 ^ _29102;
  wire _29104 = _29101 ^ _29103;
  wire _29105 = _29098 ^ _29104;
  wire _29106 = _29089 ^ _29105;
  wire _29107 = _2336 ^ _1550;
  wire _29108 = _11255 ^ _1555;
  wire _29109 = _29107 ^ _29108;
  wire _29110 = _1556 ^ _12342;
  wire _29111 = uncoded_block[1488] ^ uncoded_block[1495];
  wire _29112 = _1562 ^ _29111;
  wire _29113 = _29110 ^ _29112;
  wire _29114 = _29109 ^ _29113;
  wire _29115 = _6635 ^ _11813;
  wire _29116 = _7257 ^ _29115;
  wire _29117 = _15002 ^ _9053;
  wire _29118 = _751 ^ _754;
  wire _29119 = _29117 ^ _29118;
  wire _29120 = _29116 ^ _29119;
  wire _29121 = _29114 ^ _29120;
  wire _29122 = _7269 ^ _8473;
  wire _29123 = _3123 ^ _24994;
  wire _29124 = _29122 ^ _29123;
  wire _29125 = uncoded_block[1541] ^ uncoded_block[1545];
  wire _29126 = _3908 ^ _29125;
  wire _29127 = _8477 ^ _29126;
  wire _29128 = _29124 ^ _29127;
  wire _29129 = uncoded_block[1559] ^ uncoded_block[1565];
  wire _29130 = _7277 ^ _29129;
  wire _29131 = _8483 ^ _29130;
  wire _29132 = _4644 ^ _25895;
  wire _29133 = _15026 ^ _13478;
  wire _29134 = _29132 ^ _29133;
  wire _29135 = _29131 ^ _29134;
  wire _29136 = _29128 ^ _29135;
  wire _29137 = _29121 ^ _29136;
  wire _29138 = _29106 ^ _29137;
  wire _29139 = _29075 ^ _29138;
  wire _29140 = _1612 ^ _21826;
  wire _29141 = _2394 ^ _11295;
  wire _29142 = _29140 ^ _29141;
  wire _29143 = _24111 ^ _20896;
  wire _29144 = _29142 ^ _29143;
  wire _29145 = _804 ^ _7298;
  wire _29146 = _10182 ^ _29145;
  wire _29147 = uncoded_block[1630] ^ uncoded_block[1634];
  wire _29148 = _29147 ^ _2407;
  wire _29149 = _7301 ^ _29148;
  wire _29150 = _29146 ^ _29149;
  wire _29151 = _29144 ^ _29150;
  wire _29152 = _5394 ^ _3172;
  wire _29153 = _9106 ^ _13508;
  wire _29154 = _29152 ^ _29153;
  wire _29155 = _823 ^ _19466;
  wire _29156 = _29155 ^ _14537;
  wire _29157 = _29154 ^ _29156;
  wire _29158 = _11319 ^ _11321;
  wire _29159 = _9113 ^ _16058;
  wire _29160 = _29158 ^ _29159;
  wire _29161 = _10205 ^ _6066;
  wire _29162 = uncoded_block[1695] ^ uncoded_block[1699];
  wire _29163 = _29162 ^ _24137;
  wire _29164 = _29161 ^ _29163;
  wire _29165 = _29160 ^ _29164;
  wire _29166 = _29157 ^ _29165;
  wire _29167 = _29151 ^ _29166;
  wire _29168 = _8535 ^ _848;
  wire _29169 = _3980 ^ _854;
  wire _29170 = _29168 ^ _29169;
  wire _29171 = _20923 ^ uncoded_block[1720];
  wire _29172 = _29170 ^ _29171;
  wire _29173 = _29167 ^ _29172;
  wire _29174 = _29139 ^ _29173;
  wire _29175 = _29010 ^ _29174;
  wire _29176 = _18539 ^ _6080;
  wire _29177 = _3993 ^ _3995;
  wire _29178 = _29176 ^ _29177;
  wire _29179 = _7956 ^ _9692;
  wire _29180 = _10 ^ _11344;
  wire _29181 = _29179 ^ _29180;
  wire _29182 = _29178 ^ _29181;
  wire _29183 = _875 ^ _3227;
  wire _29184 = _29183 ^ _2467;
  wire _29185 = _885 ^ _13547;
  wire _29186 = _1700 ^ _23256;
  wire _29187 = _29185 ^ _29186;
  wire _29188 = _29184 ^ _29187;
  wire _29189 = _29182 ^ _29188;
  wire _29190 = _897 ^ _1712;
  wire _29191 = _14056 ^ _29190;
  wire _29192 = _901 ^ _18077;
  wire _29193 = _19515 ^ _7375;
  wire _29194 = _29192 ^ _29193;
  wire _29195 = _29191 ^ _29194;
  wire _29196 = _17083 ^ _19028;
  wire _29197 = uncoded_block[116] ^ uncoded_block[131];
  wire _29198 = _10816 ^ _29197;
  wire _29199 = _1736 ^ _6136;
  wire _29200 = _29198 ^ _29199;
  wire _29201 = _29196 ^ _29200;
  wire _29202 = _29195 ^ _29201;
  wire _29203 = _29189 ^ _29202;
  wire _29204 = uncoded_block[146] ^ uncoded_block[151];
  wire _29205 = _2511 ^ _29204;
  wire _29206 = _9186 ^ _24182;
  wire _29207 = _29205 ^ _29206;
  wire _29208 = uncoded_block[161] ^ uncoded_block[166];
  wire _29209 = _29208 ^ _79;
  wire _29210 = uncoded_block[169] ^ uncoded_block[174];
  wire _29211 = _29210 ^ _6149;
  wire _29212 = _29209 ^ _29211;
  wire _29213 = _29207 ^ _29212;
  wire _29214 = _10843 ^ _945;
  wire _29215 = _8010 ^ _29214;
  wire _29216 = _20006 ^ _18584;
  wire _29217 = _29215 ^ _29216;
  wire _29218 = _29213 ^ _29217;
  wire _29219 = _14622 ^ _3291;
  wire _29220 = _11405 ^ _98;
  wire _29221 = _29219 ^ _29220;
  wire _29222 = _4785 ^ _4787;
  wire _29223 = _29222 ^ _22844;
  wire _29224 = _29221 ^ _29223;
  wire _29225 = uncoded_block[230] ^ uncoded_block[233];
  wire _29226 = _29225 ^ _7423;
  wire _29227 = _10292 ^ _5505;
  wire _29228 = _29226 ^ _29227;
  wire _29229 = _4800 ^ _117;
  wire _29230 = uncoded_block[261] ^ uncoded_block[266];
  wire _29231 = _29230 ^ _4099;
  wire _29232 = _29229 ^ _29231;
  wire _29233 = _29228 ^ _29232;
  wire _29234 = _29224 ^ _29233;
  wire _29235 = _29218 ^ _29234;
  wire _29236 = _29203 ^ _29235;
  wire _29237 = _19566 ^ _19570;
  wire _29238 = uncoded_block[284] ^ uncoded_block[287];
  wire _29239 = _6194 ^ _29238;
  wire _29240 = _29237 ^ _29239;
  wire _29241 = uncoded_block[299] ^ uncoded_block[306];
  wire _29242 = _29241 ^ _3334;
  wire _29243 = _10313 ^ _29242;
  wire _29244 = _29240 ^ _29243;
  wire _29245 = uncoded_block[318] ^ uncoded_block[323];
  wire _29246 = _29245 ^ _11444;
  wire _29247 = _15672 ^ _29246;
  wire _29248 = _11983 ^ _2587;
  wire _29249 = uncoded_block[337] ^ uncoded_block[342];
  wire _29250 = _29249 ^ _4841;
  wire _29251 = _29248 ^ _29250;
  wire _29252 = _29247 ^ _29251;
  wire _29253 = _29244 ^ _29252;
  wire _29254 = _4845 ^ _19092;
  wire _29255 = _1029 ^ _12530;
  wire _29256 = _29254 ^ _29255;
  wire _29257 = uncoded_block[372] ^ uncoded_block[375];
  wire _29258 = _1838 ^ _29257;
  wire _29259 = _9795 ^ _29258;
  wire _29260 = _29256 ^ _29259;
  wire _29261 = _2612 ^ _11999;
  wire _29262 = _24235 ^ _29261;
  wire _29263 = _19601 ^ _20563;
  wire _29264 = _29262 ^ _29263;
  wire _29265 = _29260 ^ _29264;
  wire _29266 = _29253 ^ _29265;
  wire _29267 = _1048 ^ _183;
  wire _29268 = _12545 ^ _1853;
  wire _29269 = _29267 ^ _29268;
  wire _29270 = _24707 ^ _9816;
  wire _29271 = _1063 ^ _4169;
  wire _29272 = _29270 ^ _29271;
  wire _29273 = _29269 ^ _29272;
  wire _29274 = _2641 ^ _3408;
  wire _29275 = _12559 ^ _17185;
  wire _29276 = _29274 ^ _29275;
  wire _29277 = _26942 ^ _9284;
  wire _29278 = _29276 ^ _29277;
  wire _29279 = _29273 ^ _29278;
  wire _29280 = uncoded_block[471] ^ uncoded_block[476];
  wire _29281 = _29280 ^ _8693;
  wire _29282 = _8694 ^ _7516;
  wire _29283 = _29281 ^ _29282;
  wire _29284 = uncoded_block[493] ^ uncoded_block[497];
  wire _29285 = _3424 ^ _29284;
  wire _29286 = _29285 ^ _3435;
  wire _29287 = _29283 ^ _29286;
  wire _29288 = _1892 ^ _3437;
  wire _29289 = uncoded_block[512] ^ uncoded_block[517];
  wire _29290 = _29289 ^ _19638;
  wire _29291 = _29288 ^ _29290;
  wire _29292 = _237 ^ _20099;
  wire _29293 = _25171 ^ _8718;
  wire _29294 = _29292 ^ _29293;
  wire _29295 = _29291 ^ _29294;
  wire _29296 = _29287 ^ _29295;
  wire _29297 = _29279 ^ _29296;
  wire _29298 = _29266 ^ _29297;
  wire _29299 = _29236 ^ _29298;
  wire _29300 = _1908 ^ _24282;
  wire _29301 = _8720 ^ _6304;
  wire _29302 = _29300 ^ _29301;
  wire _29303 = _1916 ^ _23826;
  wire _29304 = _7550 ^ _8731;
  wire _29305 = _29303 ^ _29304;
  wire _29306 = _29302 ^ _29305;
  wire _29307 = _5641 ^ _26096;
  wire _29308 = uncoded_block[593] ^ uncoded_block[606];
  wire _29309 = _2700 ^ _29308;
  wire _29310 = _29307 ^ _29309;
  wire _29311 = uncoded_block[614] ^ uncoded_block[617];
  wire _29312 = _8739 ^ _29311;
  wire _29313 = uncoded_block[620] ^ uncoded_block[625];
  wire _29314 = _4243 ^ _29313;
  wire _29315 = _29312 ^ _29314;
  wire _29316 = _29310 ^ _29315;
  wire _29317 = _29306 ^ _29316;
  wire _29318 = uncoded_block[626] ^ uncoded_block[629];
  wire _29319 = _29318 ^ _3501;
  wire _29320 = uncoded_block[637] ^ uncoded_block[648];
  wire _29321 = _29320 ^ _14234;
  wire _29322 = _29319 ^ _29321;
  wire _29323 = _1962 ^ _21113;
  wire _29324 = _13190 ^ _8176;
  wire _29325 = _29323 ^ _29324;
  wire _29326 = _29322 ^ _29325;
  wire _29327 = _19191 ^ _10442;
  wire _29328 = _19190 ^ _29327;
  wire _29329 = _2754 ^ _18719;
  wire _29330 = _5685 ^ _4995;
  wire _29331 = _29329 ^ _29330;
  wire _29332 = _29328 ^ _29331;
  wire _29333 = _29326 ^ _29332;
  wire _29334 = _29317 ^ _29333;
  wire _29335 = _1192 ^ _4999;
  wire _29336 = _17762 ^ _21129;
  wire _29337 = _29335 ^ _29336;
  wire _29338 = _7001 ^ _1991;
  wire _29339 = uncoded_block[734] ^ uncoded_block[741];
  wire _29340 = _29339 ^ _21136;
  wire _29341 = _29338 ^ _29340;
  wire _29342 = _29337 ^ _29341;
  wire _29343 = _5013 ^ _2002;
  wire _29344 = _8779 ^ _359;
  wire _29345 = _29343 ^ _29344;
  wire _29346 = _4301 ^ _9381;
  wire _29347 = _18270 ^ _29346;
  wire _29348 = _29345 ^ _29347;
  wire _29349 = _29342 ^ _29348;
  wire _29350 = _1221 ^ _27017;
  wire _29351 = _5715 ^ _4314;
  wire _29352 = _29350 ^ _29351;
  wire _29353 = uncoded_block[796] ^ uncoded_block[807];
  wire _29354 = _29353 ^ _5041;
  wire _29355 = _2806 ^ _1241;
  wire _29356 = _29354 ^ _29355;
  wire _29357 = _29352 ^ _29356;
  wire _29358 = uncoded_block[823] ^ uncoded_block[826];
  wire _29359 = _27843 ^ _29358;
  wire _29360 = _2033 ^ _4336;
  wire _29361 = _29359 ^ _29360;
  wire _29362 = _1257 ^ _6406;
  wire _29363 = _14810 ^ _29362;
  wire _29364 = _29361 ^ _29363;
  wire _29365 = _29357 ^ _29364;
  wire _29366 = _29349 ^ _29365;
  wire _29367 = _29334 ^ _29366;
  wire _29368 = uncoded_block[854] ^ uncoded_block[857];
  wire _29369 = _29368 ^ _11614;
  wire _29370 = _17304 ^ _6416;
  wire _29371 = _29369 ^ _29370;
  wire _29372 = _9954 ^ _11624;
  wire _29373 = _10506 ^ _1277;
  wire _29374 = _29372 ^ _29373;
  wire _29375 = _29371 ^ _29374;
  wire _29376 = _2844 ^ _1281;
  wire _29377 = _17311 ^ _29376;
  wire _29378 = _6428 ^ _18775;
  wire _29379 = uncoded_block[924] ^ uncoded_block[927];
  wire _29380 = _29379 ^ _1296;
  wire _29381 = _29378 ^ _29380;
  wire _29382 = _29377 ^ _29381;
  wire _29383 = _29375 ^ _29382;
  wire _29384 = _3637 ^ _10517;
  wire _29385 = _26628 ^ _2865;
  wire _29386 = _29384 ^ _29385;
  wire _29387 = uncoded_block[947] ^ uncoded_block[950];
  wire _29388 = _29387 ^ _1303;
  wire _29389 = uncoded_block[957] ^ uncoded_block[962];
  wire _29390 = _461 ^ _29389;
  wire _29391 = _29388 ^ _29390;
  wire _29392 = _29386 ^ _29391;
  wire _29393 = _10531 ^ _7088;
  wire _29394 = _468 ^ _3657;
  wire _29395 = _29393 ^ _29394;
  wire _29396 = _10535 ^ _10538;
  wire _29397 = _29395 ^ _29396;
  wire _29398 = _29392 ^ _29397;
  wire _29399 = _29383 ^ _29398;
  wire _29400 = _8856 ^ _479;
  wire _29401 = _29400 ^ _12739;
  wire _29402 = _8866 ^ _2890;
  wire _29403 = uncoded_block[1014] ^ uncoded_block[1019];
  wire _29404 = _29403 ^ _14855;
  wire _29405 = _29402 ^ _29404;
  wire _29406 = _29401 ^ _29405;
  wire _29407 = _9455 ^ _2898;
  wire _29408 = _12198 ^ _511;
  wire _29409 = _29407 ^ _29408;
  wire _29410 = uncoded_block[1045] ^ uncoded_block[1048];
  wire _29411 = _11677 ^ _29410;
  wire _29412 = _518 ^ _12762;
  wire _29413 = _29411 ^ _29412;
  wire _29414 = _29409 ^ _29413;
  wire _29415 = _29406 ^ _29414;
  wire _29416 = _8311 ^ _19298;
  wire _29417 = _29416 ^ _8890;
  wire _29418 = _13851 ^ _5158;
  wire _29419 = _2146 ^ _5163;
  wire _29420 = _29418 ^ _29419;
  wire _29421 = _29417 ^ _29420;
  wire _29422 = uncoded_block[1087] ^ uncoded_block[1094];
  wire _29423 = _11687 ^ _29422;
  wire _29424 = _5846 ^ _8910;
  wire _29425 = _29423 ^ _29424;
  wire _29426 = uncoded_block[1105] ^ uncoded_block[1111];
  wire _29427 = uncoded_block[1117] ^ uncoded_block[1121];
  wire _29428 = _29426 ^ _29427;
  wire _29429 = _12789 ^ _18371;
  wire _29430 = _29428 ^ _29429;
  wire _29431 = _29425 ^ _29430;
  wire _29432 = _29421 ^ _29431;
  wire _29433 = _29415 ^ _29432;
  wire _29434 = _29399 ^ _29433;
  wire _29435 = _29367 ^ _29434;
  wire _29436 = _29299 ^ _29435;
  wire _29437 = _2949 ^ _564;
  wire _29438 = _29437 ^ _21243;
  wire _29439 = uncoded_block[1151] ^ uncoded_block[1154];
  wire _29440 = _29439 ^ _3728;
  wire _29441 = _6506 ^ _29440;
  wire _29442 = _29438 ^ _29441;
  wire _29443 = _578 ^ _22627;
  wire _29444 = uncoded_block[1169] ^ uncoded_block[1173];
  wire _29445 = _15907 ^ _29444;
  wire _29446 = _29443 ^ _29445;
  wire _29447 = _25798 ^ _23537;
  wire _29448 = _29446 ^ _29447;
  wire _29449 = _29442 ^ _29448;
  wire _29450 = _11719 ^ _599;
  wire _29451 = _20283 ^ _29450;
  wire _29452 = uncoded_block[1208] ^ uncoded_block[1216];
  wire _29453 = _29452 ^ _3763;
  wire _29454 = _15433 ^ _29453;
  wire _29455 = _29451 ^ _29454;
  wire _29456 = _12815 ^ _612;
  wire _29457 = _1439 ^ _15926;
  wire _29458 = _29456 ^ _29457;
  wire _29459 = _7174 ^ _6536;
  wire _29460 = _18860 ^ _2997;
  wire _29461 = _29459 ^ _29460;
  wire _29462 = _29458 ^ _29461;
  wire _29463 = _29455 ^ _29462;
  wire _29464 = _29449 ^ _29463;
  wire _29465 = _2998 ^ _22651;
  wire _29466 = _20801 ^ _5235;
  wire _29467 = _29465 ^ _29466;
  wire _29468 = uncoded_block[1276] ^ uncoded_block[1280];
  wire _29469 = _26718 ^ _29468;
  wire _29470 = _29058 ^ _29469;
  wire _29471 = _29467 ^ _29470;
  wire _29472 = uncoded_block[1281] ^ uncoded_block[1284];
  wire _29473 = _29472 ^ _639;
  wire _29474 = _29473 ^ _13381;
  wire _29475 = _3018 ^ _1479;
  wire _29476 = _13917 ^ _1483;
  wire _29477 = _29475 ^ _29476;
  wire _29478 = _29474 ^ _29477;
  wire _29479 = _29471 ^ _29478;
  wire _29480 = _23134 ^ _9555;
  wire _29481 = uncoded_block[1323] ^ uncoded_block[1327];
  wire _29482 = _29481 ^ _8997;
  wire _29483 = _29480 ^ _29482;
  wire _29484 = _14947 ^ _28674;
  wire _29485 = _29483 ^ _29484;
  wire _29486 = uncoded_block[1342] ^ uncoded_block[1345];
  wire _29487 = _29486 ^ _5268;
  wire _29488 = _670 ^ _16942;
  wire _29489 = _29487 ^ _29488;
  wire _29490 = _23581 ^ _15962;
  wire _29491 = _29490 ^ _3053;
  wire _29492 = _29489 ^ _29491;
  wire _29493 = _29485 ^ _29492;
  wire _29494 = _29479 ^ _29493;
  wire _29495 = _29464 ^ _29494;
  wire _29496 = uncoded_block[1375] ^ uncoded_block[1380];
  wire _29497 = _29496 ^ _3059;
  wire _29498 = uncoded_block[1388] ^ uncoded_block[1393];
  wire _29499 = _6596 ^ _29498;
  wire _29500 = _29497 ^ _29499;
  wire _29501 = _2299 ^ _4578;
  wire _29502 = _3067 ^ _29501;
  wire _29503 = _29500 ^ _29502;
  wire _29504 = _2300 ^ _23163;
  wire _29505 = _29504 ^ _8439;
  wire _29506 = _16463 ^ _24058;
  wire _29507 = uncoded_block[1427] ^ uncoded_block[1432];
  wire _29508 = uncoded_block[1436] ^ uncoded_block[1438];
  wire _29509 = _29507 ^ _29508;
  wire _29510 = _29506 ^ _29509;
  wire _29511 = _29505 ^ _29510;
  wire _29512 = _29503 ^ _29511;
  wire _29513 = _1541 ^ _8450;
  wire _29514 = _5976 ^ _720;
  wire _29515 = _29513 ^ _29514;
  wire _29516 = uncoded_block[1457] ^ uncoded_block[1461];
  wire _29517 = uncoded_block[1462] ^ uncoded_block[1467];
  wire _29518 = _29516 ^ _29517;
  wire _29519 = uncoded_block[1468] ^ uncoded_block[1471];
  wire _29520 = _29519 ^ _3097;
  wire _29521 = _29518 ^ _29520;
  wire _29522 = _29515 ^ _29521;
  wire _29523 = _1558 ^ _10706;
  wire _29524 = _21334 ^ _29523;
  wire _29525 = _3887 ^ _23189;
  wire _29526 = _29524 ^ _29525;
  wire _29527 = _29522 ^ _29526;
  wire _29528 = _29512 ^ _29527;
  wire _29529 = uncoded_block[1506] ^ uncoded_block[1513];
  wire _29530 = _4614 ^ _29529;
  wire _29531 = _16004 ^ _7265;
  wire _29532 = _29530 ^ _29531;
  wire _29533 = _15004 ^ _11270;
  wire _29534 = _3122 ^ _5343;
  wire _29535 = _29533 ^ _29534;
  wire _29536 = _29532 ^ _29535;
  wire _29537 = _11820 ^ _19903;
  wire _29538 = uncoded_block[1550] ^ uncoded_block[1558];
  wire _29539 = _4634 ^ _29538;
  wire _29540 = _29537 ^ _29539;
  wire _29541 = _13991 ^ _6019;
  wire _29542 = uncoded_block[1568] ^ uncoded_block[1572];
  wire _29543 = _29542 ^ _4647;
  wire _29544 = _29541 ^ _29543;
  wire _29545 = _29540 ^ _29544;
  wire _29546 = _29536 ^ _29545;
  wire _29547 = _2380 ^ _2383;
  wire _29548 = _6031 ^ _788;
  wire _29549 = _29547 ^ _29548;
  wire _29550 = uncoded_block[1597] ^ uncoded_block[1599];
  wire _29551 = _29550 ^ _1624;
  wire _29552 = _13485 ^ _29551;
  wire _29553 = _29549 ^ _29552;
  wire _29554 = _6677 ^ _5380;
  wire _29555 = _801 ^ _7297;
  wire _29556 = _29554 ^ _29555;
  wire _29557 = uncoded_block[1621] ^ uncoded_block[1626];
  wire _29558 = _29557 ^ _5388;
  wire _29559 = _3946 ^ _14009;
  wire _29560 = _29558 ^ _29559;
  wire _29561 = _29556 ^ _29560;
  wire _29562 = _29553 ^ _29561;
  wire _29563 = _29546 ^ _29562;
  wire _29564 = _29528 ^ _29563;
  wire _29565 = _29495 ^ _29564;
  wire _29566 = _3169 ^ _14530;
  wire _29567 = _18030 ^ _10760;
  wire _29568 = _29566 ^ _29567;
  wire _29569 = uncoded_block[1659] ^ uncoded_block[1661];
  wire _29570 = _29569 ^ _9666;
  wire _29571 = _6059 ^ _832;
  wire _29572 = _29570 ^ _29571;
  wire _29573 = _29568 ^ _29572;
  wire _29574 = _3187 ^ _24130;
  wire _29575 = _20428 ^ _29574;
  wire _29576 = _3968 ^ _9677;
  wire _29577 = _20436 ^ _3979;
  wire _29578 = _29576 ^ _29577;
  wire _29579 = _29575 ^ _29578;
  wire _29580 = _29573 ^ _29579;
  wire _29581 = _7337 ^ _3200;
  wire _29582 = _29581 ^ _10217;
  wire _29583 = _29580 ^ _29582;
  wire _29584 = _29565 ^ _29583;
  wire _29585 = _29436 ^ _29584;
  wire _29586 = _3210 ^ _24147;
  wire _29587 = _3995 ^ _7;
  wire _29588 = _29586 ^ _29587;
  wire _29589 = uncoded_block[13] ^ uncoded_block[20];
  wire _29590 = _29589 ^ _3219;
  wire _29591 = _5427 ^ _16;
  wire _29592 = _29590 ^ _29591;
  wire _29593 = _29588 ^ _29592;
  wire _29594 = _2466 ^ _22;
  wire _29595 = _22795 ^ _13547;
  wire _29596 = _29594 ^ _29595;
  wire _29597 = _16572 ^ _7364;
  wire _29598 = _32 ^ _25950;
  wire _29599 = _29597 ^ _29598;
  wire _29600 = _29596 ^ _29599;
  wire _29601 = _29593 ^ _29600;
  wire _29602 = _7976 ^ _19511;
  wire _29603 = _3243 ^ _28438;
  wire _29604 = _29602 ^ _29603;
  wire _29605 = _4025 ^ _15603;
  wire _29606 = _29605 ^ _19024;
  wire _29607 = _29604 ^ _29606;
  wire _29608 = _47 ^ _4745;
  wire _29609 = _4031 ^ _6123;
  wire _29610 = _29608 ^ _29609;
  wire _29611 = uncoded_block[119] ^ uncoded_block[123];
  wire _29612 = _6126 ^ _29611;
  wire _29613 = _29612 ^ _10258;
  wire _29614 = _29610 ^ _29613;
  wire _29615 = _29607 ^ _29614;
  wire _29616 = _29601 ^ _29615;
  wire _29617 = _9177 ^ _4760;
  wire _29618 = _11924 ^ _6780;
  wire _29619 = _29617 ^ _29618;
  wire _29620 = _1744 ^ _15623;
  wire _29621 = _29620 ^ _7398;
  wire _29622 = _29619 ^ _29621;
  wire _29623 = uncoded_block[158] ^ uncoded_block[165];
  wire _29624 = uncoded_block[166] ^ uncoded_block[168];
  wire _29625 = _29623 ^ _29624;
  wire _29626 = _2521 ^ _1756;
  wire _29627 = _29625 ^ _29626;
  wire _29628 = uncoded_block[184] ^ uncoded_block[189];
  wire _29629 = _941 ^ _29628;
  wire _29630 = _5483 ^ _1763;
  wire _29631 = _29629 ^ _29630;
  wire _29632 = _29627 ^ _29631;
  wire _29633 = _29622 ^ _29632;
  wire _29634 = uncoded_block[203] ^ uncoded_block[206];
  wire _29635 = _22837 ^ _29634;
  wire _29636 = _8600 ^ _4071;
  wire _29637 = _29635 ^ _29636;
  wire _29638 = _9202 ^ _14105;
  wire _29639 = _4076 ^ _11410;
  wire _29640 = _29638 ^ _29639;
  wire _29641 = _29637 ^ _29640;
  wire _29642 = uncoded_block[232] ^ uncoded_block[237];
  wire _29643 = _29642 ^ _5500;
  wire _29644 = uncoded_block[241] ^ uncoded_block[247];
  wire _29645 = uncoded_block[248] ^ uncoded_block[255];
  wire _29646 = _29644 ^ _29645;
  wire _29647 = _29643 ^ _29646;
  wire _29648 = _26000 ^ _14642;
  wire _29649 = _16630 ^ _29648;
  wire _29650 = _29647 ^ _29649;
  wire _29651 = _29641 ^ _29650;
  wire _29652 = _29633 ^ _29651;
  wire _29653 = _29616 ^ _29652;
  wire _29654 = _130 ^ _5513;
  wire _29655 = _29654 ^ _11425;
  wire _29656 = uncoded_block[299] ^ uncoded_block[302];
  wire _29657 = _1806 ^ _29656;
  wire _29658 = _19575 ^ _29657;
  wire _29659 = _29655 ^ _29658;
  wire _29660 = _8052 ^ _15668;
  wire _29661 = _13619 ^ _1006;
  wire _29662 = _29660 ^ _29661;
  wire _29663 = uncoded_block[318] ^ uncoded_block[322];
  wire _29664 = _29663 ^ _8642;
  wire _29665 = _4125 ^ _3352;
  wire _29666 = _29664 ^ _29665;
  wire _29667 = _29662 ^ _29666;
  wire _29668 = _29659 ^ _29667;
  wire _29669 = _8646 ^ _1825;
  wire _29670 = uncoded_block[346] ^ uncoded_block[354];
  wire _29671 = _1826 ^ _29670;
  wire _29672 = _29669 ^ _29671;
  wire _29673 = _6221 ^ _6866;
  wire _29674 = _9250 ^ _17163;
  wire _29675 = _29673 ^ _29674;
  wire _29676 = _29672 ^ _29675;
  wire _29677 = _4853 ^ _6233;
  wire _29678 = _20558 ^ _29677;
  wire _29679 = _7476 ^ _6876;
  wire _29680 = _11999 ^ _2615;
  wire _29681 = _29679 ^ _29680;
  wire _29682 = _29678 ^ _29681;
  wire _29683 = _29676 ^ _29682;
  wire _29684 = _29668 ^ _29683;
  wire _29685 = _3383 ^ _26042;
  wire _29686 = uncoded_block[400] ^ uncoded_block[405];
  wire _29687 = _29686 ^ _184;
  wire _29688 = _29685 ^ _29687;
  wire _29689 = _8091 ^ _7492;
  wire _29690 = _29689 ^ _9817;
  wire _29691 = _29688 ^ _29690;
  wire _29692 = _15704 ^ _2640;
  wire _29693 = _14690 ^ _21049;
  wire _29694 = _29692 ^ _29693;
  wire _29695 = uncoded_block[443] ^ uncoded_block[447];
  wire _29696 = _29695 ^ _4176;
  wire _29697 = _209 ^ _3415;
  wire _29698 = _29696 ^ _29697;
  wire _29699 = _29694 ^ _29698;
  wire _29700 = _29691 ^ _29699;
  wire _29701 = _5586 ^ _23357;
  wire _29702 = uncoded_block[473] ^ uncoded_block[476];
  wire _29703 = _29702 ^ _1085;
  wire _29704 = _29701 ^ _29703;
  wire _29705 = _4902 ^ _1093;
  wire _29706 = _10369 ^ _29705;
  wire _29707 = _29704 ^ _29706;
  wire _29708 = uncoded_block[496] ^ uncoded_block[500];
  wire _29709 = _29708 ^ _19135;
  wire _29710 = _1887 ^ _6283;
  wire _29711 = _29709 ^ _29710;
  wire _29712 = _9295 ^ _23370;
  wire _29713 = _19638 ^ _20097;
  wire _29714 = _29712 ^ _29713;
  wire _29715 = _29711 ^ _29714;
  wire _29716 = _29707 ^ _29715;
  wire _29717 = _29700 ^ _29716;
  wire _29718 = _29684 ^ _29717;
  wire _29719 = _29653 ^ _29718;
  wire _29720 = _1114 ^ _3451;
  wire _29721 = _27782 ^ _6300;
  wire _29722 = _29720 ^ _29721;
  wire _29723 = _1916 ^ _4938;
  wire _29724 = _13160 ^ _29723;
  wire _29725 = _29722 ^ _29724;
  wire _29726 = uncoded_block[562] ^ uncoded_block[568];
  wire _29727 = _29726 ^ _3472;
  wire _29728 = _29727 ^ _10968;
  wire _29729 = _22012 ^ _270;
  wire _29730 = _273 ^ _1941;
  wire _29731 = _29729 ^ _29730;
  wire _29732 = _29728 ^ _29731;
  wire _29733 = _29725 ^ _29732;
  wire _29734 = _14218 ^ _6323;
  wire _29735 = _17232 ^ _29311;
  wire _29736 = _29734 ^ _29735;
  wire _29737 = _7568 ^ _20126;
  wire _29738 = _1953 ^ _3501;
  wire _29739 = _29737 ^ _29738;
  wire _29740 = _29736 ^ _29739;
  wire _29741 = uncoded_block[636] ^ uncoded_block[642];
  wire _29742 = _29741 ^ _4972;
  wire _29743 = uncoded_block[645] ^ uncoded_block[648];
  wire _29744 = _29743 ^ _301;
  wire _29745 = _29742 ^ _29744;
  wire _29746 = _6974 ^ _14755;
  wire _29747 = _18705 ^ _13726;
  wire _29748 = _29746 ^ _29747;
  wire _29749 = _29745 ^ _29748;
  wire _29750 = _29740 ^ _29749;
  wire _29751 = _29733 ^ _29750;
  wire _29752 = _7586 ^ _1178;
  wire _29753 = _10434 ^ _10440;
  wire _29754 = _29752 ^ _29753;
  wire _29755 = _18249 ^ _13735;
  wire _29756 = uncoded_block[693] ^ uncoded_block[696];
  wire _29757 = _29756 ^ _4990;
  wire _29758 = _29755 ^ _29757;
  wire _29759 = _29754 ^ _29758;
  wire _29760 = _3533 ^ _19688;
  wire _29761 = uncoded_block[712] ^ uncoded_block[716];
  wire _29762 = _29761 ^ _17762;
  wire _29763 = _29760 ^ _29762;
  wire _29764 = _9369 ^ _1988;
  wire _29765 = uncoded_block[727] ^ uncoded_block[732];
  wire _29766 = _29765 ^ _5006;
  wire _29767 = _29764 ^ _29766;
  wire _29768 = _29763 ^ _29767;
  wire _29769 = _29759 ^ _29768;
  wire _29770 = _23425 ^ _23870;
  wire _29771 = _29770 ^ _12656;
  wire _29772 = _2775 ^ _24331;
  wire _29773 = _2778 ^ _4298;
  wire _29774 = _29772 ^ _29773;
  wire _29775 = _29771 ^ _29774;
  wire _29776 = _4299 ^ _2783;
  wire _29777 = _5709 ^ _7617;
  wire _29778 = _29776 ^ _29777;
  wire _29779 = _20165 ^ _5715;
  wire _29780 = _8790 ^ _374;
  wire _29781 = _29779 ^ _29780;
  wire _29782 = _29778 ^ _29781;
  wire _29783 = _29775 ^ _29782;
  wire _29784 = _29769 ^ _29783;
  wire _29785 = _29751 ^ _29784;
  wire _29786 = _11591 ^ _2801;
  wire _29787 = _29786 ^ _25240;
  wire _29788 = uncoded_block[817] ^ uncoded_block[820];
  wire _29789 = _2808 ^ _29788;
  wire _29790 = _25702 ^ _29789;
  wire _29791 = _29787 ^ _29790;
  wire _29792 = _7037 ^ _29358;
  wire _29793 = _2812 ^ _12686;
  wire _29794 = _29792 ^ _29793;
  wire _29795 = _13783 ^ _3599;
  wire _29796 = _12689 ^ _29795;
  wire _29797 = _29794 ^ _29796;
  wire _29798 = _29791 ^ _29797;
  wire _29799 = _12146 ^ _2823;
  wire _29800 = uncoded_block[862] ^ uncoded_block[865];
  wire _29801 = _29800 ^ _12150;
  wire _29802 = _29799 ^ _29801;
  wire _29803 = uncoded_block[878] ^ uncoded_block[881];
  wire _29804 = _15826 ^ _29803;
  wire _29805 = _29804 ^ _20197;
  wire _29806 = _29802 ^ _29805;
  wire _29807 = _1273 ^ _14827;
  wire _29808 = uncoded_block[894] ^ uncoded_block[899];
  wire _29809 = uncoded_block[900] ^ uncoded_block[903];
  wire _29810 = _29808 ^ _29809;
  wire _29811 = _29807 ^ _29810;
  wire _29812 = _8254 ^ _6428;
  wire _29813 = _12708 ^ _5092;
  wire _29814 = _29812 ^ _29813;
  wire _29815 = _29811 ^ _29814;
  wire _29816 = _29806 ^ _29815;
  wire _29817 = _29798 ^ _29816;
  wire _29818 = _15350 ^ _439;
  wire _29819 = _445 ^ _8834;
  wire _29820 = _29818 ^ _29819;
  wire _29821 = _1296 ^ _24837;
  wire _29822 = _6439 ^ _24840;
  wire _29823 = _29821 ^ _29822;
  wire _29824 = _29820 ^ _29823;
  wire _29825 = _4384 ^ _464;
  wire _29826 = _4383 ^ _29825;
  wire _29827 = _11646 ^ _2093;
  wire _29828 = _7088 ^ _19268;
  wire _29829 = _29827 ^ _29828;
  wire _29830 = _29826 ^ _29829;
  wire _29831 = _29824 ^ _29830;
  wire _29832 = uncoded_block[980] ^ uncoded_block[983];
  wire _29833 = _5114 ^ _29832;
  wire _29834 = _29833 ^ _18331;
  wire _29835 = uncoded_block[991] ^ uncoded_block[996];
  wire _29836 = _16338 ^ _29835;
  wire _29837 = _22584 ^ _483;
  wire _29838 = _29836 ^ _29837;
  wire _29839 = _29834 ^ _29838;
  wire _29840 = _24400 ^ _487;
  wire _29841 = uncoded_block[1012] ^ uncoded_block[1021];
  wire _29842 = _29841 ^ _19766;
  wire _29843 = _29840 ^ _29842;
  wire _29844 = uncoded_block[1030] ^ uncoded_block[1036];
  wire _29845 = _1339 ^ _29844;
  wire _29846 = uncoded_block[1039] ^ uncoded_block[1043];
  wire _29847 = _29846 ^ _8309;
  wire _29848 = _29845 ^ _29847;
  wire _29849 = _29843 ^ _29848;
  wire _29850 = _29839 ^ _29849;
  wire _29851 = _29831 ^ _29850;
  wire _29852 = _29817 ^ _29851;
  wire _29853 = _29785 ^ _29852;
  wire _29854 = _29719 ^ _29853;
  wire _29855 = _5148 ^ _4432;
  wire _29856 = _9475 ^ _527;
  wire _29857 = _23502 ^ _29856;
  wire _29858 = _29855 ^ _29857;
  wire _29859 = uncoded_block[1076] ^ uncoded_block[1079];
  wire _29860 = _8893 ^ _29859;
  wire _29861 = _5163 ^ _15401;
  wire _29862 = _29860 ^ _29861;
  wire _29863 = _1374 ^ _22610;
  wire _29864 = uncoded_block[1096] ^ uncoded_block[1102];
  wire _29865 = _3698 ^ _29864;
  wire _29866 = _29863 ^ _29865;
  wire _29867 = _29862 ^ _29866;
  wire _29868 = _29858 ^ _29867;
  wire _29869 = _25323 ^ _1388;
  wire _29870 = _23976 ^ _29869;
  wire _29871 = uncoded_block[1125] ^ uncoded_block[1131];
  wire _29872 = _5176 ^ _29871;
  wire _29873 = uncoded_block[1132] ^ uncoded_block[1139];
  wire _29874 = _29873 ^ _7743;
  wire _29875 = _29872 ^ _29874;
  wire _29876 = _29870 ^ _29875;
  wire _29877 = _4465 ^ _8933;
  wire _29878 = uncoded_block[1156] ^ uncoded_block[1158];
  wire _29879 = _3727 ^ _29878;
  wire _29880 = _29877 ^ _29879;
  wire _29881 = _7149 ^ _3736;
  wire _29882 = _1408 ^ _3739;
  wire _29883 = _29881 ^ _29882;
  wire _29884 = _29880 ^ _29883;
  wire _29885 = _29876 ^ _29884;
  wire _29886 = _29868 ^ _29885;
  wire _29887 = uncoded_block[1178] ^ uncoded_block[1183];
  wire _29888 = _585 ^ _29887;
  wire _29889 = _23097 ^ _4488;
  wire _29890 = _29888 ^ _29889;
  wire _29891 = _11721 ^ _8370;
  wire _29892 = _2978 ^ _6530;
  wire _29893 = _29891 ^ _29892;
  wire _29894 = _29890 ^ _29893;
  wire _29895 = _2217 ^ _2219;
  wire _29896 = _12815 ^ _2986;
  wire _29897 = _29895 ^ _29896;
  wire _29898 = _14919 ^ _5219;
  wire _29899 = uncoded_block[1236] ^ uncoded_block[1242];
  wire _29900 = _29899 ^ _19829;
  wire _29901 = _29898 ^ _29900;
  wire _29902 = _29897 ^ _29901;
  wire _29903 = _29894 ^ _29902;
  wire _29904 = uncoded_block[1250] ^ uncoded_block[1256];
  wire _29905 = _1451 ^ _29904;
  wire _29906 = uncoded_block[1263] ^ uncoded_block[1266];
  wire _29907 = _5234 ^ _29906;
  wire _29908 = _29905 ^ _29907;
  wire _29909 = _3008 ^ _9538;
  wire _29910 = _29909 ^ _23563;
  wire _29911 = _29908 ^ _29910;
  wire _29912 = uncoded_block[1283] ^ uncoded_block[1288];
  wire _29913 = uncoded_block[1289] ^ uncoded_block[1295];
  wire _29914 = _29912 ^ _29913;
  wire _29915 = _7184 ^ _29914;
  wire _29916 = _645 ^ _16424;
  wire _29917 = _29916 ^ _25833;
  wire _29918 = _29915 ^ _29917;
  wire _29919 = _29911 ^ _29918;
  wire _29920 = _29903 ^ _29919;
  wire _29921 = _29886 ^ _29920;
  wire _29922 = _14430 ^ _5253;
  wire _29923 = _9555 ^ _4543;
  wire _29924 = _29922 ^ _29923;
  wire _29925 = _7201 ^ _8997;
  wire _29926 = _24036 ^ _2277;
  wire _29927 = _29925 ^ _29926;
  wire _29928 = _29924 ^ _29927;
  wire _29929 = _14950 ^ _664;
  wire _29930 = uncoded_block[1351] ^ uncoded_block[1357];
  wire _29931 = _29930 ^ _6588;
  wire _29932 = _29929 ^ _29931;
  wire _29933 = _5275 ^ _10665;
  wire _29934 = uncoded_block[1367] ^ uncoded_block[1370];
  wire _29935 = _29934 ^ _8423;
  wire _29936 = _29933 ^ _29935;
  wire _29937 = _29932 ^ _29936;
  wire _29938 = _29928 ^ _29937;
  wire _29939 = uncoded_block[1378] ^ uncoded_block[1382];
  wire _29940 = _5284 ^ _29939;
  wire _29941 = _29940 ^ _16454;
  wire _29942 = _13412 ^ _694;
  wire _29943 = _2296 ^ _5293;
  wire _29944 = _29942 ^ _29943;
  wire _29945 = _29941 ^ _29944;
  wire _29946 = _4578 ^ _2300;
  wire _29947 = _8436 ^ _17461;
  wire _29948 = _29946 ^ _29947;
  wire _29949 = _27167 ^ _14975;
  wire _29950 = _29948 ^ _29949;
  wire _29951 = _29945 ^ _29950;
  wire _29952 = _29938 ^ _29951;
  wire _29953 = _14466 ^ _5968;
  wire _29954 = _1533 ^ _21324;
  wire _29955 = _29953 ^ _29954;
  wire _29956 = _716 ^ _2322;
  wire _29957 = _719 ^ _5309;
  wire _29958 = _29956 ^ _29957;
  wire _29959 = _29955 ^ _29958;
  wire _29960 = _723 ^ _3870;
  wire _29961 = _2336 ^ _18469;
  wire _29962 = _29960 ^ _29961;
  wire _29963 = _25423 ^ _23181;
  wire _29964 = _10706 ^ _740;
  wire _29965 = _29963 ^ _29964;
  wire _29966 = _29962 ^ _29965;
  wire _29967 = _29959 ^ _29966;
  wire _29968 = _3108 ^ _11260;
  wire _29969 = _1572 ^ _7262;
  wire _29970 = _29968 ^ _29969;
  wire _29971 = _5334 ^ _5336;
  wire _29972 = _29971 ^ _10150;
  wire _29973 = _29970 ^ _29972;
  wire _29974 = _20874 ^ _13979;
  wire _29975 = _20386 ^ _7274;
  wire _29976 = _29974 ^ _29975;
  wire _29977 = uncoded_block[1547] ^ uncoded_block[1553];
  wire _29978 = _29977 ^ _3131;
  wire _29979 = _6016 ^ _3139;
  wire _29980 = _29978 ^ _29979;
  wire _29981 = _29976 ^ _29980;
  wire _29982 = _29973 ^ _29981;
  wire _29983 = _29967 ^ _29982;
  wire _29984 = _29952 ^ _29983;
  wire _29985 = _29921 ^ _29984;
  wire _29986 = uncoded_block[1565] ^ uncoded_block[1568];
  wire _29987 = uncoded_block[1569] ^ uncoded_block[1571];
  wire _29988 = _29986 ^ _29987;
  wire _29989 = _29988 ^ _17008;
  wire _29990 = _6663 ^ _1612;
  wire _29991 = _1615 ^ _3146;
  wire _29992 = _29990 ^ _29991;
  wire _29993 = _29989 ^ _29992;
  wire _29994 = _2394 ^ _6674;
  wire _29995 = _12937 ^ _3153;
  wire _29996 = _29994 ^ _29995;
  wire _29997 = uncoded_block[1614] ^ uncoded_block[1617];
  wire _29998 = _3937 ^ _29997;
  wire _29999 = uncoded_block[1618] ^ uncoded_block[1622];
  wire _30000 = uncoded_block[1626] ^ uncoded_block[1632];
  wire _30001 = _29999 ^ _30000;
  wire _30002 = _29998 ^ _30001;
  wire _30003 = _29996 ^ _30002;
  wire _30004 = _29993 ^ _30003;
  wire _30005 = _3946 ^ _12949;
  wire _30006 = _27651 ^ _18516;
  wire _30007 = _30005 ^ _30006;
  wire _30008 = uncoded_block[1653] ^ uncoded_block[1657];
  wire _30009 = _30008 ^ _1653;
  wire _30010 = _28408 ^ _30009;
  wire _30011 = _30007 ^ _30010;
  wire _30012 = _19470 ^ _3182;
  wire _30013 = _22762 ^ _30012;
  wire _30014 = uncoded_block[1672] ^ uncoded_block[1674];
  wire _30015 = _30014 ^ _3183;
  wire _30016 = _17538 ^ _3965;
  wire _30017 = _30015 ^ _30016;
  wire _30018 = _30013 ^ _30017;
  wire _30019 = _30011 ^ _30018;
  wire _30020 = _30004 ^ _30019;
  wire _30021 = _13519 ^ _6707;
  wire _30022 = _6066 ^ _1669;
  wire _30023 = _30021 ^ _30022;
  wire _30024 = _3975 ^ _847;
  wire _30025 = _30024 ^ _3198;
  wire _30026 = _30023 ^ _30025;
  wire _30027 = uncoded_block[1713] ^ uncoded_block[1715];
  wire _30028 = _30027 ^ _13528;
  wire _30029 = _30028 ^ uncoded_block[1720];
  wire _30030 = _30026 ^ _30029;
  wire _30031 = _30020 ^ _30030;
  wire _30032 = _29985 ^ _30031;
  wire _30033 = _29854 ^ _30032;
  wire _30034 = uncoded_block[7] ^ uncoded_block[11];
  wire _30035 = _21861 ^ _30034;
  wire _30036 = uncoded_block[18] ^ uncoded_block[21];
  wire _30037 = _7956 ^ _30036;
  wire _30038 = _30035 ^ _30037;
  wire _30039 = uncoded_block[28] ^ uncoded_block[32];
  wire _30040 = _30039 ^ _18;
  wire _30041 = _4002 ^ _30040;
  wire _30042 = _30038 ^ _30041;
  wire _30043 = _19 ^ _15591;
  wire _30044 = _30043 ^ _28005;
  wire _30045 = uncoded_block[56] ^ uncoded_block[64];
  wire _30046 = _30045 ^ _34;
  wire _30047 = _21878 ^ _30046;
  wire _30048 = _30044 ^ _30047;
  wire _30049 = _30042 ^ _30048;
  wire _30050 = _896 ^ _14583;
  wire _30051 = uncoded_block[79] ^ uncoded_block[84];
  wire _30052 = _901 ^ _30051;
  wire _30053 = _30050 ^ _30052;
  wire _30054 = _2487 ^ _6115;
  wire _30055 = _11909 ^ _19025;
  wire _30056 = _30054 ^ _30055;
  wire _30057 = _30053 ^ _30056;
  wire _30058 = _16589 ^ _6128;
  wire _30059 = _11914 ^ _30058;
  wire _30060 = _12451 ^ _20961;
  wire _30061 = _57 ^ _3263;
  wire _30062 = _30060 ^ _30061;
  wire _30063 = _30059 ^ _30062;
  wire _30064 = _30057 ^ _30063;
  wire _30065 = _30049 ^ _30064;
  wire _30066 = _927 ^ _5461;
  wire _30067 = _2511 ^ _67;
  wire _30068 = _30066 ^ _30067;
  wire _30069 = _4048 ^ _9188;
  wire _30070 = _29620 ^ _30069;
  wire _30071 = _30068 ^ _30070;
  wire _30072 = _16108 ^ _13029;
  wire _30073 = _938 ^ _13032;
  wire _30074 = _1757 ^ _4062;
  wire _30075 = _30073 ^ _30074;
  wire _30076 = _30072 ^ _30075;
  wire _30077 = _30071 ^ _30076;
  wire _30078 = uncoded_block[190] ^ uncoded_block[193];
  wire _30079 = _30078 ^ _7411;
  wire _30080 = _16116 ^ _6805;
  wire _30081 = _30079 ^ _30080;
  wire _30082 = uncoded_block[207] ^ uncoded_block[212];
  wire _30083 = _30082 ^ _1767;
  wire _30084 = _15639 ^ _30083;
  wire _30085 = _30081 ^ _30084;
  wire _30086 = _8606 ^ _10854;
  wire _30087 = uncoded_block[231] ^ uncoded_block[234];
  wire _30088 = _10287 ^ _30087;
  wire _30089 = _30086 ^ _30088;
  wire _30090 = _10289 ^ _970;
  wire _30091 = _10860 ^ _11952;
  wire _30092 = _30090 ^ _30091;
  wire _30093 = _30089 ^ _30092;
  wire _30094 = _30085 ^ _30093;
  wire _30095 = _30077 ^ _30094;
  wire _30096 = _30065 ^ _30095;
  wire _30097 = _7432 ^ _3309;
  wire _30098 = _3311 ^ _13055;
  wire _30099 = _30097 ^ _30098;
  wire _30100 = uncoded_block[260] ^ uncoded_block[268];
  wire _30101 = _30100 ^ _2566;
  wire _30102 = _30101 ^ _10873;
  wire _30103 = _30099 ^ _30102;
  wire _30104 = uncoded_block[280] ^ uncoded_block[284];
  wire _30105 = _4814 ^ _30104;
  wire _30106 = uncoded_block[286] ^ uncoded_block[291];
  wire _30107 = _30106 ^ _4819;
  wire _30108 = _30105 ^ _30107;
  wire _30109 = uncoded_block[300] ^ uncoded_block[306];
  wire _30110 = _4110 ^ _30109;
  wire _30111 = uncoded_block[310] ^ uncoded_block[314];
  wire _30112 = _3334 ^ _30111;
  wire _30113 = _30110 ^ _30112;
  wire _30114 = _30108 ^ _30113;
  wire _30115 = _30103 ^ _30114;
  wire _30116 = uncoded_block[319] ^ uncoded_block[322];
  wire _30117 = uncoded_block[326] ^ uncoded_block[328];
  wire _30118 = _30116 ^ _30117;
  wire _30119 = _4831 ^ _30118;
  wire _30120 = _8065 ^ _4129;
  wire _30121 = _17153 ^ _30120;
  wire _30122 = _30119 ^ _30121;
  wire _30123 = uncoded_block[349] ^ uncoded_block[353];
  wire _30124 = _18621 ^ _30123;
  wire _30125 = _8069 ^ _8073;
  wire _30126 = _30124 ^ _30125;
  wire _30127 = _3366 ^ _7470;
  wire _30128 = _8076 ^ _13094;
  wire _30129 = _30127 ^ _30128;
  wire _30130 = _30126 ^ _30129;
  wire _30131 = _30122 ^ _30130;
  wire _30132 = _30115 ^ _30131;
  wire _30133 = _6233 ^ _4857;
  wire _30134 = _30133 ^ _4150;
  wire _30135 = uncoded_block[391] ^ uncoded_block[398];
  wire _30136 = _6239 ^ _30135;
  wire _30137 = _181 ^ _183;
  wire _30138 = _30136 ^ _30137;
  wire _30139 = _30134 ^ _30138;
  wire _30140 = _12545 ^ _24243;
  wire _30141 = _19612 ^ _3396;
  wire _30142 = _30140 ^ _30141;
  wire _30143 = _4163 ^ _2633;
  wire _30144 = _2637 ^ _4167;
  wire _30145 = _30143 ^ _30144;
  wire _30146 = _30142 ^ _30145;
  wire _30147 = _30139 ^ _30146;
  wire _30148 = _6255 ^ _16187;
  wire _30149 = _28852 ^ _30148;
  wire _30150 = _5579 ^ _26056;
  wire _30151 = _30149 ^ _30150;
  wire _30152 = uncoded_block[455] ^ uncoded_block[459];
  wire _30153 = _30152 ^ _2653;
  wire _30154 = _13661 ^ _30153;
  wire _30155 = uncoded_block[463] ^ uncoded_block[466];
  wire _30156 = _30155 ^ _9283;
  wire _30157 = _8686 ^ _4189;
  wire _30158 = _30156 ^ _30157;
  wire _30159 = _30154 ^ _30158;
  wire _30160 = _30151 ^ _30159;
  wire _30161 = _30147 ^ _30160;
  wire _30162 = _30132 ^ _30161;
  wire _30163 = _30096 ^ _30162;
  wire _30164 = _1085 ^ _3423;
  wire _30165 = _7516 ^ _4902;
  wire _30166 = _30164 ^ _30165;
  wire _30167 = uncoded_block[494] ^ uncoded_block[498];
  wire _30168 = _30167 ^ _228;
  wire _30169 = _30168 ^ _23810;
  wire _30170 = _30166 ^ _30169;
  wire _30171 = uncoded_block[515] ^ uncoded_block[522];
  wire _30172 = _17694 ^ _30171;
  wire _30173 = _4921 ^ _16711;
  wire _30174 = _30172 ^ _30173;
  wire _30175 = _16215 ^ _24279;
  wire _30176 = _14198 ^ _2684;
  wire _30177 = _30175 ^ _30176;
  wire _30178 = _30174 ^ _30177;
  wire _30179 = _30170 ^ _30178;
  wire _30180 = _3459 ^ _8724;
  wire _30181 = _30180 ^ _26523;
  wire _30182 = uncoded_block[568] ^ uncoded_block[575];
  wire _30183 = _20110 ^ _30182;
  wire _30184 = _30183 ^ _1134;
  wire _30185 = _30181 ^ _30184;
  wire _30186 = _4947 ^ _18222;
  wire _30187 = uncoded_block[597] ^ uncoded_block[602];
  wire _30188 = _15247 ^ _30187;
  wire _30189 = _30186 ^ _30188;
  wire _30190 = _3489 ^ _2713;
  wire _30191 = _7563 ^ _3494;
  wire _30192 = _30190 ^ _30191;
  wire _30193 = _30189 ^ _30192;
  wire _30194 = _30185 ^ _30193;
  wire _30195 = _30179 ^ _30194;
  wire _30196 = _4963 ^ _10418;
  wire _30197 = _287 ^ _12071;
  wire _30198 = _30196 ^ _30197;
  wire _30199 = uncoded_block[631] ^ uncoded_block[634];
  wire _30200 = _30199 ^ _11543;
  wire _30201 = _9343 ^ _3505;
  wire _30202 = _30200 ^ _30201;
  wire _30203 = _30198 ^ _30202;
  wire _30204 = _301 ^ _2738;
  wire _30205 = _4261 ^ _15768;
  wire _30206 = _30204 ^ _30205;
  wire _30207 = _10990 ^ _10434;
  wire _30208 = _8179 ^ _4271;
  wire _30209 = _30207 ^ _30208;
  wire _30210 = _30206 ^ _30209;
  wire _30211 = _30203 ^ _30210;
  wire _30212 = uncoded_block[692] ^ uncoded_block[696];
  wire _30213 = _6357 ^ _30212;
  wire _30214 = uncoded_block[697] ^ uncoded_block[701];
  wire _30215 = _30214 ^ _18721;
  wire _30216 = _30213 ^ _30215;
  wire _30217 = _3533 ^ _10448;
  wire _30218 = _10452 ^ _1195;
  wire _30219 = _30217 ^ _30218;
  wire _30220 = _30216 ^ _30219;
  wire _30221 = uncoded_block[720] ^ uncoded_block[722];
  wire _30222 = _30221 ^ _344;
  wire _30223 = _7603 ^ _7002;
  wire _30224 = _30222 ^ _30223;
  wire _30225 = _7605 ^ _1207;
  wire _30226 = _1998 ^ _12107;
  wire _30227 = _30225 ^ _30226;
  wire _30228 = _30224 ^ _30227;
  wire _30229 = _30220 ^ _30228;
  wire _30230 = _30211 ^ _30229;
  wire _30231 = _30195 ^ _30230;
  wire _30232 = uncoded_block[753] ^ uncoded_block[756];
  wire _30233 = _30232 ^ _8781;
  wire _30234 = uncoded_block[767] ^ uncoded_block[772];
  wire _30235 = _4301 ^ _30234;
  wire _30236 = _30233 ^ _30235;
  wire _30237 = _2012 ^ _2014;
  wire _30238 = uncoded_block[781] ^ uncoded_block[787];
  wire _30239 = _368 ^ _30238;
  wire _30240 = _30237 ^ _30239;
  wire _30241 = _30236 ^ _30240;
  wire _30242 = _5033 ^ _14282;
  wire _30243 = _7628 ^ _5039;
  wire _30244 = _30242 ^ _30243;
  wire _30245 = _3581 ^ _2806;
  wire _30246 = _7634 ^ _5051;
  wire _30247 = _30245 ^ _30246;
  wire _30248 = _30244 ^ _30247;
  wire _30249 = _30241 ^ _30248;
  wire _30250 = _4328 ^ _5734;
  wire _30251 = _1250 ^ _11607;
  wire _30252 = _30250 ^ _30251;
  wire _30253 = _2036 ^ _14812;
  wire _30254 = _3599 ^ _14814;
  wire _30255 = _30253 ^ _30254;
  wire _30256 = _30252 ^ _30255;
  wire _30257 = _2821 ^ _3600;
  wire _30258 = _5747 ^ _9948;
  wire _30259 = _30257 ^ _30258;
  wire _30260 = uncoded_block[868] ^ uncoded_block[872];
  wire _30261 = _30260 ^ _3608;
  wire _30262 = _22087 ^ _30261;
  wire _30263 = _30259 ^ _30262;
  wire _30264 = _30256 ^ _30263;
  wire _30265 = _30249 ^ _30264;
  wire _30266 = _29803 ^ _423;
  wire _30267 = uncoded_block[888] ^ uncoded_block[896];
  wire _30268 = _11059 ^ _30267;
  wire _30269 = _30266 ^ _30268;
  wire _30270 = uncoded_block[908] ^ uncoded_block[911];
  wire _30271 = _5089 ^ _30270;
  wire _30272 = uncoded_block[912] ^ uncoded_block[918];
  wire _30273 = _30272 ^ _439;
  wire _30274 = _30271 ^ _30273;
  wire _30275 = _30269 ^ _30274;
  wire _30276 = uncoded_block[923] ^ uncoded_block[926];
  wire _30277 = _30276 ^ _446;
  wire _30278 = _5773 ^ _24837;
  wire _30279 = _30277 ^ _30278;
  wire _30280 = _12171 ^ _2086;
  wire _30281 = _30280 ^ _21192;
  wire _30282 = _30279 ^ _30281;
  wire _30283 = _30275 ^ _30282;
  wire _30284 = _4384 ^ _7680;
  wire _30285 = _30284 ^ _27063;
  wire _30286 = _2093 ^ _3656;
  wire _30287 = uncoded_block[973] ^ uncoded_block[977];
  wire _30288 = _30287 ^ _2100;
  wire _30289 = _30286 ^ _30288;
  wire _30290 = _30285 ^ _30289;
  wire _30291 = uncoded_block[981] ^ uncoded_block[986];
  wire _30292 = _30291 ^ _8859;
  wire _30293 = _2883 ^ _11101;
  wire _30294 = _30292 ^ _30293;
  wire _30295 = _15858 ^ _8866;
  wire _30296 = _30295 ^ _22589;
  wire _30297 = _30294 ^ _30296;
  wire _30298 = _30290 ^ _30297;
  wire _30299 = _30283 ^ _30298;
  wire _30300 = _30265 ^ _30299;
  wire _30301 = _30231 ^ _30300;
  wire _30302 = _30163 ^ _30301;
  wire _30303 = _9996 ^ _11663;
  wire _30304 = _2120 ^ _5137;
  wire _30305 = _30303 ^ _30304;
  wire _30306 = uncoded_block[1032] ^ uncoded_block[1037];
  wire _30307 = _2898 ^ _30306;
  wire _30308 = _511 ^ _17855;
  wire _30309 = _30307 ^ _30308;
  wire _30310 = _30305 ^ _30309;
  wire _30311 = _2136 ^ _8884;
  wire _30312 = _11120 ^ _8889;
  wire _30313 = _30311 ^ _30312;
  wire _30314 = _5158 ^ _5162;
  wire _30315 = _7724 ^ _533;
  wire _30316 = _30314 ^ _30315;
  wire _30317 = _30313 ^ _30316;
  wire _30318 = _30310 ^ _30317;
  wire _30319 = _11687 ^ _1374;
  wire _30320 = _536 ^ _7129;
  wire _30321 = _30319 ^ _30320;
  wire _30322 = _546 ^ _3708;
  wire _30323 = _22612 ^ _30322;
  wire _30324 = _30321 ^ _30323;
  wire _30325 = _2164 ^ _14882;
  wire _30326 = uncoded_block[1116] ^ uncoded_block[1121];
  wire _30327 = _30326 ^ _2942;
  wire _30328 = _30325 ^ _30327;
  wire _30329 = uncoded_block[1134] ^ uncoded_block[1140];
  wire _30330 = _30329 ^ _5859;
  wire _30331 = _23083 ^ _30330;
  wire _30332 = _30328 ^ _30331;
  wire _30333 = _30324 ^ _30332;
  wire _30334 = _30318 ^ _30333;
  wire _30335 = _3724 ^ _15902;
  wire _30336 = _2186 ^ _3728;
  wire _30337 = _30335 ^ _30336;
  wire _30338 = _578 ^ _7748;
  wire _30339 = _22627 ^ _6511;
  wire _30340 = _30338 ^ _30339;
  wire _30341 = _30337 ^ _30340;
  wire _30342 = _4481 ^ _3747;
  wire _30343 = _27538 ^ _30342;
  wire _30344 = uncoded_block[1198] ^ uncoded_block[1205];
  wire _30345 = _3749 ^ _30344;
  wire _30346 = uncoded_block[1206] ^ uncoded_block[1210];
  wire _30347 = _30346 ^ _26694;
  wire _30348 = _30345 ^ _30347;
  wire _30349 = _30343 ^ _30348;
  wire _30350 = _30341 ^ _30349;
  wire _30351 = uncoded_block[1213] ^ uncoded_block[1216];
  wire _30352 = uncoded_block[1217] ^ uncoded_block[1220];
  wire _30353 = _30351 ^ _30352;
  wire _30354 = _30353 ^ _4503;
  wire _30355 = uncoded_block[1242] ^ uncoded_block[1249];
  wire _30356 = _615 ^ _30355;
  wire _30357 = _13358 ^ _30356;
  wire _30358 = _30354 ^ _30357;
  wire _30359 = _7778 ^ _22651;
  wire _30360 = _30359 ^ _7782;
  wire _30361 = uncoded_block[1261] ^ uncoded_block[1263];
  wire _30362 = _30361 ^ _6550;
  wire _30363 = uncoded_block[1268] ^ uncoded_block[1271];
  wire _30364 = _30363 ^ _9538;
  wire _30365 = _30362 ^ _30364;
  wire _30366 = _30360 ^ _30365;
  wire _30367 = _30358 ^ _30366;
  wire _30368 = _30350 ^ _30367;
  wire _30369 = _30334 ^ _30368;
  wire _30370 = _5908 ^ _19365;
  wire _30371 = _11195 ^ _7194;
  wire _30372 = _30370 ^ _30371;
  wire _30373 = _646 ^ _22665;
  wire _30374 = _8991 ^ _7804;
  wire _30375 = _30373 ^ _30374;
  wire _30376 = _30372 ^ _30375;
  wire _30377 = _18426 ^ _4543;
  wire _30378 = _10655 ^ _2269;
  wire _30379 = _30377 ^ _30378;
  wire _30380 = _23576 ^ _13927;
  wire _30381 = _9003 ^ _5268;
  wire _30382 = _30380 ^ _30381;
  wire _30383 = _30379 ^ _30382;
  wire _30384 = _30376 ^ _30383;
  wire _30385 = _672 ^ _1504;
  wire _30386 = _2284 ^ _11226;
  wire _30387 = _30385 ^ _30386;
  wire _30388 = _2289 ^ _20334;
  wire _30389 = _11781 ^ _12311;
  wire _30390 = _30388 ^ _30389;
  wire _30391 = _30387 ^ _30390;
  wire _30392 = _3838 ^ _4568;
  wire _30393 = _20340 ^ _4572;
  wire _30394 = _30392 ^ _30393;
  wire _30395 = _2297 ^ _2299;
  wire _30396 = _30395 ^ _5958;
  wire _30397 = _30394 ^ _30396;
  wire _30398 = _30391 ^ _30397;
  wire _30399 = _30384 ^ _30398;
  wire _30400 = _4580 ^ _15492;
  wire _30401 = _2306 ^ _13428;
  wire _30402 = _30400 ^ _30401;
  wire _30403 = uncoded_block[1428] ^ uncoded_block[1431];
  wire _30404 = _709 ^ _30403;
  wire _30405 = _4586 ^ _2314;
  wire _30406 = _30404 ^ _30405;
  wire _30407 = _30402 ^ _30406;
  wire _30408 = _17470 ^ _20355;
  wire _30409 = uncoded_block[1450] ^ uncoded_block[1457];
  wire _30410 = _16969 ^ _30409;
  wire _30411 = _30408 ^ _30410;
  wire _30412 = _7241 ^ _22703;
  wire _30413 = _7247 ^ _22707;
  wire _30414 = _30412 ^ _30413;
  wire _30415 = _30411 ^ _30414;
  wire _30416 = _30407 ^ _30415;
  wire _30417 = _3101 ^ _1565;
  wire _30418 = _20864 ^ _30417;
  wire _30419 = uncoded_block[1495] ^ uncoded_block[1498];
  wire _30420 = _30419 ^ _747;
  wire _30421 = _3111 ^ _3894;
  wire _30422 = _30420 ^ _30421;
  wire _30423 = _30418 ^ _30422;
  wire _30424 = _23624 ^ _1575;
  wire _30425 = uncoded_block[1514] ^ uncoded_block[1520];
  wire _30426 = _30425 ^ _8473;
  wire _30427 = _30424 ^ _30426;
  wire _30428 = _4623 ^ _1582;
  wire _30429 = uncoded_block[1537] ^ uncoded_block[1542];
  wire _30430 = _11820 ^ _30429;
  wire _30431 = _30428 ^ _30430;
  wire _30432 = _30427 ^ _30431;
  wire _30433 = _30423 ^ _30432;
  wire _30434 = _30416 ^ _30433;
  wire _30435 = _30399 ^ _30434;
  wire _30436 = _30369 ^ _30435;
  wire _30437 = uncoded_block[1543] ^ uncoded_block[1547];
  wire _30438 = _30437 ^ _13472;
  wire _30439 = _30438 ^ _771;
  wire _30440 = _26794 ^ _5361;
  wire _30441 = _29986 ^ _25895;
  wire _30442 = _30440 ^ _30441;
  wire _30443 = _30439 ^ _30442;
  wire _30444 = _15026 ^ _4647;
  wire _30445 = _4648 ^ _4651;
  wire _30446 = _30444 ^ _30445;
  wire _30447 = _12369 ^ _3145;
  wire _30448 = _3146 ^ _2394;
  wire _30449 = _30447 ^ _30448;
  wire _30450 = _30446 ^ _30449;
  wire _30451 = _30443 ^ _30450;
  wire _30452 = _3934 ^ _3151;
  wire _30453 = _30452 ^ _6678;
  wire _30454 = _18020 ^ _13494;
  wire _30455 = uncoded_block[1631] ^ uncoded_block[1635];
  wire _30456 = _18511 ^ _30455;
  wire _30457 = _30454 ^ _30456;
  wire _30458 = _30453 ^ _30457;
  wire _30459 = _18969 ^ _1650;
  wire _30460 = _16532 ^ _30459;
  wire _30461 = _10760 ^ _3174;
  wire _30462 = _3958 ^ _7319;
  wire _30463 = _30461 ^ _30462;
  wire _30464 = _30460 ^ _30463;
  wire _30465 = _30458 ^ _30464;
  wire _30466 = _30451 ^ _30465;
  wire _30467 = _4687 ^ _19471;
  wire _30468 = _30467 ^ _17037;
  wire _30469 = _7936 ^ _20434;
  wire _30470 = _30468 ^ _30469;
  wire _30471 = _16550 ^ _12406;
  wire _30472 = _25487 ^ _17554;
  wire _30473 = _30471 ^ _30472;
  wire _30474 = _30470 ^ _30473;
  wire _30475 = _30466 ^ _30474;
  wire _30476 = _30436 ^ _30475;
  wire _30477 = _30302 ^ _30476;
  wire _30478 = _3 ^ _3213;
  wire _30479 = _3211 ^ _30478;
  wire _30480 = _28748 ^ _3221;
  wire _30481 = _30479 ^ _30480;
  wire _30482 = _7959 ^ _2461;
  wire _30483 = _15 ^ _8549;
  wire _30484 = _30482 ^ _30483;
  wire _30485 = uncoded_block[43] ^ uncoded_block[47];
  wire _30486 = _21871 ^ _30485;
  wire _30487 = _1699 ^ _25;
  wire _30488 = _30486 ^ _30487;
  wire _30489 = _30484 ^ _30488;
  wire _30490 = _30481 ^ _30489;
  wire _30491 = _15087 ^ _7364;
  wire _30492 = _8559 ^ _7367;
  wire _30493 = _30491 ^ _30492;
  wire _30494 = _14058 ^ _1712;
  wire _30495 = _28765 ^ _2483;
  wire _30496 = _30494 ^ _30495;
  wire _30497 = _30493 ^ _30496;
  wire _30498 = uncoded_block[92] ^ uncoded_block[96];
  wire _30499 = _30498 ^ _6116;
  wire _30500 = _19021 ^ _30499;
  wire _30501 = _17583 ^ _6122;
  wire _30502 = _20957 ^ _6126;
  wire _30503 = _30501 ^ _30502;
  wire _30504 = _30500 ^ _30503;
  wire _30505 = _30497 ^ _30504;
  wire _30506 = _30490 ^ _30505;
  wire _30507 = _2495 ^ _4750;
  wire _30508 = _10256 ^ _57;
  wire _30509 = _30507 ^ _30508;
  wire _30510 = _4754 ^ _924;
  wire _30511 = uncoded_block[138] ^ uncoded_block[142];
  wire _30512 = _20969 ^ _30511;
  wire _30513 = _30510 ^ _30512;
  wire _30514 = _30509 ^ _30513;
  wire _30515 = _7392 ^ _15622;
  wire _30516 = uncoded_block[153] ^ uncoded_block[157];
  wire _30517 = _1745 ^ _30516;
  wire _30518 = _30515 ^ _30517;
  wire _30519 = uncoded_block[163] ^ uncoded_block[167];
  wire _30520 = _9188 ^ _30519;
  wire _30521 = _1752 ^ _19539;
  wire _30522 = _30520 ^ _30521;
  wire _30523 = _30518 ^ _30522;
  wire _30524 = _30514 ^ _30523;
  wire _30525 = _28037 ^ _15631;
  wire _30526 = _7404 ^ _30525;
  wire _30527 = _5483 ^ _18583;
  wire _30528 = uncoded_block[201] ^ uncoded_block[207];
  wire _30529 = _6801 ^ _30528;
  wire _30530 = _30527 ^ _30529;
  wire _30531 = _30526 ^ _30530;
  wire _30532 = _97 ^ _956;
  wire _30533 = _9202 ^ _3299;
  wire _30534 = _30532 ^ _30533;
  wire _30535 = _4084 ^ _10860;
  wire _30536 = _22381 ^ _30535;
  wire _30537 = _30534 ^ _30536;
  wire _30538 = _30531 ^ _30537;
  wire _30539 = _30524 ^ _30538;
  wire _30540 = _30506 ^ _30539;
  wire _30541 = _11952 ^ _974;
  wire _30542 = _13053 ^ _3311;
  wire _30543 = _30541 ^ _30542;
  wire _30544 = _13055 ^ _120;
  wire _30545 = _6188 ^ _127;
  wire _30546 = _30544 ^ _30545;
  wire _30547 = _30543 ^ _30546;
  wire _30548 = uncoded_block[270] ^ uncoded_block[274];
  wire _30549 = _30548 ^ _1795;
  wire _30550 = _12506 ^ _7446;
  wire _30551 = _30549 ^ _30550;
  wire _30552 = _5524 ^ _999;
  wire _30553 = _9773 ^ _30552;
  wire _30554 = _30551 ^ _30553;
  wire _30555 = _30547 ^ _30554;
  wire _30556 = _17639 ^ _21017;
  wire _30557 = uncoded_block[311] ^ uncoded_block[318];
  wire _30558 = _30557 ^ _6850;
  wire _30559 = _30556 ^ _30558;
  wire _30560 = _15677 ^ _1014;
  wire _30561 = _4837 ^ _1821;
  wire _30562 = _30560 ^ _30561;
  wire _30563 = _30559 ^ _30562;
  wire _30564 = uncoded_block[343] ^ uncoded_block[347];
  wire _30565 = _30564 ^ _3359;
  wire _30566 = _12525 ^ _30565;
  wire _30567 = uncoded_block[355] ^ uncoded_block[359];
  wire _30568 = _30567 ^ _12530;
  wire _30569 = uncoded_block[365] ^ uncoded_block[370];
  wire _30570 = _5548 ^ _30569;
  wire _30571 = _30568 ^ _30570;
  wire _30572 = _30566 ^ _30571;
  wire _30573 = _30563 ^ _30572;
  wire _30574 = _30555 ^ _30573;
  wire _30575 = _4140 ^ _7474;
  wire _30576 = _30575 ^ _29679;
  wire _30577 = _1039 ^ _2613;
  wire _30578 = _21504 ^ _6881;
  wire _30579 = _30577 ^ _30578;
  wire _30580 = _30576 ^ _30579;
  wire _30581 = _2622 ^ _12545;
  wire _30582 = _4867 ^ _14682;
  wire _30583 = _30581 ^ _30582;
  wire _30584 = _8671 ^ _9816;
  wire _30585 = _4167 ^ _200;
  wire _30586 = _30584 ^ _30585;
  wire _30587 = _30583 ^ _30586;
  wire _30588 = _30580 ^ _30587;
  wire _30589 = _21049 ^ _12559;
  wire _30590 = _30589 ^ _17183;
  wire _30591 = uncoded_block[456] ^ uncoded_block[464];
  wire _30592 = _2645 ^ _30591;
  wire _30593 = _8683 ^ _21523;
  wire _30594 = _30592 ^ _30593;
  wire _30595 = _30590 ^ _30594;
  wire _30596 = _15211 ^ _8111;
  wire _30597 = _19127 ^ _30596;
  wire _30598 = _9833 ^ _9836;
  wire _30599 = _30597 ^ _30598;
  wire _30600 = _30595 ^ _30599;
  wire _30601 = _30588 ^ _30600;
  wire _30602 = _30574 ^ _30601;
  wire _30603 = _30540 ^ _30602;
  wire _30604 = uncoded_block[501] ^ uncoded_block[506];
  wire _30605 = uncoded_block[507] ^ uncoded_block[511];
  wire _30606 = _30604 ^ _30605;
  wire _30607 = _15220 ^ _8706;
  wire _30608 = _30606 ^ _30607;
  wire _30609 = uncoded_block[528] ^ uncoded_block[534];
  wire _30610 = _1900 ^ _30609;
  wire _30611 = _3446 ^ _30610;
  wire _30612 = _30608 ^ _30611;
  wire _30613 = _5619 ^ _6293;
  wire _30614 = _1908 ^ _22934;
  wire _30615 = _30613 ^ _30614;
  wire _30616 = _20110 ^ _20615;
  wire _30617 = _4939 ^ _30616;
  wire _30618 = _30615 ^ _30617;
  wire _30619 = _30612 ^ _30618;
  wire _30620 = uncoded_block[580] ^ uncoded_block[587];
  wire _30621 = _30620 ^ _271;
  wire _30622 = _1932 ^ _30621;
  wire _30623 = _4236 ^ _4952;
  wire _30624 = uncoded_block[601] ^ uncoded_block[611];
  wire _30625 = _30624 ^ _7563;
  wire _30626 = _30623 ^ _30625;
  wire _30627 = _30622 ^ _30626;
  wire _30628 = _1149 ^ _6959;
  wire _30629 = _1154 ^ _30199;
  wire _30630 = _30628 ^ _30629;
  wire _30631 = _29741 ^ _4256;
  wire _30632 = _30631 ^ _9883;
  wire _30633 = _30630 ^ _30632;
  wire _30634 = _30627 ^ _30633;
  wire _30635 = _30619 ^ _30634;
  wire _30636 = _13726 ^ _7586;
  wire _30637 = _16750 ^ _30636;
  wire _30638 = _17745 ^ _1968;
  wire _30639 = _30638 ^ _9360;
  wire _30640 = _30637 ^ _30639;
  wire _30641 = uncoded_block[695] ^ uncoded_block[699];
  wire _30642 = _30641 ^ _333;
  wire _30643 = _19681 ^ _30642;
  wire _30644 = _3535 ^ _19201;
  wire _30645 = uncoded_block[719] ^ uncoded_block[722];
  wire _30646 = _1195 ^ _30645;
  wire _30647 = _30644 ^ _30646;
  wire _30648 = _30643 ^ _30647;
  wire _30649 = _30640 ^ _30648;
  wire _30650 = _6374 ^ _10457;
  wire _30651 = uncoded_block[730] ^ uncoded_block[734];
  wire _30652 = _30651 ^ _350;
  wire _30653 = _30650 ^ _30652;
  wire _30654 = _5704 ^ _13754;
  wire _30655 = _27820 ^ _30654;
  wire _30656 = _30653 ^ _30655;
  wire _30657 = uncoded_block[759] ^ uncoded_block[763];
  wire _30658 = _30657 ^ _10470;
  wire _30659 = uncoded_block[769] ^ uncoded_block[772];
  wire _30660 = _30659 ^ _5711;
  wire _30661 = _30658 ^ _30660;
  wire _30662 = _2014 ^ _2018;
  wire _30663 = _1225 ^ _21614;
  wire _30664 = _30662 ^ _30663;
  wire _30665 = _30661 ^ _30664;
  wire _30666 = _30656 ^ _30665;
  wire _30667 = _30649 ^ _30666;
  wire _30668 = _30635 ^ _30667;
  wire _30669 = _4316 ^ _26589;
  wire _30670 = _8793 ^ _10485;
  wire _30671 = _30669 ^ _30670;
  wire _30672 = _19717 ^ _14290;
  wire _30673 = _1246 ^ _5052;
  wire _30674 = _30672 ^ _30673;
  wire _30675 = _30671 ^ _30674;
  wire _30676 = _16801 ^ _4337;
  wire _30677 = _5737 ^ _14812;
  wire _30678 = _30676 ^ _30677;
  wire _30679 = _5741 ^ _11048;
  wire _30680 = uncoded_block[855] ^ uncoded_block[858];
  wire _30681 = _30680 ^ _9948;
  wire _30682 = _30679 ^ _30681;
  wire _30683 = _30678 ^ _30682;
  wire _30684 = _30675 ^ _30683;
  wire _30685 = _26171 ^ _12150;
  wire _30686 = _30685 ^ _14307;
  wire _30687 = _2835 ^ _3610;
  wire _30688 = _30687 ^ _5084;
  wire _30689 = _30686 ^ _30688;
  wire _30690 = _5085 ^ _3617;
  wire _30691 = _8827 ^ _3623;
  wire _30692 = _30690 ^ _30691;
  wire _30693 = _17318 ^ _4368;
  wire _30694 = _25730 ^ _30693;
  wire _30695 = _30692 ^ _30694;
  wire _30696 = _30689 ^ _30695;
  wire _30697 = _30684 ^ _30696;
  wire _30698 = _1295 ^ _9968;
  wire _30699 = uncoded_block[932] ^ uncoded_block[939];
  wire _30700 = _30699 ^ _453;
  wire _30701 = _30698 ^ _30700;
  wire _30702 = _13263 ^ _23926;
  wire _30703 = _8274 ^ _12726;
  wire _30704 = _30702 ^ _30703;
  wire _30705 = _30701 ^ _30704;
  wire _30706 = _4385 ^ _12180;
  wire _30707 = _6447 ^ _4390;
  wire _30708 = _30706 ^ _30707;
  wire _30709 = _471 ^ _5792;
  wire _30710 = _6451 ^ _16338;
  wire _30711 = _30709 ^ _30710;
  wire _30712 = _30708 ^ _30711;
  wire _30713 = _30705 ^ _30712;
  wire _30714 = _3663 ^ _5798;
  wire _30715 = _30714 ^ _9450;
  wire _30716 = uncoded_block[1017] ^ uncoded_block[1025];
  wire _30717 = _2117 ^ _30716;
  wire _30718 = _488 ^ _30717;
  wire _30719 = _30715 ^ _30718;
  wire _30720 = _4417 ^ _12198;
  wire _30721 = _8876 ^ _30720;
  wire _30722 = _6475 ^ _8309;
  wire _30723 = _2134 ^ _518;
  wire _30724 = _30722 ^ _30723;
  wire _30725 = _30721 ^ _30724;
  wire _30726 = _30719 ^ _30725;
  wire _30727 = _30713 ^ _30726;
  wire _30728 = _30697 ^ _30727;
  wire _30729 = _30668 ^ _30728;
  wire _30730 = _30603 ^ _30729;
  wire _30731 = uncoded_block[1055] ^ uncoded_block[1060];
  wire _30732 = _1359 ^ _30731;
  wire _30733 = _10569 ^ _11122;
  wire _30734 = _30732 ^ _30733;
  wire _30735 = _8892 ^ _5831;
  wire _30736 = _30735 ^ _8324;
  wire _30737 = _30734 ^ _30736;
  wire _30738 = uncoded_block[1083] ^ uncoded_block[1087];
  wire _30739 = _7724 ^ _30738;
  wire _30740 = uncoded_block[1088] ^ uncoded_block[1092];
  wire _30741 = _30740 ^ _10026;
  wire _30742 = _30739 ^ _30741;
  wire _30743 = _545 ^ _11142;
  wire _30744 = _3708 ^ _550;
  wire _30745 = _30743 ^ _30744;
  wire _30746 = _30742 ^ _30745;
  wire _30747 = _30737 ^ _30746;
  wire _30748 = uncoded_block[1116] ^ uncoded_block[1122];
  wire _30749 = _8917 ^ _30748;
  wire _30750 = _1392 ^ _4460;
  wire _30751 = _30749 ^ _30750;
  wire _30752 = _23084 ^ _7139;
  wire _30753 = _30751 ^ _30752;
  wire _30754 = _7141 ^ _8351;
  wire _30755 = _30754 ^ _24901;
  wire _30756 = uncoded_block[1164] ^ uncoded_block[1168];
  wire _30757 = _8356 ^ _30756;
  wire _30758 = _9506 ^ _3739;
  wire _30759 = _30757 ^ _30758;
  wire _30760 = _30755 ^ _30759;
  wire _30761 = _30753 ^ _30760;
  wire _30762 = _30747 ^ _30761;
  wire _30763 = _585 ^ _589;
  wire _30764 = _590 ^ _5200;
  wire _30765 = _30763 ^ _30764;
  wire _30766 = _3747 ^ _10612;
  wire _30767 = _12810 ^ _7162;
  wire _30768 = _30766 ^ _30767;
  wire _30769 = _30765 ^ _30768;
  wire _30770 = _2209 ^ _2216;
  wire _30771 = _1427 ^ _3762;
  wire _30772 = _30770 ^ _30771;
  wire _30773 = uncoded_block[1223] ^ uncoded_block[1226];
  wire _30774 = _14407 ^ _30773;
  wire _30775 = _13357 ^ _18400;
  wire _30776 = _30774 ^ _30775;
  wire _30777 = _30772 ^ _30776;
  wire _30778 = _30769 ^ _30777;
  wire _30779 = _5219 ^ _3771;
  wire _30780 = _3772 ^ _2994;
  wire _30781 = _30779 ^ _30780;
  wire _30782 = _6538 ^ _5229;
  wire _30783 = _5901 ^ _3780;
  wire _30784 = _30782 ^ _30783;
  wire _30785 = _30781 ^ _30784;
  wire _30786 = _6550 ^ _9532;
  wire _30787 = _11743 ^ _30786;
  wire _30788 = _2245 ^ _4523;
  wire _30789 = uncoded_block[1275] ^ uncoded_block[1278];
  wire _30790 = _30789 ^ _631;
  wire _30791 = _30788 ^ _30790;
  wire _30792 = _30787 ^ _30791;
  wire _30793 = _30785 ^ _30792;
  wire _30794 = _30778 ^ _30793;
  wire _30795 = _30762 ^ _30794;
  wire _30796 = _6557 ^ _11195;
  wire _30797 = uncoded_block[1292] ^ uncoded_block[1294];
  wire _30798 = _30797 ^ _4532;
  wire _30799 = _30796 ^ _30798;
  wire _30800 = uncoded_block[1310] ^ uncoded_block[1314];
  wire _30801 = _2259 ^ _30800;
  wire _30802 = _21748 ^ _23134;
  wire _30803 = _30801 ^ _30802;
  wire _30804 = _30799 ^ _30803;
  wire _30805 = _9555 ^ _656;
  wire _30806 = _10655 ^ _1494;
  wire _30807 = _30805 ^ _30806;
  wire _30808 = _18431 ^ _9563;
  wire _30809 = _30808 ^ _1499;
  wire _30810 = _30807 ^ _30809;
  wire _30811 = _30804 ^ _30810;
  wire _30812 = _21302 ^ _28331;
  wire _30813 = _23581 ^ _27157;
  wire _30814 = _5281 ^ _3832;
  wire _30815 = _30813 ^ _30814;
  wire _30816 = _30812 ^ _30815;
  wire _30817 = _13410 ^ _3835;
  wire _30818 = uncoded_block[1392] ^ uncoded_block[1396];
  wire _30819 = _24511 ^ _30818;
  wire _30820 = _30817 ^ _30819;
  wire _30821 = uncoded_block[1397] ^ uncoded_block[1403];
  wire _30822 = _30821 ^ _4578;
  wire _30823 = _701 ^ _8436;
  wire _30824 = _30822 ^ _30823;
  wire _30825 = _30820 ^ _30824;
  wire _30826 = _30816 ^ _30825;
  wire _30827 = _30811 ^ _30826;
  wire _30828 = uncoded_block[1411] ^ uncoded_block[1416];
  wire _30829 = _30828 ^ _10120;
  wire _30830 = _9588 ^ _14466;
  wire _30831 = _30829 ^ _30830;
  wire _30832 = _2314 ^ _3861;
  wire _30833 = _12326 ^ _30832;
  wire _30834 = _30831 ^ _30833;
  wire _30835 = _6613 ^ _8450;
  wire _30836 = uncoded_block[1452] ^ uncoded_block[1462];
  wire _30837 = _3865 ^ _30836;
  wire _30838 = _30835 ^ _30837;
  wire _30839 = _22254 ^ _11255;
  wire _30840 = _5316 ^ _13446;
  wire _30841 = _30839 ^ _30840;
  wire _30842 = _30838 ^ _30841;
  wire _30843 = _30834 ^ _30842;
  wire _30844 = uncoded_block[1485] ^ uncoded_block[1491];
  wire _30845 = _23181 ^ _30844;
  wire _30846 = _2350 ^ _2352;
  wire _30847 = _30845 ^ _30846;
  wire _30848 = uncoded_block[1502] ^ uncoded_block[1505];
  wire _30849 = _30848 ^ _3112;
  wire _30850 = _6637 ^ _19429;
  wire _30851 = _30849 ^ _30850;
  wire _30852 = _30847 ^ _30851;
  wire _30853 = _5337 ^ _15004;
  wire _30854 = uncoded_block[1526] ^ uncoded_block[1530];
  wire _30855 = _16988 ^ _30854;
  wire _30856 = _30853 ^ _30855;
  wire _30857 = _28375 ^ _3909;
  wire _30858 = uncoded_block[1544] ^ uncoded_block[1548];
  wire _30859 = _30858 ^ _14496;
  wire _30860 = _30857 ^ _30859;
  wire _30861 = _30856 ^ _30860;
  wire _30862 = _30852 ^ _30861;
  wire _30863 = _30843 ^ _30862;
  wire _30864 = _30827 ^ _30863;
  wire _30865 = _30795 ^ _30864;
  wire _30866 = _769 ^ _6016;
  wire _30867 = _4640 ^ _5361;
  wire _30868 = _30866 ^ _30867;
  wire _30869 = _20392 ^ _16510;
  wire _30870 = uncoded_block[1571] ^ uncoded_block[1573];
  wire _30871 = _30870 ^ _4648;
  wire _30872 = _30869 ^ _30871;
  wire _30873 = _30868 ^ _30872;
  wire _30874 = _6663 ^ _17009;
  wire _30875 = uncoded_block[1589] ^ uncoded_block[1594];
  wire _30876 = _30875 ^ _13486;
  wire _30877 = _30874 ^ _30876;
  wire _30878 = _26343 ^ _3157;
  wire _30879 = _10181 ^ _12376;
  wire _30880 = _30878 ^ _30879;
  wire _30881 = _30877 ^ _30880;
  wire _30882 = _30873 ^ _30881;
  wire _30883 = _14525 ^ _1639;
  wire _30884 = _24573 ^ _30883;
  wire _30885 = _812 ^ _10754;
  wire _30886 = _3948 ^ _815;
  wire _30887 = _30885 ^ _30886;
  wire _30888 = _30884 ^ _30887;
  wire _30889 = uncoded_block[1648] ^ uncoded_block[1658];
  wire _30890 = _816 ^ _30889;
  wire _30891 = uncoded_block[1661] ^ uncoded_block[1666];
  wire _30892 = _30891 ^ _8521;
  wire _30893 = _30890 ^ _30892;
  wire _30894 = _7323 ^ _10766;
  wire _30895 = _17040 ^ _3965;
  wire _30896 = _30894 ^ _30895;
  wire _30897 = _30893 ^ _30896;
  wire _30898 = _30888 ^ _30897;
  wire _30899 = _30882 ^ _30898;
  wire _30900 = uncoded_block[1688] ^ uncoded_block[1691];
  wire _30901 = _30900 ^ _840;
  wire _30902 = _844 ^ _24137;
  wire _30903 = _30901 ^ _30902;
  wire _30904 = _8535 ^ _5412;
  wire _30905 = _851 ^ _7337;
  wire _30906 = _30904 ^ _30905;
  wire _30907 = _30903 ^ _30906;
  wire _30908 = uncoded_block[1713] ^ uncoded_block[1716];
  wire _30909 = _30908 ^ _20923;
  wire _30910 = _30909 ^ uncoded_block[1720];
  wire _30911 = _30907 ^ _30910;
  wire _30912 = _30899 ^ _30911;
  wire _30913 = _30865 ^ _30912;
  wire _30914 = _30730 ^ _30913;
  wire _30915 = _3995 ^ _19001;
  wire _30916 = _22325 ^ _30915;
  wire _30917 = _871 ^ _10226;
  wire _30918 = uncoded_block[22] ^ uncoded_block[28];
  wire _30919 = _1690 ^ _30918;
  wire _30920 = _30917 ^ _30919;
  wire _30921 = _30916 ^ _30920;
  wire _30922 = _5429 ^ _19501;
  wire _30923 = _14571 ^ _6736;
  wire _30924 = _30922 ^ _30923;
  wire _30925 = _5433 ^ _8556;
  wire _30926 = _20465 ^ _10806;
  wire _30927 = _30925 ^ _30926;
  wire _30928 = _30924 ^ _30927;
  wire _30929 = _30921 ^ _30928;
  wire _30930 = _896 ^ _4733;
  wire _30931 = _25510 ^ _30930;
  wire _30932 = _7979 ^ _41;
  wire _30933 = _2484 ^ _9713;
  wire _30934 = _30932 ^ _30933;
  wire _30935 = _30931 ^ _30934;
  wire _30936 = _903 ^ _10251;
  wire _30937 = _6122 ^ _2491;
  wire _30938 = _30936 ^ _30937;
  wire _30939 = _5453 ^ _7990;
  wire _30940 = _30939 ^ _12452;
  wire _30941 = _30938 ^ _30940;
  wire _30942 = _30935 ^ _30941;
  wire _30943 = _30929 ^ _30942;
  wire _30944 = _8579 ^ _15112;
  wire _30945 = uncoded_block[143] ^ uncoded_block[146];
  wire _30946 = _9180 ^ _30945;
  wire _30947 = _30944 ^ _30946;
  wire _30948 = _14082 ^ _3269;
  wire _30949 = _30948 ^ _7398;
  wire _30950 = _30947 ^ _30949;
  wire _30951 = uncoded_block[158] ^ uncoded_block[161];
  wire _30952 = _30951 ^ _4054;
  wire _30953 = _29624 ^ _8591;
  wire _30954 = _30952 ^ _30953;
  wire _30955 = _14614 ^ _6149;
  wire _30956 = uncoded_block[183] ^ uncoded_block[187];
  wire _30957 = _11933 ^ _30956;
  wire _30958 = _30955 ^ _30957;
  wire _30959 = _30954 ^ _30958;
  wire _30960 = _30950 ^ _30959;
  wire _30961 = _18583 ^ _6801;
  wire _30962 = _23288 ^ _30961;
  wire _30963 = uncoded_block[207] ^ uncoded_block[211];
  wire _30964 = _30963 ^ _3295;
  wire _30965 = _17610 ^ _30964;
  wire _30966 = _30962 ^ _30965;
  wire _30967 = _28046 ^ _9206;
  wire _30968 = _6169 ^ _9208;
  wire _30969 = _30967 ^ _30968;
  wire _30970 = _112 ^ _3308;
  wire _30971 = _4088 ^ _119;
  wire _30972 = _30970 ^ _30971;
  wire _30973 = _30969 ^ _30972;
  wire _30974 = _30966 ^ _30973;
  wire _30975 = _30960 ^ _30974;
  wire _30976 = _30943 ^ _30975;
  wire _30977 = _6831 ^ _6188;
  wire _30978 = _127 ^ _130;
  wire _30979 = _30977 ^ _30978;
  wire _30980 = _12506 ^ _4105;
  wire _30981 = _30980 ^ _26902;
  wire _30982 = _30979 ^ _30981;
  wire _30983 = _10876 ^ _2573;
  wire _30984 = _138 ^ _8052;
  wire _30985 = _30983 ^ _30984;
  wire _30986 = _1002 ^ _3337;
  wire _30987 = _15671 ^ _4830;
  wire _30988 = _30986 ^ _30987;
  wire _30989 = _30985 ^ _30988;
  wire _30990 = _30982 ^ _30989;
  wire _30991 = uncoded_block[321] ^ uncoded_block[329];
  wire _30992 = _30991 ^ _4125;
  wire _30993 = _30992 ^ _9787;
  wire _30994 = _9242 ^ _1021;
  wire _30995 = _4131 ^ _1023;
  wire _30996 = _30994 ^ _30995;
  wire _30997 = _30993 ^ _30996;
  wire _30998 = _6864 ^ _26032;
  wire _30999 = uncoded_block[367] ^ uncoded_block[374];
  wire _31000 = _30999 ^ _4854;
  wire _31001 = _30998 ^ _31000;
  wire _31002 = _26030 ^ _31001;
  wire _31003 = _30997 ^ _31002;
  wire _31004 = _30990 ^ _31003;
  wire _31005 = uncoded_block[385] ^ uncoded_block[388];
  wire _31006 = _31005 ^ _6879;
  wire _31007 = _3378 ^ _31006;
  wire _31008 = _26925 ^ _1051;
  wire _31009 = _26479 ^ _31008;
  wire _31010 = _31007 ^ _31009;
  wire _31011 = uncoded_block[408] ^ uncoded_block[418];
  wire _31012 = _31011 ^ _4872;
  wire _31013 = _4164 ^ _8672;
  wire _31014 = _31012 ^ _31013;
  wire _31015 = _9816 ^ _4167;
  wire _31016 = _31015 ^ _26052;
  wire _31017 = _31014 ^ _31016;
  wire _31018 = _31010 ^ _31017;
  wire _31019 = _21974 ^ _16191;
  wire _31020 = _21973 ^ _31019;
  wire _31021 = _1870 ^ _10926;
  wire _31022 = _19622 ^ _31021;
  wire _31023 = _31020 ^ _31022;
  wire _31024 = uncoded_block[467] ^ uncoded_block[472];
  wire _31025 = _7507 ^ _31024;
  wire _31026 = _31025 ^ _1087;
  wire _31027 = _1090 ^ _5600;
  wire _31028 = _1093 ^ _2667;
  wire _31029 = _31027 ^ _31028;
  wire _31030 = _31026 ^ _31029;
  wire _31031 = _31023 ^ _31030;
  wire _31032 = _31018 ^ _31031;
  wire _31033 = _31004 ^ _31032;
  wire _31034 = _30976 ^ _31033;
  wire _31035 = uncoded_block[502] ^ uncoded_block[506];
  wire _31036 = _31035 ^ _8701;
  wire _31037 = _31036 ^ _23371;
  wire _31038 = uncoded_block[519] ^ uncoded_block[523];
  wire _31039 = _31038 ^ _20602;
  wire _31040 = _240 ^ _27375;
  wire _31041 = _31039 ^ _31040;
  wire _31042 = _31037 ^ _31041;
  wire _31043 = _14721 ^ _24282;
  wire _31044 = _1913 ^ _8721;
  wire _31045 = _31043 ^ _31044;
  wire _31046 = _8724 ^ _4937;
  wire _31047 = _4938 ^ _3464;
  wire _31048 = _31046 ^ _31047;
  wire _31049 = _31045 ^ _31048;
  wire _31050 = _31042 ^ _31049;
  wire _31051 = _262 ^ _6947;
  wire _31052 = _5636 ^ _31051;
  wire _31053 = _266 ^ _4950;
  wire _31054 = _1938 ^ _8149;
  wire _31055 = _31053 ^ _31054;
  wire _31056 = _31052 ^ _31055;
  wire _31057 = _2707 ^ _2709;
  wire _31058 = _5647 ^ _6957;
  wire _31059 = _31057 ^ _31058;
  wire _31060 = uncoded_block[619] ^ uncoded_block[623];
  wire _31061 = _7567 ^ _31060;
  wire _31062 = _287 ^ _30199;
  wire _31063 = _31061 ^ _31062;
  wire _31064 = _31059 ^ _31063;
  wire _31065 = _31056 ^ _31064;
  wire _31066 = _31050 ^ _31065;
  wire _31067 = _28527 ^ _17243;
  wire _31068 = _2730 ^ _301;
  wire _31069 = _14755 ^ _3514;
  wire _31070 = _31068 ^ _31069;
  wire _31071 = _31067 ^ _31070;
  wire _31072 = uncoded_block[668] ^ uncoded_block[672];
  wire _31073 = _9885 ^ _31072;
  wire _31074 = _3519 ^ _13731;
  wire _31075 = _31073 ^ _31074;
  wire _31076 = uncoded_block[686] ^ uncoded_block[689];
  wire _31077 = _6352 ^ _31076;
  wire _31078 = _31077 ^ _15283;
  wire _31079 = _31075 ^ _31078;
  wire _31080 = _31071 ^ _31079;
  wire _31081 = _25218 ^ _4995;
  wire _31082 = _15285 ^ _31081;
  wire _31083 = _8190 ^ _2762;
  wire _31084 = _10452 ^ _17266;
  wire _31085 = _31083 ^ _31084;
  wire _31086 = _31082 ^ _31085;
  wire _31087 = _6367 ^ _9369;
  wire _31088 = _6374 ^ _5693;
  wire _31089 = _31087 ^ _31088;
  wire _31090 = _2768 ^ _4287;
  wire _31091 = _1995 ^ _350;
  wire _31092 = _31090 ^ _31091;
  wire _31093 = _31089 ^ _31092;
  wire _31094 = _31086 ^ _31093;
  wire _31095 = _31080 ^ _31094;
  wire _31096 = _31066 ^ _31095;
  wire _31097 = _2774 ^ _4293;
  wire _31098 = uncoded_block[754] ^ uncoded_block[759];
  wire _31099 = _1214 ^ _31098;
  wire _31100 = _31097 ^ _31099;
  wire _31101 = _9914 ^ _1217;
  wire _31102 = _4301 ^ _9917;
  wire _31103 = _31101 ^ _31102;
  wire _31104 = _31100 ^ _31103;
  wire _31105 = _1221 ^ _2014;
  wire _31106 = uncoded_block[781] ^ uncoded_block[785];
  wire _31107 = _7021 ^ _31106;
  wire _31108 = _31105 ^ _31107;
  wire _31109 = _3574 ^ _2021;
  wire _31110 = _5034 ^ _31109;
  wire _31111 = _31108 ^ _31110;
  wire _31112 = _31104 ^ _31111;
  wire _31113 = _15813 ^ _16287;
  wire _31114 = _2026 ^ _4324;
  wire _31115 = uncoded_block[816] ^ uncoded_block[822];
  wire _31116 = _31115 ^ _1247;
  wire _31117 = _31114 ^ _31116;
  wire _31118 = _31113 ^ _31117;
  wire _31119 = _7039 ^ _400;
  wire _31120 = _4336 ^ _14809;
  wire _31121 = _31119 ^ _31120;
  wire _31122 = _8808 ^ _3600;
  wire _31123 = uncoded_block[860] ^ uncoded_block[864];
  wire _31124 = _31123 ^ _414;
  wire _31125 = _31122 ^ _31124;
  wire _31126 = _31121 ^ _31125;
  wire _31127 = _31118 ^ _31126;
  wire _31128 = _31112 ^ _31127;
  wire _31129 = uncoded_block[867] ^ uncoded_block[871];
  wire _31130 = _31129 ^ _417;
  wire _31131 = uncoded_block[878] ^ uncoded_block[882];
  wire _31132 = uncoded_block[883] ^ uncoded_block[886];
  wire _31133 = _31131 ^ _31132;
  wire _31134 = _31130 ^ _31133;
  wire _31135 = _28962 ^ _4355;
  wire _31136 = _31135 ^ _4359;
  wire _31137 = _31134 ^ _31136;
  wire _31138 = _8254 ^ _30270;
  wire _31139 = _1287 ^ _3628;
  wire _31140 = _31138 ^ _31139;
  wire _31141 = uncoded_block[923] ^ uncoded_block[927];
  wire _31142 = _17318 ^ _31141;
  wire _31143 = _4371 ^ _5096;
  wire _31144 = _31142 ^ _31143;
  wire _31145 = _31140 ^ _31144;
  wire _31146 = _31137 ^ _31145;
  wire _31147 = _455 ^ _23926;
  wire _31148 = _454 ^ _31147;
  wire _31149 = _4381 ^ _12726;
  wire _31150 = _7086 ^ _7088;
  wire _31151 = _31149 ^ _31150;
  wire _31152 = _31148 ^ _31151;
  wire _31153 = _2877 ^ _28233;
  wire _31154 = _31153 ^ _4396;
  wire _31155 = uncoded_block[984] ^ uncoded_block[988];
  wire _31156 = _31155 ^ _2882;
  wire _31157 = _4401 ^ _479;
  wire _31158 = _31156 ^ _31157;
  wire _31159 = _31154 ^ _31158;
  wire _31160 = _31152 ^ _31159;
  wire _31161 = _31146 ^ _31160;
  wire _31162 = _31128 ^ _31161;
  wire _31163 = _31096 ^ _31162;
  wire _31164 = _31034 ^ _31163;
  wire _31165 = uncoded_block[996] ^ uncoded_block[999];
  wire _31166 = uncoded_block[1000] ^ uncoded_block[1004];
  wire _31167 = _31165 ^ _31166;
  wire _31168 = _31167 ^ _6460;
  wire _31169 = _2893 ^ _1334;
  wire _31170 = _5132 ^ _31169;
  wire _31171 = _31168 ^ _31170;
  wire _31172 = uncoded_block[1028] ^ uncoded_block[1032];
  wire _31173 = _1338 ^ _31172;
  wire _31174 = _2129 ^ _6475;
  wire _31175 = _31173 ^ _31174;
  wire _31176 = _11677 ^ _8309;
  wire _31177 = _2134 ^ _12762;
  wire _31178 = _31176 ^ _31177;
  wire _31179 = _31175 ^ _31178;
  wire _31180 = _31171 ^ _31179;
  wire _31181 = _5816 ^ _2140;
  wire _31182 = _31181 ^ _12769;
  wire _31183 = _2143 ^ _2146;
  wire _31184 = _6486 ^ _5834;
  wire _31185 = _31183 ^ _31184;
  wire _31186 = _31182 ^ _31185;
  wire _31187 = uncoded_block[1083] ^ uncoded_block[1088];
  wire _31188 = _7724 ^ _31187;
  wire _31189 = uncoded_block[1090] ^ uncoded_block[1094];
  wire _31190 = _31189 ^ _8330;
  wire _31191 = _31188 ^ _31190;
  wire _31192 = uncoded_block[1103] ^ uncoded_block[1107];
  wire _31193 = _4444 ^ _31192;
  wire _31194 = _2164 ^ _4451;
  wire _31195 = _31193 ^ _31194;
  wire _31196 = _31191 ^ _31195;
  wire _31197 = _31186 ^ _31196;
  wire _31198 = _31180 ^ _31197;
  wire _31199 = _29869 ^ _9490;
  wire _31200 = _6499 ^ _2174;
  wire _31201 = uncoded_block[1136] ^ uncoded_block[1142];
  wire _31202 = _31201 ^ _5861;
  wire _31203 = _31200 ^ _31202;
  wire _31204 = _31199 ^ _31203;
  wire _31205 = _8354 ^ _5190;
  wire _31206 = _20271 ^ _31205;
  wire _31207 = _1404 ^ _22627;
  wire _31208 = _7151 ^ _11161;
  wire _31209 = _31207 ^ _31208;
  wire _31210 = _31206 ^ _31209;
  wire _31211 = _31204 ^ _31210;
  wire _31212 = _17890 ^ _590;
  wire _31213 = _592 ^ _5201;
  wire _31214 = _31212 ^ _31213;
  wire _31215 = _13346 ^ _1420;
  wire _31216 = _8951 ^ _1424;
  wire _31217 = _31215 ^ _31216;
  wire _31218 = _31214 ^ _31217;
  wire _31219 = uncoded_block[1215] ^ uncoded_block[1219];
  wire _31220 = _10617 ^ _31219;
  wire _31221 = _18394 ^ _31220;
  wire _31222 = _4502 ^ _30773;
  wire _31223 = _31222 ^ _13895;
  wire _31224 = _31221 ^ _31223;
  wire _31225 = _31218 ^ _31224;
  wire _31226 = _31211 ^ _31225;
  wire _31227 = _31198 ^ _31226;
  wire _31228 = uncoded_block[1232] ^ uncoded_block[1233];
  wire _31229 = uncoded_block[1235] ^ uncoded_block[1239];
  wire _31230 = _31228 ^ _31229;
  wire _31231 = uncoded_block[1240] ^ uncoded_block[1243];
  wire _31232 = _31231 ^ _13365;
  wire _31233 = _31230 ^ _31232;
  wire _31234 = _5229 ^ _8385;
  wire _31235 = _5231 ^ _3783;
  wire _31236 = _31234 ^ _31235;
  wire _31237 = _31233 ^ _31236;
  wire _31238 = _24015 ^ _11189;
  wire _31239 = _9538 ^ _5907;
  wire _31240 = _4525 ^ _23124;
  wire _31241 = _31239 ^ _31240;
  wire _31242 = _31238 ^ _31241;
  wire _31243 = _31237 ^ _31242;
  wire _31244 = _3801 ^ _28321;
  wire _31245 = _7187 ^ _31244;
  wire _31246 = _22665 ^ _2259;
  wire _31247 = uncoded_block[1309] ^ uncoded_block[1313];
  wire _31248 = _31247 ^ _3811;
  wire _31249 = _31246 ^ _31248;
  wire _31250 = _31245 ^ _31249;
  wire _31251 = _3814 ^ _8994;
  wire _31252 = _31251 ^ _19849;
  wire _31253 = _2276 ^ _5266;
  wire _31254 = uncoded_block[1349] ^ uncoded_block[1353];
  wire _31255 = _5268 ^ _31254;
  wire _31256 = _31253 ^ _31255;
  wire _31257 = _31252 ^ _31256;
  wire _31258 = _31250 ^ _31257;
  wire _31259 = _31243 ^ _31258;
  wire _31260 = _12857 ^ _5273;
  wire _31261 = _31260 ^ _6590;
  wire _31262 = _9572 ^ _7824;
  wire _31263 = _23151 ^ _31262;
  wire _31264 = _31261 ^ _31263;
  wire _31265 = _687 ^ _17953;
  wire _31266 = _7828 ^ _694;
  wire _31267 = _31265 ^ _31266;
  wire _31268 = _1516 ^ _5293;
  wire _31269 = _3846 ^ _18452;
  wire _31270 = _31268 ^ _31269;
  wire _31271 = _31267 ^ _31270;
  wire _31272 = _31264 ^ _31271;
  wire _31273 = _7229 ^ _704;
  wire _31274 = uncoded_block[1423] ^ uncoded_block[1427];
  wire _31275 = _3072 ^ _31274;
  wire _31276 = _31273 ^ _31275;
  wire _31277 = _30403 ^ _1533;
  wire _31278 = _2314 ^ _24521;
  wire _31279 = _31277 ^ _31278;
  wire _31280 = _31276 ^ _31279;
  wire _31281 = _2319 ^ _2321;
  wire _31282 = _2322 ^ _2325;
  wire _31283 = _31281 ^ _31282;
  wire _31284 = _2326 ^ _6622;
  wire _31285 = _3088 ^ _724;
  wire _31286 = _31284 ^ _31285;
  wire _31287 = _31283 ^ _31286;
  wire _31288 = _31280 ^ _31287;
  wire _31289 = _31272 ^ _31288;
  wire _31290 = _31259 ^ _31289;
  wire _31291 = _31227 ^ _31290;
  wire _31292 = _18919 ^ _9608;
  wire _31293 = _23612 ^ _31292;
  wire _31294 = uncoded_block[1478] ^ uncoded_block[1480];
  wire _31295 = _4603 ^ _31294;
  wire _31296 = _9042 ^ _5321;
  wire _31297 = _31295 ^ _31296;
  wire _31298 = _31293 ^ _31297;
  wire _31299 = _1563 ^ _4610;
  wire _31300 = _747 ^ _7259;
  wire _31301 = _31299 ^ _31300;
  wire _31302 = uncoded_block[1511] ^ uncoded_block[1515];
  wire _31303 = _7262 ^ _31302;
  wire _31304 = _7265 ^ _1579;
  wire _31305 = _31303 ^ _31304;
  wire _31306 = _31301 ^ _31305;
  wire _31307 = _31298 ^ _31306;
  wire _31308 = _13459 ^ _6002;
  wire _31309 = uncoded_block[1534] ^ uncoded_block[1538];
  wire _31310 = _31309 ^ _16010;
  wire _31311 = _31308 ^ _31310;
  wire _31312 = _767 ^ _3131;
  wire _31313 = _13473 ^ _31312;
  wire _31314 = _31311 ^ _31313;
  wire _31315 = _11281 ^ _1597;
  wire _31316 = _7889 ^ _25895;
  wire _31317 = _31315 ^ _31316;
  wire _31318 = _25450 ^ _15535;
  wire _31319 = _5368 ^ _14512;
  wire _31320 = _31318 ^ _31319;
  wire _31321 = _31317 ^ _31320;
  wire _31322 = _31314 ^ _31321;
  wire _31323 = _31307 ^ _31322;
  wire _31324 = _26808 ^ _798;
  wire _31325 = _31324 ^ _2397;
  wire _31326 = _7908 ^ _9094;
  wire _31327 = _31326 ^ _16040;
  wire _31328 = _31325 ^ _31327;
  wire _31329 = uncoded_block[1629] ^ uncoded_block[1635];
  wire _31330 = _31329 ^ _1642;
  wire _31331 = _27651 ^ _816;
  wire _31332 = _31330 ^ _31331;
  wire _31333 = uncoded_block[1649] ^ uncoded_block[1654];
  wire _31334 = _31333 ^ _1653;
  wire _31335 = _6055 ^ _19466;
  wire _31336 = _31334 ^ _31335;
  wire _31337 = _31332 ^ _31336;
  wire _31338 = _31328 ^ _31337;
  wire _31339 = uncoded_block[1674] ^ uncoded_block[1679];
  wire _31340 = _8521 ^ _31339;
  wire _31341 = _23671 ^ _6705;
  wire _31342 = _31340 ^ _31341;
  wire _31343 = uncoded_block[1692] ^ uncoded_block[1699];
  wire _31344 = _7935 ^ _31343;
  wire _31345 = _15063 ^ _2437;
  wire _31346 = _31344 ^ _31345;
  wire _31347 = _31342 ^ _31346;
  wire _31348 = _3200 ^ _2443;
  wire _31349 = _31348 ^ _5416;
  wire _31350 = _31347 ^ _31349;
  wire _31351 = _31338 ^ _31350;
  wire _31352 = _31323 ^ _31351;
  wire _31353 = _31291 ^ _31352;
  wire _31354 = _31164 ^ _31353;
  wire _31355 = _16560 ^ _3212;
  wire _31356 = uncoded_block[9] ^ uncoded_block[15];
  wire _31357 = _31356 ^ _871;
  wire _31358 = _31355 ^ _31357;
  wire _31359 = _13537 ^ _10791;
  wire _31360 = _7959 ^ _9143;
  wire _31361 = _31359 ^ _31360;
  wire _31362 = _31358 ^ _31361;
  wire _31363 = uncoded_block[30] ^ uncoded_block[32];
  wire _31364 = _31363 ^ _6095;
  wire _31365 = uncoded_block[39] ^ uncoded_block[43];
  wire _31366 = _15590 ^ _31365;
  wire _31367 = _31364 ^ _31366;
  wire _31368 = _10234 ^ _3233;
  wire _31369 = _14575 ^ _7969;
  wire _31370 = _31368 ^ _31369;
  wire _31371 = _31367 ^ _31370;
  wire _31372 = _31362 ^ _31371;
  wire _31373 = _13553 ^ _12435;
  wire _31374 = _25950 ^ _1711;
  wire _31375 = _31373 ^ _31374;
  wire _31376 = _4733 ^ _7979;
  wire _31377 = _11364 ^ _2484;
  wire _31378 = _31376 ^ _31377;
  wire _31379 = _31375 ^ _31378;
  wire _31380 = _6116 ^ _4031;
  wire _31381 = _17081 ^ _31380;
  wire _31382 = uncoded_block[109] ^ uncoded_block[113];
  wire _31383 = _1722 ^ _31382;
  wire _31384 = _10816 ^ _16592;
  wire _31385 = _31383 ^ _31384;
  wire _31386 = _31381 ^ _31385;
  wire _31387 = _31379 ^ _31386;
  wire _31388 = _31372 ^ _31387;
  wire _31389 = _4754 ^ _1736;
  wire _31390 = _20483 ^ _31389;
  wire _31391 = _11918 ^ _15114;
  wire _31392 = uncoded_block[145] ^ uncoded_block[149];
  wire _31393 = uncoded_block[150] ^ uncoded_block[153];
  wire _31394 = _31392 ^ _31393;
  wire _31395 = _31391 ^ _31394;
  wire _31396 = _31390 ^ _31395;
  wire _31397 = _30951 ^ _1749;
  wire _31398 = _7398 ^ _31397;
  wire _31399 = _8589 ^ _8591;
  wire _31400 = _938 ^ _6149;
  wire _31401 = _31399 ^ _31400;
  wire _31402 = _31398 ^ _31401;
  wire _31403 = _31396 ^ _31402;
  wire _31404 = _86 ^ _18111;
  wire _31405 = _11934 ^ _31404;
  wire _31406 = _15636 ^ _8019;
  wire _31407 = _31405 ^ _31406;
  wire _31408 = _3291 ^ _4071;
  wire _31409 = _5491 ^ _2543;
  wire _31410 = _31408 ^ _31409;
  wire _31411 = _29225 ^ _10289;
  wire _31412 = _22844 ^ _31411;
  wire _31413 = _31410 ^ _31412;
  wire _31414 = _31407 ^ _31413;
  wire _31415 = _31403 ^ _31414;
  wire _31416 = _31388 ^ _31415;
  wire _31417 = _6824 ^ _113;
  wire _31418 = _31417 ^ _7433;
  wire _31419 = _26000 ^ _7441;
  wire _31420 = _18599 ^ _31419;
  wire _31421 = _31418 ^ _31420;
  wire _31422 = uncoded_block[277] ^ uncoded_block[280];
  wire _31423 = _130 ^ _31422;
  wire _31424 = _988 ^ _11428;
  wire _31425 = _31423 ^ _31424;
  wire _31426 = _9772 ^ _994;
  wire _31427 = _2573 ^ _138;
  wire _31428 = _31426 ^ _31427;
  wire _31429 = _31425 ^ _31428;
  wire _31430 = _31421 ^ _31429;
  wire _31431 = _30111 ^ _4830;
  wire _31432 = _11974 ^ _31431;
  wire _31433 = _22870 ^ _21948;
  wire _31434 = _31432 ^ _31433;
  wire _31435 = _4838 ^ _2593;
  wire _31436 = _31435 ^ _16656;
  wire _31437 = _9790 ^ _15179;
  wire _31438 = _2601 ^ _21497;
  wire _31439 = _31437 ^ _31438;
  wire _31440 = _31436 ^ _31439;
  wire _31441 = _31434 ^ _31440;
  wire _31442 = _31430 ^ _31441;
  wire _31443 = _6866 ^ _7470;
  wire _31444 = _31443 ^ _18628;
  wire _31445 = _8079 ^ _14150;
  wire _31446 = _6876 ^ _9255;
  wire _31447 = _31445 ^ _31446;
  wire _31448 = _31444 ^ _31447;
  wire _31449 = _18633 ^ _9806;
  wire _31450 = _2623 ^ _5559;
  wire _31451 = _31449 ^ _31450;
  wire _31452 = _15697 ^ _3391;
  wire _31453 = _1054 ^ _3396;
  wire _31454 = _31452 ^ _31453;
  wire _31455 = _31451 ^ _31454;
  wire _31456 = _31448 ^ _31455;
  wire _31457 = _1059 ^ _8671;
  wire _31458 = _31457 ^ _15705;
  wire _31459 = uncoded_block[441] ^ uncoded_block[445];
  wire _31460 = _31459 ^ _10356;
  wire _31461 = _24250 ^ _31460;
  wire _31462 = _31458 ^ _31461;
  wire _31463 = _4176 ^ _4883;
  wire _31464 = _31463 ^ _22435;
  wire _31465 = _30155 ^ _14175;
  wire _31466 = _4182 ^ _31465;
  wire _31467 = _31464 ^ _31466;
  wire _31468 = _31462 ^ _31467;
  wire _31469 = _31456 ^ _31468;
  wire _31470 = _31442 ^ _31469;
  wire _31471 = _31416 ^ _31470;
  wire _31472 = _8686 ^ _2657;
  wire _31473 = _1085 ^ _13135;
  wire _31474 = _31472 ^ _31473;
  wire _31475 = _9832 ^ _6919;
  wire _31476 = _31475 ^ _1098;
  wire _31477 = _31474 ^ _31476;
  wire _31478 = _1892 ^ _231;
  wire _31479 = _9295 ^ _20598;
  wire _31480 = _31478 ^ _31479;
  wire _31481 = _3444 ^ _3447;
  wire _31482 = _6931 ^ _1905;
  wire _31483 = _31481 ^ _31482;
  wire _31484 = _31480 ^ _31483;
  wire _31485 = _31477 ^ _31484;
  wire _31486 = _13688 ^ _1909;
  wire _31487 = _6300 ^ _8721;
  wire _31488 = _31486 ^ _31487;
  wire _31489 = _8724 ^ _256;
  wire _31490 = uncoded_block[563] ^ uncoded_block[567];
  wire _31491 = _31490 ^ _3468;
  wire _31492 = _31489 ^ _31491;
  wire _31493 = _31488 ^ _31492;
  wire _31494 = _262 ^ _22012;
  wire _31495 = _4950 ^ _8148;
  wire _31496 = _31494 ^ _31495;
  wire _31497 = _4952 ^ _9332;
  wire _31498 = _3489 ^ _16233;
  wire _31499 = _31497 ^ _31498;
  wire _31500 = _31496 ^ _31499;
  wire _31501 = _31493 ^ _31500;
  wire _31502 = _31485 ^ _31501;
  wire _31503 = _18232 ^ _21098;
  wire _31504 = _31503 ^ _6961;
  wire _31505 = _4246 ^ _7570;
  wire _31506 = uncoded_block[635] ^ uncoded_block[638];
  wire _31507 = _8749 ^ _31506;
  wire _31508 = _31505 ^ _31507;
  wire _31509 = _31504 ^ _31508;
  wire _31510 = _6335 ^ _8751;
  wire _31511 = _6338 ^ _19177;
  wire _31512 = _31510 ^ _31511;
  wire _31513 = _29746 ^ _14239;
  wire _31514 = _31512 ^ _31513;
  wire _31515 = _31509 ^ _31514;
  wire _31516 = _10990 ^ _1177;
  wire _31517 = _31516 ^ _1969;
  wire _31518 = _12636 ^ _325;
  wire _31519 = _4272 ^ _328;
  wire _31520 = _31518 ^ _31519;
  wire _31521 = _31517 ^ _31520;
  wire _31522 = _14249 ^ _20654;
  wire _31523 = _10448 ^ _3535;
  wire _31524 = _31522 ^ _31523;
  wire _31525 = uncoded_block[712] ^ uncoded_block[715];
  wire _31526 = _31525 ^ _17762;
  wire _31527 = _341 ^ _343;
  wire _31528 = _31526 ^ _31527;
  wire _31529 = _31524 ^ _31528;
  wire _31530 = _31521 ^ _31529;
  wire _31531 = _31515 ^ _31530;
  wire _31532 = _31502 ^ _31531;
  wire _31533 = uncoded_block[730] ^ uncoded_block[733];
  wire _31534 = _5693 ^ _31533;
  wire _31535 = _7605 ^ _1996;
  wire _31536 = _31534 ^ _31535;
  wire _31537 = uncoded_block[748] ^ uncoded_block[752];
  wire _31538 = _353 ^ _31537;
  wire _31539 = _7013 ^ _7015;
  wire _31540 = _31538 ^ _31539;
  wire _31541 = _31536 ^ _31540;
  wire _31542 = uncoded_block[768] ^ uncoded_block[773];
  wire _31543 = _13762 ^ _31542;
  wire _31544 = _26141 ^ _31543;
  wire _31545 = uncoded_block[775] ^ uncoded_block[780];
  wire _31546 = _31545 ^ _3570;
  wire _31547 = _8215 ^ _5033;
  wire _31548 = _31546 ^ _31547;
  wire _31549 = _31544 ^ _31548;
  wire _31550 = _31541 ^ _31549;
  wire _31551 = uncoded_block[797] ^ uncoded_block[801];
  wire _31552 = _31551 ^ _386;
  wire _31553 = _18753 ^ _31552;
  wire _31554 = _2806 ^ _2808;
  wire _31555 = _391 ^ _31554;
  wire _31556 = _31553 ^ _31555;
  wire _31557 = _2028 ^ _14802;
  wire _31558 = _23896 ^ _26160;
  wire _31559 = _31557 ^ _31558;
  wire _31560 = _9938 ^ _2815;
  wire _31561 = uncoded_block[845] ^ uncoded_block[853];
  wire _31562 = _31561 ^ _30680;
  wire _31563 = _31560 ^ _31562;
  wire _31564 = _31559 ^ _31563;
  wire _31565 = _31556 ^ _31564;
  wire _31566 = _31550 ^ _31565;
  wire _31567 = _20192 ^ _22541;
  wire _31568 = _416 ^ _6416;
  wire _31569 = _12151 ^ _7062;
  wire _31570 = _31568 ^ _31569;
  wire _31571 = _31567 ^ _31570;
  wire _31572 = _423 ^ _11059;
  wire _31573 = _20701 ^ _4355;
  wire _31574 = _31572 ^ _31573;
  wire _31575 = _5758 ^ _2843;
  wire _31576 = _11062 ^ _3628;
  wire _31577 = _31575 ^ _31576;
  wire _31578 = _31574 ^ _31577;
  wire _31579 = _31571 ^ _31578;
  wire _31580 = _3629 ^ _29379;
  wire _31581 = uncoded_block[934] ^ uncoded_block[937];
  wire _31582 = _18316 ^ _31581;
  wire _31583 = _31580 ^ _31582;
  wire _31584 = _26189 ^ _9975;
  wire _31585 = _8274 ^ _7680;
  wire _31586 = _31584 ^ _31585;
  wire _31587 = _31583 ^ _31586;
  wire _31588 = _4385 ^ _5108;
  wire _31589 = _11649 ^ _471;
  wire _31590 = _31588 ^ _31589;
  wire _31591 = _1317 ^ _23939;
  wire _31592 = _11095 ^ _31591;
  wire _31593 = _31590 ^ _31592;
  wire _31594 = _31587 ^ _31593;
  wire _31595 = _31579 ^ _31594;
  wire _31596 = _31566 ^ _31595;
  wire _31597 = _31532 ^ _31596;
  wire _31598 = _31471 ^ _31597;
  wire _31599 = _2107 ^ _1326;
  wire _31600 = _9445 ^ _31599;
  wire _31601 = _5129 ^ _13283;
  wire _31602 = _2117 ^ _7703;
  wire _31603 = _31601 ^ _31602;
  wire _31604 = _31600 ^ _31603;
  wire _31605 = _5135 ^ _4415;
  wire _31606 = _2898 ^ _1345;
  wire _31607 = _31605 ^ _31606;
  wire _31608 = _1359 ^ _10566;
  wire _31609 = _31176 ^ _31608;
  wire _31610 = _31607 ^ _31609;
  wire _31611 = _31604 ^ _31610;
  wire _31612 = _11681 ^ _11123;
  wire _31613 = _7722 ^ _6486;
  wire _31614 = _31613 ^ _12773;
  wire _31615 = _31612 ^ _31614;
  wire _31616 = _17363 ^ _31189;
  wire _31617 = _543 ^ _11142;
  wire _31618 = _31616 ^ _31617;
  wire _31619 = _4451 ^ _7133;
  wire _31620 = _19312 ^ _31619;
  wire _31621 = _31618 ^ _31620;
  wire _31622 = _31615 ^ _31621;
  wire _31623 = _31611 ^ _31622;
  wire _31624 = _6499 ^ _27526;
  wire _31625 = _31624 ^ _28627;
  wire _31626 = _23082 ^ _31625;
  wire _31627 = _10597 ^ _2956;
  wire _31628 = _10037 ^ _31627;
  wire _31629 = uncoded_block[1160] ^ uncoded_block[1164];
  wire _31630 = _578 ^ _31629;
  wire _31631 = _30336 ^ _31630;
  wire _31632 = _31628 ^ _31631;
  wire _31633 = _31626 ^ _31632;
  wire _31634 = _17390 ^ _10046;
  wire _31635 = _7154 ^ _13339;
  wire _31636 = _31634 ^ _31635;
  wire _31637 = uncoded_block[1177] ^ uncoded_block[1182];
  wire _31638 = _31637 ^ _4486;
  wire _31639 = _31638 ^ _23538;
  wire _31640 = _31636 ^ _31639;
  wire _31641 = _2206 ^ _6529;
  wire _31642 = _1422 ^ _31641;
  wire _31643 = _4498 ^ _3765;
  wire _31644 = _13891 ^ _31643;
  wire _31645 = _31642 ^ _31644;
  wire _31646 = _31640 ^ _31645;
  wire _31647 = _31633 ^ _31646;
  wire _31648 = _31623 ^ _31647;
  wire _31649 = _7168 ^ _1436;
  wire _31650 = _3769 ^ _5219;
  wire _31651 = _31649 ^ _31650;
  wire _31652 = _11181 ^ _4509;
  wire _31653 = uncoded_block[1244] ^ uncoded_block[1250];
  wire _31654 = _31653 ^ _7778;
  wire _31655 = _31652 ^ _31654;
  wire _31656 = _31651 ^ _31655;
  wire _31657 = _2235 ^ _3783;
  wire _31658 = _31657 ^ _24015;
  wire _31659 = _1460 ^ _4524;
  wire _31660 = _31658 ^ _31659;
  wire _31661 = _31656 ^ _31660;
  wire _31662 = _1463 ^ _12837;
  wire _31663 = uncoded_block[1285] ^ uncoded_block[1289];
  wire _31664 = _31663 ^ _1468;
  wire _31665 = _31662 ^ _31664;
  wire _31666 = _12843 ^ _2254;
  wire _31667 = _29064 ^ _31666;
  wire _31668 = _31665 ^ _31667;
  wire _31669 = uncoded_block[1307] ^ uncoded_block[1312];
  wire _31670 = _648 ^ _31669;
  wire _31671 = uncoded_block[1316] ^ uncoded_block[1327];
  wire _31672 = _2261 ^ _31671;
  wire _31673 = _31670 ^ _31672;
  wire _31674 = _1490 ^ _5931;
  wire _31675 = uncoded_block[1336] ^ uncoded_block[1341];
  wire _31676 = uncoded_block[1342] ^ uncoded_block[1346];
  wire _31677 = _31675 ^ _31676;
  wire _31678 = _31674 ^ _31677;
  wire _31679 = _31673 ^ _31678;
  wire _31680 = _31668 ^ _31679;
  wire _31681 = _31661 ^ _31680;
  wire _31682 = _17446 ^ _18437;
  wire _31683 = _5940 ^ _7821;
  wire _31684 = _31683 ^ _11225;
  wire _31685 = _31682 ^ _31684;
  wire _31686 = uncoded_block[1368] ^ uncoded_block[1371];
  wire _31687 = _31686 ^ _9572;
  wire _31688 = _12866 ^ _3059;
  wire _31689 = _31687 ^ _31688;
  wire _31690 = _691 ^ _4569;
  wire _31691 = _31690 ^ _7226;
  wire _31692 = _31689 ^ _31691;
  wire _31693 = _31685 ^ _31692;
  wire _31694 = _5293 ^ _14457;
  wire _31695 = _13420 ^ _7229;
  wire _31696 = _31694 ^ _31695;
  wire _31697 = _704 ^ _5964;
  wire _31698 = uncoded_block[1423] ^ uncoded_block[1428];
  wire _31699 = _31698 ^ _9591;
  wire _31700 = _31697 ^ _31699;
  wire _31701 = _31696 ^ _31700;
  wire _31702 = _2314 ^ _17470;
  wire _31703 = _20355 ^ _5305;
  wire _31704 = _31702 ^ _31703;
  wire _31705 = uncoded_block[1452] ^ uncoded_block[1459];
  wire _31706 = _1543 ^ _31705;
  wire _31707 = _20361 ^ _9602;
  wire _31708 = _31706 ^ _31707;
  wire _31709 = _31704 ^ _31708;
  wire _31710 = _31701 ^ _31709;
  wire _31711 = _31693 ^ _31710;
  wire _31712 = _31681 ^ _31711;
  wire _31713 = _31648 ^ _31712;
  wire _31714 = _31294 ^ _5320;
  wire _31715 = _10702 ^ _31714;
  wire _31716 = _5321 ^ _1563;
  wire _31717 = uncoded_block[1494] ^ uncoded_block[1502];
  wire _31718 = _31717 ^ _7259;
  wire _31719 = _31716 ^ _31718;
  wire _31720 = _31715 ^ _31719;
  wire _31721 = _23624 ^ _31302;
  wire _31722 = _31721 ^ _31304;
  wire _31723 = _3122 ^ _11272;
  wire _31724 = uncoded_block[1531] ^ uncoded_block[1538];
  wire _31725 = _31724 ^ _16010;
  wire _31726 = _31723 ^ _31725;
  wire _31727 = _31722 ^ _31726;
  wire _31728 = _31720 ^ _31727;
  wire _31729 = _16499 ^ _13471;
  wire _31730 = _13472 ^ _3131;
  wire _31731 = _31729 ^ _31730;
  wire _31732 = uncoded_block[1557] ^ uncoded_block[1560];
  wire _31733 = _31732 ^ _2372;
  wire _31734 = _24102 ^ _7892;
  wire _31735 = _31733 ^ _31734;
  wire _31736 = _31731 ^ _31735;
  wire _31737 = _784 ^ _9083;
  wire _31738 = _24565 ^ _3934;
  wire _31739 = _31737 ^ _31738;
  wire _31740 = uncoded_block[1608] ^ uncoded_block[1611];
  wire _31741 = _800 ^ _31740;
  wire _31742 = _10739 ^ _31741;
  wire _31743 = _31739 ^ _31742;
  wire _31744 = _31736 ^ _31743;
  wire _31745 = _31728 ^ _31744;
  wire _31746 = uncoded_block[1622] ^ uncoded_block[1624];
  wire _31747 = _31746 ^ _12947;
  wire _31748 = _18021 ^ _31747;
  wire _31749 = uncoded_block[1628] ^ uncoded_block[1631];
  wire _31750 = _31749 ^ _7914;
  wire _31751 = _31750 ^ _15556;
  wire _31752 = _31748 ^ _31751;
  wire _31753 = _27651 ^ _5394;
  wire _31754 = _6691 ^ _17529;
  wire _31755 = _31753 ^ _31754;
  wire _31756 = _12957 ^ _29569;
  wire _31757 = _16049 ^ _5399;
  wire _31758 = _31756 ^ _31757;
  wire _31759 = _31755 ^ _31758;
  wire _31760 = _31752 ^ _31759;
  wire _31761 = _7928 ^ _6059;
  wire _31762 = _11321 ^ _4691;
  wire _31763 = _31761 ^ _31762;
  wire _31764 = _4693 ^ _6705;
  wire _31765 = _31764 ^ _29576;
  wire _31766 = _31763 ^ _31765;
  wire _31767 = _24137 ^ _15063;
  wire _31768 = _31767 ^ _2439;
  wire _31769 = _31348 ^ uncoded_block[1720];
  wire _31770 = _31768 ^ _31769;
  wire _31771 = _31766 ^ _31770;
  wire _31772 = _31760 ^ _31771;
  wire _31773 = _31745 ^ _31772;
  wire _31774 = _31713 ^ _31773;
  wire _31775 = _31598 ^ _31774;
  wire _31776 = _3993 ^ _4713;
  wire _31777 = _4711 ^ _31776;
  wire _31778 = _5423 ^ _4716;
  wire _31779 = _10 ^ _6093;
  wire _31780 = _31778 ^ _31779;
  wire _31781 = _31777 ^ _31780;
  wire _31782 = _875 ^ _8549;
  wire _31783 = _19 ^ _20457;
  wire _31784 = _31782 ^ _31783;
  wire _31785 = _15594 ^ _9150;
  wire _31786 = _5436 ^ _1703;
  wire _31787 = _31785 ^ _31786;
  wire _31788 = _31784 ^ _31787;
  wire _31789 = _31781 ^ _31788;
  wire _31790 = uncoded_block[59] ^ uncoded_block[63];
  wire _31791 = _31790 ^ _12435;
  wire _31792 = _31791 ^ _6746;
  wire _31793 = _4733 ^ _6109;
  wire _31794 = _31793 ^ _4736;
  wire _31795 = _31792 ^ _31794;
  wire _31796 = _17578 ^ _6113;
  wire _31797 = _31796 ^ _9165;
  wire _31798 = _7377 ^ _7986;
  wire _31799 = _17584 ^ _8572;
  wire _31800 = _31798 ^ _31799;
  wire _31801 = _31797 ^ _31800;
  wire _31802 = _31795 ^ _31801;
  wire _31803 = _31789 ^ _31802;
  wire _31804 = _6769 ^ _10819;
  wire _31805 = _10821 ^ _25073;
  wire _31806 = _31804 ^ _31805;
  wire _31807 = _924 ^ _22819;
  wire _31808 = _7999 ^ _17097;
  wire _31809 = _31807 ^ _31808;
  wire _31810 = _31806 ^ _31809;
  wire _31811 = _27279 ^ _22827;
  wire _31812 = _6785 ^ _79;
  wire _31813 = uncoded_block[171] ^ uncoded_block[174];
  wire _31814 = _31813 ^ _82;
  wire _31815 = _31812 ^ _31814;
  wire _31816 = _31811 ^ _31815;
  wire _31817 = _31810 ^ _31816;
  wire _31818 = _1759 ^ _13588;
  wire _31819 = _20981 ^ _31818;
  wire _31820 = _2532 ^ _8018;
  wire _31821 = _10852 ^ _956;
  wire _31822 = _31820 ^ _31821;
  wire _31823 = _31819 ^ _31822;
  wire _31824 = _8606 ^ _5492;
  wire _31825 = _5497 ^ _20990;
  wire _31826 = _31824 ^ _31825;
  wire _31827 = _1778 ^ _21465;
  wire _31828 = _6180 ^ _2556;
  wire _31829 = _31827 ^ _31828;
  wire _31830 = _31826 ^ _31829;
  wire _31831 = _31823 ^ _31830;
  wire _31832 = _31817 ^ _31831;
  wire _31833 = _31803 ^ _31832;
  wire _31834 = uncoded_block[252] ^ uncoded_block[255];
  wire _31835 = _31834 ^ _1788;
  wire _31836 = _120 ^ _6188;
  wire _31837 = _31835 ^ _31836;
  wire _31838 = uncoded_block[268] ^ uncoded_block[273];
  wire _31839 = _31838 ^ _5515;
  wire _31840 = _31839 ^ _18138;
  wire _31841 = _31837 ^ _31840;
  wire _31842 = uncoded_block[289] ^ uncoded_block[293];
  wire _31843 = uncoded_block[294] ^ uncoded_block[298];
  wire _31844 = _31842 ^ _31843;
  wire _31845 = _29656 ^ _1000;
  wire _31846 = _31844 ^ _31845;
  wire _31847 = uncoded_block[306] ^ uncoded_block[309];
  wire _31848 = _31847 ^ _8056;
  wire _31849 = _17642 ^ _1008;
  wire _31850 = _31848 ^ _31849;
  wire _31851 = _31846 ^ _31850;
  wire _31852 = _31841 ^ _31851;
  wire _31853 = _13625 ^ _8058;
  wire _31854 = _4125 ^ _1017;
  wire _31855 = _31853 ^ _31854;
  wire _31856 = _4840 ^ _6218;
  wire _31857 = _4844 ^ _11454;
  wire _31858 = _31856 ^ _31857;
  wire _31859 = _31855 ^ _31858;
  wire _31860 = _1833 ^ _6228;
  wire _31861 = _31860 ^ _6230;
  wire _31862 = uncoded_block[370] ^ uncoded_block[373];
  wire _31863 = uncoded_block[374] ^ uncoded_block[380];
  wire _31864 = _31862 ^ _31863;
  wire _31865 = _28090 ^ _12541;
  wire _31866 = _31864 ^ _31865;
  wire _31867 = _31861 ^ _31866;
  wire _31868 = _31859 ^ _31867;
  wire _31869 = _31852 ^ _31868;
  wire _31870 = uncoded_block[395] ^ uncoded_block[397];
  wire _31871 = _31870 ^ _25141;
  wire _31872 = _4867 ^ _11473;
  wire _31873 = _31871 ^ _31872;
  wire _31874 = _1060 ^ _9271;
  wire _31875 = _10346 ^ _31874;
  wire _31876 = _31873 ^ _31875;
  wire _31877 = _7497 ^ _205;
  wire _31878 = uncoded_block[447] ^ uncoded_block[453];
  wire _31879 = _1864 ^ _31878;
  wire _31880 = _31877 ^ _31879;
  wire _31881 = _215 ^ _1079;
  wire _31882 = _24257 ^ _31881;
  wire _31883 = _31880 ^ _31882;
  wire _31884 = _31876 ^ _31883;
  wire _31885 = _3418 ^ _7509;
  wire _31886 = _2657 ^ _1086;
  wire _31887 = _31885 ^ _31886;
  wire _31888 = _1090 ^ _2664;
  wire _31889 = _7520 ^ _5607;
  wire _31890 = _31888 ^ _31889;
  wire _31891 = _31887 ^ _31890;
  wire _31892 = _30605 ^ _8122;
  wire _31893 = _236 ^ _1898;
  wire _31894 = _31892 ^ _31893;
  wire _31895 = _4921 ^ _14716;
  wire _31896 = _10384 ^ _1905;
  wire _31897 = _31895 ^ _31896;
  wire _31898 = _31894 ^ _31897;
  wire _31899 = _31891 ^ _31898;
  wire _31900 = _31884 ^ _31899;
  wire _31901 = _31869 ^ _31900;
  wire _31902 = _31833 ^ _31901;
  wire _31903 = _3451 ^ _1909;
  wire _31904 = uncoded_block[549] ^ uncoded_block[551];
  wire _31905 = _31904 ^ _8721;
  wire _31906 = _31903 ^ _31905;
  wire _31907 = uncoded_block[559] ^ uncoded_block[562];
  wire _31908 = _15740 ^ _31907;
  wire _31909 = uncoded_block[564] ^ uncoded_block[568];
  wire _31910 = _31909 ^ _6942;
  wire _31911 = _31908 ^ _31910;
  wire _31912 = _31906 ^ _31911;
  wire _31913 = _4224 ^ _18684;
  wire _31914 = _31913 ^ _28513;
  wire _31915 = uncoded_block[583] ^ uncoded_block[586];
  wire _31916 = _31915 ^ _271;
  wire _31917 = _25640 ^ _3487;
  wire _31918 = _31916 ^ _31917;
  wire _31919 = _31914 ^ _31918;
  wire _31920 = _31912 ^ _31919;
  wire _31921 = _2710 ^ _4242;
  wire _31922 = _7564 ^ _13713;
  wire _31923 = _31921 ^ _31922;
  wire _31924 = uncoded_block[621] ^ uncoded_block[626];
  wire _31925 = _4960 ^ _31924;
  wire _31926 = _17238 ^ _14228;
  wire _31927 = _31925 ^ _31926;
  wire _31928 = _31923 ^ _31927;
  wire _31929 = uncoded_block[639] ^ uncoded_block[643];
  wire _31930 = _6331 ^ _31929;
  wire _31931 = _31930 ^ _2731;
  wire _31932 = _20134 ^ _3513;
  wire _31933 = _15768 ^ _7586;
  wire _31934 = _31932 ^ _31933;
  wire _31935 = _31931 ^ _31934;
  wire _31936 = _31928 ^ _31935;
  wire _31937 = _31920 ^ _31936;
  wire _31938 = _15775 ^ _8177;
  wire _31939 = _6352 ^ _18247;
  wire _31940 = _31938 ^ _31939;
  wire _31941 = _2751 ^ _11556;
  wire _31942 = _17752 ^ _31941;
  wire _31943 = _31940 ^ _31942;
  wire _31944 = _333 ^ _3533;
  wire _31945 = _15285 ^ _31944;
  wire _31946 = _1192 ^ _3536;
  wire _31947 = _18726 ^ _4283;
  wire _31948 = _31946 ^ _31947;
  wire _31949 = _31945 ^ _31948;
  wire _31950 = _31943 ^ _31949;
  wire _31951 = _11006 ^ _7002;
  wire _31952 = uncoded_block[734] ^ uncoded_block[740];
  wire _31953 = _31952 ^ _17272;
  wire _31954 = _31951 ^ _31953;
  wire _31955 = _5013 ^ _24331;
  wire _31956 = _2778 ^ _23879;
  wire _31957 = _31955 ^ _31956;
  wire _31958 = _31954 ^ _31957;
  wire _31959 = _8781 ^ _13215;
  wire _31960 = _7019 ^ _3567;
  wire _31961 = _31959 ^ _31960;
  wire _31962 = _2015 ^ _3570;
  wire _31963 = uncoded_block[786] ^ uncoded_block[791];
  wire _31964 = _31963 ^ _1232;
  wire _31965 = _31962 ^ _31964;
  wire _31966 = _31961 ^ _31965;
  wire _31967 = _31958 ^ _31966;
  wire _31968 = _31950 ^ _31967;
  wire _31969 = _31937 ^ _31968;
  wire _31970 = _11591 ^ _16790;
  wire _31971 = uncoded_block[814] ^ uncoded_block[818];
  wire _31972 = _15318 ^ _31971;
  wire _31973 = _31970 ^ _31972;
  wire _31974 = _397 ^ _4331;
  wire _31975 = _31974 ^ _25250;
  wire _31976 = _31973 ^ _31975;
  wire _31977 = _4339 ^ _1257;
  wire _31978 = _25711 ^ _7049;
  wire _31979 = _31977 ^ _31978;
  wire _31980 = _6410 ^ _29800;
  wire _31981 = _5071 ^ _2830;
  wire _31982 = _31980 ^ _31981;
  wire _31983 = _31979 ^ _31982;
  wire _31984 = _31976 ^ _31983;
  wire _31985 = _417 ^ _3608;
  wire _31986 = _5079 ^ _2058;
  wire _31987 = _31985 ^ _31986;
  wire _31988 = uncoded_block[896] ^ uncoded_block[902];
  wire _31989 = _24367 ^ _31988;
  wire _31990 = _9961 ^ _16312;
  wire _31991 = _31989 ^ _31990;
  wire _31992 = _31987 ^ _31991;
  wire _31993 = _1287 ^ _21644;
  wire _31994 = _31993 ^ _3633;
  wire _31995 = uncoded_block[923] ^ uncoded_block[925];
  wire _31996 = _31995 ^ _4371;
  wire _31997 = uncoded_block[930] ^ uncoded_block[936];
  wire _31998 = _31997 ^ _4375;
  wire _31999 = _31996 ^ _31998;
  wire _32000 = _31994 ^ _31999;
  wire _32001 = _31992 ^ _32000;
  wire _32002 = _31984 ^ _32001;
  wire _32003 = _13263 ^ _456;
  wire _32004 = _32003 ^ _9436;
  wire _32005 = _22564 ^ _4385;
  wire _32006 = _1310 ^ _2092;
  wire _32007 = _32005 ^ _32006;
  wire _32008 = _32004 ^ _32007;
  wire _32009 = uncoded_block[971] ^ uncoded_block[974];
  wire _32010 = _6447 ^ _32009;
  wire _32011 = _11091 ^ _2100;
  wire _32012 = _32010 ^ _32011;
  wire _32013 = _8855 ^ _12186;
  wire _32014 = _32013 ^ _28601;
  wire _32015 = _32012 ^ _32014;
  wire _32016 = _32008 ^ _32015;
  wire _32017 = _29835 ^ _28241;
  wire _32018 = _20730 ^ _13282;
  wire _32019 = _32017 ^ _32018;
  wire _32020 = _492 ^ _9998;
  wire _32021 = _20228 ^ _32020;
  wire _32022 = _32019 ^ _32021;
  wire _32023 = _28995 ^ _8306;
  wire _32024 = _15866 ^ _32023;
  wire _32025 = _2914 ^ _519;
  wire _32026 = _5815 ^ _32025;
  wire _32027 = _32024 ^ _32026;
  wire _32028 = _32022 ^ _32027;
  wire _32029 = _32016 ^ _32028;
  wire _32030 = _32002 ^ _32029;
  wire _32031 = _31969 ^ _32030;
  wire _32032 = _31902 ^ _32031;
  wire _32033 = _13849 ^ _14357;
  wire _32034 = _32033 ^ _11123;
  wire _32035 = uncoded_block[1072] ^ uncoded_block[1077];
  wire _32036 = _32035 ^ _5162;
  wire _32037 = _7724 ^ _534;
  wire _32038 = _32036 ^ _32037;
  wire _32039 = _32034 ^ _32038;
  wire _32040 = _8906 ^ _537;
  wire _32041 = _32040 ^ _11140;
  wire _32042 = uncoded_block[1106] ^ uncoded_block[1110];
  wire _32043 = _2160 ^ _32042;
  wire _32044 = _2938 ^ _1388;
  wire _32045 = _32043 ^ _32044;
  wire _32046 = _32041 ^ _32045;
  wire _32047 = _32039 ^ _32046;
  wire _32048 = _3714 ^ _557;
  wire _32049 = _12791 ^ _8343;
  wire _32050 = _32048 ^ _32049;
  wire _32051 = _1393 ^ _15896;
  wire _32052 = _20266 ^ _8930;
  wire _32053 = _32051 ^ _32052;
  wire _32054 = _32050 ^ _32053;
  wire _32055 = _2179 ^ _5184;
  wire _32056 = uncoded_block[1152] ^ uncoded_block[1155];
  wire _32057 = _4466 ^ _32056;
  wire _32058 = _32055 ^ _32057;
  wire _32059 = _3728 ^ _29028;
  wire _32060 = _32059 ^ _16897;
  wire _32061 = _32058 ^ _32060;
  wire _32062 = _32054 ^ _32061;
  wire _32063 = _32047 ^ _32062;
  wire _32064 = uncoded_block[1172] ^ uncoded_block[1176];
  wire _32065 = _1408 ^ _32064;
  wire _32066 = _589 ^ _3742;
  wire _32067 = _32065 ^ _32066;
  wire _32068 = _16902 ^ _28637;
  wire _32069 = _32067 ^ _32068;
  wire _32070 = _13347 ^ _7758;
  wire _32071 = _1425 ^ _2217;
  wire _32072 = _32070 ^ _32071;
  wire _32073 = _1428 ^ _2982;
  wire _32074 = _3763 ^ _5215;
  wire _32075 = _32073 ^ _32074;
  wire _32076 = _32072 ^ _32075;
  wire _32077 = _32069 ^ _32076;
  wire _32078 = _5891 ^ _11180;
  wire _32079 = _3771 ^ _11734;
  wire _32080 = _32078 ^ _32079;
  wire _32081 = _2997 ^ _5901;
  wire _32082 = uncoded_block[1255] ^ uncoded_block[1257];
  wire _32083 = _32082 ^ _3003;
  wire _32084 = _32081 ^ _32083;
  wire _32085 = _32080 ^ _32084;
  wire _32086 = _13371 ^ _22656;
  wire _32087 = _10638 ^ _29472;
  wire _32088 = _7797 ^ _30797;
  wire _32089 = _32087 ^ _32088;
  wire _32090 = _32086 ^ _32089;
  wire _32091 = _32085 ^ _32090;
  wire _32092 = _32077 ^ _32091;
  wire _32093 = _32063 ^ _32092;
  wire _32094 = _3015 ^ _18870;
  wire _32095 = _2254 ^ _2259;
  wire _32096 = _32094 ^ _32095;
  wire _32097 = _1480 ^ _20314;
  wire _32098 = _9555 ^ _8411;
  wire _32099 = _32097 ^ _32098;
  wire _32100 = _32096 ^ _32099;
  wire _32101 = _14437 ^ _7814;
  wire _32102 = uncoded_block[1344] ^ uncoded_block[1350];
  wire _32103 = _7815 ^ _32102;
  wire _32104 = _32101 ^ _32103;
  wire _32105 = _670 ^ _12857;
  wire _32106 = uncoded_block[1360] ^ uncoded_block[1366];
  wire _32107 = _32106 ^ _11226;
  wire _32108 = _32105 ^ _32107;
  wire _32109 = _32104 ^ _32108;
  wire _32110 = _32100 ^ _32109;
  wire _32111 = _12305 ^ _4564;
  wire _32112 = _10108 ^ _7222;
  wire _32113 = _32111 ^ _32112;
  wire _32114 = _2293 ^ _20340;
  wire _32115 = _3066 ^ _26749;
  wire _32116 = _32114 ^ _32115;
  wire _32117 = _32113 ^ _32116;
  wire _32118 = _701 ^ _7229;
  wire _32119 = _20347 ^ _705;
  wire _32120 = _32118 ^ _32119;
  wire _32121 = _10120 ^ _2308;
  wire _32122 = _2311 ^ _18459;
  wire _32123 = _32121 ^ _32122;
  wire _32124 = _32120 ^ _32123;
  wire _32125 = _32117 ^ _32124;
  wire _32126 = _32110 ^ _32125;
  wire _32127 = _17470 ^ _4590;
  wire _32128 = _3084 ^ _3864;
  wire _32129 = _32127 ^ _32128;
  wire _32130 = uncoded_block[1454] ^ uncoded_block[1460];
  wire _32131 = _16970 ^ _32130;
  wire _32132 = _3871 ^ _10136;
  wire _32133 = _32131 ^ _32132;
  wire _32134 = _32129 ^ _32133;
  wire _32135 = _733 ^ _735;
  wire _32136 = _12889 ^ _32135;
  wire _32137 = _15994 ^ _1562;
  wire _32138 = _9044 ^ _7864;
  wire _32139 = _32137 ^ _32138;
  wire _32140 = _32136 ^ _32139;
  wire _32141 = _32134 ^ _32140;
  wire _32142 = _3112 ^ _5333;
  wire _32143 = _10144 ^ _32142;
  wire _32144 = _13458 ^ _3900;
  wire _32145 = _29971 ^ _32144;
  wire _32146 = _32143 ^ _32145;
  wire _32147 = _6001 ^ _16008;
  wire _32148 = _5348 ^ _6008;
  wire _32149 = _32147 ^ _32148;
  wire _32150 = uncoded_block[1549] ^ uncoded_block[1553];
  wire _32151 = _32150 ^ _22731;
  wire _32152 = _4635 ^ _32151;
  wire _32153 = _32149 ^ _32152;
  wire _32154 = _32146 ^ _32153;
  wire _32155 = _32141 ^ _32154;
  wire _32156 = _32126 ^ _32155;
  wire _32157 = _32093 ^ _32156;
  wire _32158 = _774 ^ _2376;
  wire _32159 = _11284 ^ _2377;
  wire _32160 = _32158 ^ _32159;
  wire _32161 = _2379 ^ _3920;
  wire _32162 = uncoded_block[1580] ^ uncoded_block[1584];
  wire _32163 = _32162 ^ _2386;
  wire _32164 = _32161 ^ _32163;
  wire _32165 = _32160 ^ _32164;
  wire _32166 = _14512 ^ _792;
  wire _32167 = _17012 ^ _32166;
  wire _32168 = _1620 ^ _3936;
  wire _32169 = _32168 ^ _20896;
  wire _32170 = _32167 ^ _32169;
  wire _32171 = _32165 ^ _32170;
  wire _32172 = _18020 ^ _3941;
  wire _32173 = _4665 ^ _4667;
  wire _32174 = _32172 ^ _32173;
  wire _32175 = _7306 ^ _3948;
  wire _32176 = _32175 ^ _26351;
  wire _32177 = _32174 ^ _32176;
  wire _32178 = uncoded_block[1651] ^ uncoded_block[1653];
  wire _32179 = _10757 ^ _32178;
  wire _32180 = _10761 ^ _3175;
  wire _32181 = _32179 ^ _32180;
  wire _32182 = _8522 ^ _10766;
  wire _32183 = _18976 ^ _32182;
  wire _32184 = _32181 ^ _32183;
  wire _32185 = _32177 ^ _32184;
  wire _32186 = _32171 ^ _32185;
  wire _32187 = uncoded_block[1682] ^ uncoded_block[1689];
  wire _32188 = _32187 ^ _7331;
  wire _32189 = uncoded_block[1694] ^ uncoded_block[1699];
  wire _32190 = _9675 ^ _32189;
  wire _32191 = _32188 ^ _32190;
  wire _32192 = _20436 ^ _2438;
  wire _32193 = uncoded_block[1716] ^ uncoded_block[1721];
  wire _32194 = _11333 ^ _32193;
  wire _32195 = _32192 ^ _32194;
  wire _32196 = _32191 ^ _32195;
  wire _32197 = _32196 ^ uncoded_block[1722];
  wire _32198 = _32186 ^ _32197;
  wire _32199 = _32157 ^ _32198;
  wire _32200 = _32032 ^ _32199;
  wire _32201 = uncoded_block[4] ^ uncoded_block[6];
  wire _32202 = _3209 ^ _32201;
  wire _32203 = _6724 ^ _7;
  wire _32204 = _32202 ^ _32203;
  wire _32205 = _19496 ^ _3220;
  wire _32206 = _7352 ^ _32205;
  wire _32207 = _32204 ^ _32206;
  wire _32208 = _6728 ^ _14569;
  wire _32209 = _880 ^ _882;
  wire _32210 = _32208 ^ _32209;
  wire _32211 = uncoded_block[44] ^ uncoded_block[48];
  wire _32212 = uncoded_block[49] ^ uncoded_block[53];
  wire _32213 = _32211 ^ _32212;
  wire _32214 = _7969 ^ _1705;
  wire _32215 = _32213 ^ _32214;
  wire _32216 = _32210 ^ _32215;
  wire _32217 = _32207 ^ _32216;
  wire _32218 = _7367 ^ _30051;
  wire _32219 = _25957 ^ _1718;
  wire _32220 = _32218 ^ _32219;
  wire _32221 = _20952 ^ _21429;
  wire _32222 = _6120 ^ _6122;
  wire _32223 = _32221 ^ _32222;
  wire _32224 = _32220 ^ _32223;
  wire _32225 = _2491 ^ _6763;
  wire _32226 = _6769 ^ _2497;
  wire _32227 = _32225 ^ _32226;
  wire _32228 = _15613 ^ _25523;
  wire _32229 = _32227 ^ _32228;
  wire _32230 = _32224 ^ _32229;
  wire _32231 = _32217 ^ _32230;
  wire _32232 = uncoded_block[134] ^ uncoded_block[140];
  wire _32233 = _21898 ^ _32232;
  wire _32234 = _5461 ^ _24178;
  wire _32235 = _32233 ^ _32234;
  wire _32236 = uncoded_block[150] ^ uncoded_block[154];
  wire _32237 = _6780 ^ _32236;
  wire _32238 = _932 ^ _15118;
  wire _32239 = _32237 ^ _32238;
  wire _32240 = _32235 ^ _32239;
  wire _32241 = _10838 ^ _2523;
  wire _32242 = _6794 ^ _86;
  wire _32243 = _13588 ^ _20500;
  wire _32244 = _32242 ^ _32243;
  wire _32245 = _32241 ^ _32244;
  wire _32246 = _32240 ^ _32245;
  wire _32247 = _94 ^ _6801;
  wire _32248 = uncoded_block[200] ^ uncoded_block[203];
  wire _32249 = _32248 ^ _4070;
  wire _32250 = _32247 ^ _32249;
  wire _32251 = uncoded_block[216] ^ uncoded_block[224];
  wire _32252 = _2540 ^ _32251;
  wire _32253 = _14102 ^ _32252;
  wire _32254 = _32250 ^ _32253;
  wire _32255 = _967 ^ _9208;
  wire _32256 = _12488 ^ _32255;
  wire _32257 = _2552 ^ _10860;
  wire _32258 = _11952 ^ _116;
  wire _32259 = _32257 ^ _32258;
  wire _32260 = _32256 ^ _32259;
  wire _32261 = _32254 ^ _32260;
  wire _32262 = _32246 ^ _32261;
  wire _32263 = _32231 ^ _32262;
  wire _32264 = _4095 ^ _4099;
  wire _32265 = _22385 ^ _32264;
  wire _32266 = _6192 ^ _5515;
  wire _32267 = _11424 ^ _5522;
  wire _32268 = _32266 ^ _32267;
  wire _32269 = _32265 ^ _32268;
  wire _32270 = _9226 ^ _995;
  wire _32271 = _7452 ^ _143;
  wire _32272 = _32270 ^ _32271;
  wire _32273 = _13074 ^ _15670;
  wire _32274 = uncoded_block[314] ^ uncoded_block[319];
  wire _32275 = _32274 ^ _30117;
  wire _32276 = _32273 ^ _32275;
  wire _32277 = _32272 ^ _32276;
  wire _32278 = _32269 ^ _32277;
  wire _32279 = _20547 ^ _3359;
  wire _32280 = _8647 ^ _32279;
  wire _32281 = _3362 ^ _10331;
  wire _32282 = _22878 ^ _32281;
  wire _32283 = _32280 ^ _32282;
  wire _32284 = _13093 ^ _27334;
  wire _32285 = _32284 ^ _7477;
  wire _32286 = _16169 ^ _176;
  wire _32287 = _2616 ^ _1048;
  wire _32288 = _32286 ^ _32287;
  wire _32289 = _32285 ^ _32288;
  wire _32290 = _32283 ^ _32289;
  wire _32291 = _32278 ^ _32290;
  wire _32292 = _26045 ^ _1054;
  wire _32293 = _20565 ^ _32292;
  wire _32294 = _1055 ^ _15197;
  wire _32295 = _32294 ^ _21045;
  wire _32296 = _32293 ^ _32295;
  wire _32297 = uncoded_block[429] ^ uncoded_block[433];
  wire _32298 = _32297 ^ _201;
  wire _32299 = _32298 ^ _21973;
  wire _32300 = _15709 ^ _1866;
  wire _32301 = _1867 ^ _3415;
  wire _32302 = _32300 ^ _32301;
  wire _32303 = _32299 ^ _32302;
  wire _32304 = _32296 ^ _32303;
  wire _32305 = uncoded_block[468] ^ uncoded_block[475];
  wire _32306 = _32305 ^ _8688;
  wire _32307 = _26062 ^ _32306;
  wire _32308 = _5593 ^ _15212;
  wire _32309 = uncoded_block[485] ^ uncoded_block[490];
  wire _32310 = _32309 ^ _6277;
  wire _32311 = _32308 ^ _32310;
  wire _32312 = _32307 ^ _32311;
  wire _32313 = _19135 ^ _2671;
  wire _32314 = _7529 ^ _27369;
  wire _32315 = _32313 ^ _32314;
  wire _32316 = _17702 ^ _31038;
  wire _32317 = _32316 ^ _24737;
  wire _32318 = _32315 ^ _32317;
  wire _32319 = _32312 ^ _32318;
  wire _32320 = _32304 ^ _32319;
  wire _32321 = _32291 ^ _32320;
  wire _32322 = _32263 ^ _32321;
  wire _32323 = _28879 ^ _6292;
  wire _32324 = uncoded_block[541] ^ uncoded_block[546];
  wire _32325 = _32324 ^ _23382;
  wire _32326 = _32323 ^ _32325;
  wire _32327 = uncoded_block[564] ^ uncoded_block[566];
  wire _32328 = _9319 ^ _32327;
  wire _32329 = _19152 ^ _32328;
  wire _32330 = _32326 ^ _32329;
  wire _32331 = _13697 ^ _4224;
  wire _32332 = _18684 ^ _1933;
  wire _32333 = _32331 ^ _32332;
  wire _32334 = _6316 ^ _3487;
  wire _32335 = _4951 ^ _32334;
  wire _32336 = _32333 ^ _32335;
  wire _32337 = _32330 ^ _32336;
  wire _32338 = _1146 ^ _1149;
  wire _32339 = _281 ^ _3495;
  wire _32340 = _32338 ^ _32339;
  wire _32341 = _8161 ^ _5661;
  wire _32342 = _12619 ^ _32341;
  wire _32343 = _32340 ^ _32342;
  wire _32344 = uncoded_block[641] ^ uncoded_block[647];
  wire _32345 = _11543 ^ _32344;
  wire _32346 = _3507 ^ _19674;
  wire _32347 = _32345 ^ _32346;
  wire _32348 = _9885 ^ _15275;
  wire _32349 = _2748 ^ _1968;
  wire _32350 = _32348 ^ _32349;
  wire _32351 = _32347 ^ _32350;
  wire _32352 = _32343 ^ _32351;
  wire _32353 = _32337 ^ _32352;
  wire _32354 = _1971 ^ _10442;
  wire _32355 = _11556 ^ _8186;
  wire _32356 = _32354 ^ _32355;
  wire _32357 = _6360 ^ _10447;
  wire _32358 = _16761 ^ _2762;
  wire _32359 = _32357 ^ _32358;
  wire _32360 = _32356 ^ _32359;
  wire _32361 = _19201 ^ _340;
  wire _32362 = _32361 ^ _24324;
  wire _32363 = _1988 ^ _4286;
  wire _32364 = _30651 ^ _1995;
  wire _32365 = _32363 ^ _32364;
  wire _32366 = _32362 ^ _32365;
  wire _32367 = _32360 ^ _32366;
  wire _32368 = _5699 ^ _2775;
  wire _32369 = uncoded_block[752] ^ uncoded_block[759];
  wire _32370 = _1210 ^ _32369;
  wire _32371 = _32368 ^ _32370;
  wire _32372 = uncoded_block[760] ^ uncoded_block[765];
  wire _32373 = _32372 ^ _17776;
  wire _32374 = _1221 ^ _2792;
  wire _32375 = _32373 ^ _32374;
  wire _32376 = _32371 ^ _32375;
  wire _32377 = _3567 ^ _2015;
  wire _32378 = _14793 ^ _5032;
  wire _32379 = _32377 ^ _32378;
  wire _32380 = _1225 ^ _6391;
  wire _32381 = uncoded_block[802] ^ uncoded_block[808];
  wire _32382 = _7628 ^ _32381;
  wire _32383 = _32380 ^ _32382;
  wire _32384 = _32379 ^ _32383;
  wire _32385 = _32376 ^ _32384;
  wire _32386 = _32367 ^ _32385;
  wire _32387 = _32353 ^ _32386;
  wire _32388 = uncoded_block[815] ^ uncoded_block[819];
  wire _32389 = _11029 ^ _32388;
  wire _32390 = _32389 ^ _5053;
  wire _32391 = _400 ^ _13781;
  wire _32392 = _2035 ^ _1254;
  wire _32393 = _32391 ^ _32392;
  wire _32394 = _32390 ^ _32393;
  wire _32395 = _5058 ^ _3597;
  wire _32396 = _2820 ^ _12146;
  wire _32397 = _32395 ^ _32396;
  wire _32398 = _3600 ^ _20692;
  wire _32399 = _13244 ^ _7054;
  wire _32400 = _32398 ^ _32399;
  wire _32401 = _32397 ^ _32400;
  wire _32402 = _32394 ^ _32401;
  wire _32403 = _1269 ^ _2835;
  wire _32404 = uncoded_block[887] ^ uncoded_block[896];
  wire _32405 = _8820 ^ _32404;
  wire _32406 = _32403 ^ _32405;
  wire _32407 = _2843 ^ _8254;
  wire _32408 = _3623 ^ _30270;
  wire _32409 = _32407 ^ _32408;
  wire _32410 = _32406 ^ _32409;
  wire _32411 = uncoded_block[916] ^ uncoded_block[922];
  wire _32412 = _32411 ^ _5766;
  wire _32413 = _24377 ^ _2858;
  wire _32414 = _32412 ^ _32413;
  wire _32415 = uncoded_block[946] ^ uncoded_block[950];
  wire _32416 = _1300 ^ _32415;
  wire _32417 = _26627 ^ _32416;
  wire _32418 = _32414 ^ _32417;
  wire _32419 = _32410 ^ _32418;
  wire _32420 = _32402 ^ _32419;
  wire _32421 = _9437 ^ _1308;
  wire _32422 = uncoded_block[963] ^ uncoded_block[966];
  wire _32423 = _10529 ^ _32422;
  wire _32424 = _32421 ^ _32423;
  wire _32425 = uncoded_block[974] ^ uncoded_block[976];
  wire _32426 = _467 ^ _32425;
  wire _32427 = uncoded_block[977] ^ uncoded_block[980];
  wire _32428 = _32427 ^ _476;
  wire _32429 = _32426 ^ _32428;
  wire _32430 = _32424 ^ _32429;
  wire _32431 = uncoded_block[997] ^ uncoded_block[1001];
  wire _32432 = _22575 ^ _32431;
  wire _32433 = _1319 ^ _32432;
  wire _32434 = _2112 ^ _487;
  wire _32435 = _2893 ^ _8299;
  wire _32436 = _32434 ^ _32435;
  wire _32437 = _32433 ^ _32436;
  wire _32438 = _32430 ^ _32437;
  wire _32439 = _2121 ^ _2898;
  wire _32440 = _32439 ^ _8880;
  wire _32441 = _502 ^ _6475;
  wire _32442 = _32441 ^ _11115;
  wire _32443 = _32440 ^ _32442;
  wire _32444 = _1359 ^ _8311;
  wire _32445 = _2916 ^ _2142;
  wire _32446 = _32444 ^ _32445;
  wire _32447 = _7724 ^ _2928;
  wire _32448 = _31183 ^ _32447;
  wire _32449 = _32446 ^ _32448;
  wire _32450 = _32443 ^ _32449;
  wire _32451 = _32438 ^ _32450;
  wire _32452 = _32420 ^ _32451;
  wire _32453 = _32387 ^ _32452;
  wire _32454 = _32322 ^ _32453;
  wire _32455 = _5839 ^ _536;
  wire _32456 = _5842 ^ _13316;
  wire _32457 = _32455 ^ _32456;
  wire _32458 = _1385 ^ _3713;
  wire _32459 = _21690 ^ _32458;
  wire _32460 = _32457 ^ _32459;
  wire _32461 = _11147 ^ _12789;
  wire _32462 = _5854 ^ _15894;
  wire _32463 = _32461 ^ _32462;
  wire _32464 = _8343 ^ _13866;
  wire _32465 = _32464 ^ _13870;
  wire _32466 = _32463 ^ _32465;
  wire _32467 = _32460 ^ _32466;
  wire _32468 = uncoded_block[1145] ^ uncoded_block[1150];
  wire _32469 = _2179 ^ _32468;
  wire _32470 = _32469 ^ _2187;
  wire _32471 = _10043 ^ _1407;
  wire _32472 = _5193 ^ _10046;
  wire _32473 = _32471 ^ _32472;
  wire _32474 = _32470 ^ _32473;
  wire _32475 = _7154 ^ _3739;
  wire _32476 = _17396 ^ _6519;
  wire _32477 = _32475 ^ _32476;
  wire _32478 = _2195 ^ _2200;
  wire _32479 = _21257 ^ _21259;
  wire _32480 = _32478 ^ _32479;
  wire _32481 = _32477 ^ _32480;
  wire _32482 = _32474 ^ _32481;
  wire _32483 = _32467 ^ _32482;
  wire _32484 = uncoded_block[1199] ^ uncoded_block[1204];
  wire _32485 = _32484 ^ _2210;
  wire _32486 = _32485 ^ _5210;
  wire _32487 = _1428 ^ _2219;
  wire _32488 = _2220 ^ _608;
  wire _32489 = _32487 ^ _32488;
  wire _32490 = _32486 ^ _32489;
  wire _32491 = _5891 ^ _8377;
  wire _32492 = _15926 ^ _3771;
  wire _32493 = _32491 ^ _32492;
  wire _32494 = _16915 ^ _8963;
  wire _32495 = _5229 ^ _24010;
  wire _32496 = _32494 ^ _32495;
  wire _32497 = _32493 ^ _32496;
  wire _32498 = _32490 ^ _32497;
  wire _32499 = _22195 ^ _30362;
  wire _32500 = uncoded_block[1270] ^ uncoded_block[1275];
  wire _32501 = _9532 ^ _32500;
  wire _32502 = _32501 ^ _11194;
  wire _32503 = _32499 ^ _32502;
  wire _32504 = _12838 ^ _10647;
  wire _32505 = _32504 ^ _11199;
  wire _32506 = uncoded_block[1307] ^ uncoded_block[1311];
  wire _32507 = _32506 ^ _4540;
  wire _32508 = _32507 ^ _20319;
  wire _32509 = _32505 ^ _32508;
  wire _32510 = _32503 ^ _32509;
  wire _32511 = _32498 ^ _32510;
  wire _32512 = _32483 ^ _32511;
  wire _32513 = uncoded_block[1329] ^ uncoded_block[1331];
  wire _32514 = _656 ^ _32513;
  wire _32515 = _21753 ^ _5259;
  wire _32516 = _32514 ^ _32515;
  wire _32517 = _1497 ^ _5268;
  wire _32518 = uncoded_block[1350] ^ uncoded_block[1354];
  wire _32519 = _32518 ^ _12857;
  wire _32520 = _32517 ^ _32519;
  wire _32521 = _32516 ^ _32520;
  wire _32522 = _6588 ^ _3052;
  wire _32523 = _9572 ^ _3055;
  wire _32524 = _32522 ^ _32523;
  wire _32525 = uncoded_block[1383] ^ uncoded_block[1389];
  wire _32526 = _3058 ^ _32525;
  wire _32527 = _2293 ^ _1516;
  wire _32528 = _32526 ^ _32527;
  wire _32529 = _32524 ^ _32528;
  wire _32530 = _32521 ^ _32529;
  wire _32531 = uncoded_block[1404] ^ uncoded_block[1409];
  wire _32532 = _32531 ^ _3069;
  wire _32533 = _30395 ^ _32532;
  wire _32534 = _13429 ^ _1533;
  wire _32535 = _7231 ^ _32534;
  wire _32536 = _32533 ^ _32535;
  wire _32537 = _3861 ^ _2319;
  wire _32538 = _20357 ^ _26309;
  wire _32539 = _32537 ^ _32538;
  wire _32540 = _724 ^ _24071;
  wire _32541 = _20853 ^ _32540;
  wire _32542 = _32539 ^ _32541;
  wire _32543 = _32536 ^ _32542;
  wire _32544 = _32530 ^ _32543;
  wire _32545 = _22707 ^ _2342;
  wire _32546 = _3884 ^ _7861;
  wire _32547 = _32545 ^ _32546;
  wire _32548 = _25426 ^ _9614;
  wire _32549 = uncoded_block[1505] ^ uncoded_block[1514];
  wire _32550 = _1572 ^ _32549;
  wire _32551 = _32548 ^ _32550;
  wire _32552 = _32547 ^ _32551;
  wire _32553 = _5337 ^ _2357;
  wire _32554 = _1581 ^ _6647;
  wire _32555 = _32553 ^ _32554;
  wire _32556 = _26789 ^ _6652;
  wire _32557 = _32555 ^ _32556;
  wire _32558 = _32552 ^ _32557;
  wire _32559 = _1590 ^ _5355;
  wire _32560 = _32559 ^ _13473;
  wire _32561 = _9070 ^ _1597;
  wire _32562 = _10161 ^ _15026;
  wire _32563 = _32561 ^ _32562;
  wire _32564 = _32560 ^ _32563;
  wire _32565 = uncoded_block[1575] ^ uncoded_block[1580];
  wire _32566 = _4647 ^ _32565;
  wire _32567 = uncoded_block[1581] ^ uncoded_block[1586];
  wire _32568 = _32567 ^ _11841;
  wire _32569 = _32566 ^ _32568;
  wire _32570 = _13996 ^ _11847;
  wire _32571 = _798 ^ _5380;
  wire _32572 = _32570 ^ _32571;
  wire _32573 = _32569 ^ _32572;
  wire _32574 = _32564 ^ _32573;
  wire _32575 = _32558 ^ _32574;
  wire _32576 = _32544 ^ _32575;
  wire _32577 = _32512 ^ _32576;
  wire _32578 = _18020 ^ _31746;
  wire _32579 = _27974 ^ _32578;
  wire _32580 = _3942 ^ _3166;
  wire _32581 = _7914 ^ _5392;
  wire _32582 = _32580 ^ _32581;
  wire _32583 = _32579 ^ _32582;
  wire _32584 = _3951 ^ _10757;
  wire _32585 = _32584 ^ _4679;
  wire _32586 = _822 ^ _10196;
  wire _32587 = _1654 ^ _7319;
  wire _32588 = _32586 ^ _32587;
  wire _32589 = _32585 ^ _32588;
  wire _32590 = _32583 ^ _32589;
  wire _32591 = _11319 ^ _5406;
  wire _32592 = _6701 ^ _32591;
  wire _32593 = _17040 ^ _3187;
  wire _32594 = _20429 ^ _3972;
  wire _32595 = _32593 ^ _32594;
  wire _32596 = _32592 ^ _32595;
  wire _32597 = _11327 ^ _845;
  wire _32598 = _3976 ^ _2437;
  wire _32599 = _32597 ^ _32598;
  wire _32600 = uncoded_block[1711] ^ uncoded_block[1716];
  wire _32601 = _32600 ^ _20923;
  wire _32602 = _32601 ^ uncoded_block[1722];
  wire _32603 = _32599 ^ _32602;
  wire _32604 = _32596 ^ _32603;
  wire _32605 = _32590 ^ _32604;
  wire _32606 = _32577 ^ _32605;
  wire _32607 = _32454 ^ _32606;
  wire _32608 = _1 ^ _4712;
  wire _32609 = uncoded_block[7] ^ uncoded_block[12];
  wire _32610 = _32609 ^ _6086;
  wire _32611 = _32608 ^ _32610;
  wire _32612 = _4716 ^ _9694;
  wire _32613 = uncoded_block[30] ^ uncoded_block[40];
  wire _32614 = _6093 ^ _32613;
  wire _32615 = _32612 ^ _32614;
  wire _32616 = _32611 ^ _32615;
  wire _32617 = _20457 ^ _12425;
  wire _32618 = _32617 ^ _8555;
  wire _32619 = _13547 ^ _888;
  wire _32620 = _13552 ^ _894;
  wire _32621 = _32619 ^ _32620;
  wire _32622 = _32618 ^ _32621;
  wire _32623 = _32616 ^ _32622;
  wire _32624 = _34 ^ _3241;
  wire _32625 = _32624 ^ _17076;
  wire _32626 = _41 ^ _18077;
  wire _32627 = _8566 ^ _4741;
  wire _32628 = _32626 ^ _32627;
  wire _32629 = _32625 ^ _32628;
  wire _32630 = _4031 ^ _7990;
  wire _32631 = _1729 ^ _3255;
  wire _32632 = _32630 ^ _32631;
  wire _32633 = _1730 ^ _1733;
  wire _32634 = uncoded_block[129] ^ uncoded_block[132];
  wire _32635 = _32634 ^ _15112;
  wire _32636 = _32633 ^ _32635;
  wire _32637 = _32632 ^ _32636;
  wire _32638 = _32629 ^ _32637;
  wire _32639 = _32623 ^ _32638;
  wire _32640 = _5461 ^ _7392;
  wire _32641 = _19529 ^ _32640;
  wire _32642 = _15622 ^ _9186;
  wire _32643 = _1748 ^ _19536;
  wire _32644 = _32642 ^ _32643;
  wire _32645 = _32641 ^ _32644;
  wire _32646 = _6788 ^ _15123;
  wire _32647 = _32646 ^ _25089;
  wire _32648 = _941 ^ _20004;
  wire _32649 = _2529 ^ _89;
  wire _32650 = _32648 ^ _32649;
  wire _32651 = _32647 ^ _32650;
  wire _32652 = _32645 ^ _32651;
  wire _32653 = _94 ^ _9745;
  wire _32654 = _29634 ^ _8600;
  wire _32655 = _32653 ^ _32654;
  wire _32656 = _2540 ^ _17613;
  wire _32657 = _17617 ^ _6814;
  wire _32658 = _32656 ^ _32657;
  wire _32659 = _32655 ^ _32658;
  wire _32660 = _25993 ^ _968;
  wire _32661 = _32660 ^ _11413;
  wire _32662 = _17127 ^ _6180;
  wire _32663 = _7432 ^ _4800;
  wire _32664 = _32662 ^ _32663;
  wire _32665 = _32661 ^ _32664;
  wire _32666 = _32659 ^ _32665;
  wire _32667 = _32652 ^ _32666;
  wire _32668 = _32639 ^ _32667;
  wire _32669 = _1788 ^ _6187;
  wire _32670 = _13607 ^ _32669;
  wire _32671 = _26443 ^ _30549;
  wire _32672 = _32670 ^ _32671;
  wire _32673 = _8632 ^ _10876;
  wire _32674 = _11968 ^ _32673;
  wire _32675 = _2573 ^ _2577;
  wire _32676 = uncoded_block[301] ^ uncoded_block[307];
  wire _32677 = _32676 ^ _5528;
  wire _32678 = _32675 ^ _32677;
  wire _32679 = _32674 ^ _32678;
  wire _32680 = _32672 ^ _32679;
  wire _32681 = _4117 ^ _1006;
  wire _32682 = uncoded_block[324] ^ uncoded_block[328];
  wire _32683 = _1008 ^ _32682;
  wire _32684 = _32681 ^ _32683;
  wire _32685 = uncoded_block[330] ^ uncoded_block[337];
  wire _32686 = _32685 ^ _9242;
  wire _32687 = uncoded_block[341] ^ uncoded_block[346];
  wire _32688 = _32687 ^ _15684;
  wire _32689 = _32686 ^ _32688;
  wire _32690 = _32684 ^ _32689;
  wire _32691 = _168 ^ _6873;
  wire _32692 = _10899 ^ _10901;
  wire _32693 = _32691 ^ _32692;
  wire _32694 = _28091 ^ _5554;
  wire _32695 = _32694 ^ _23782;
  wire _32696 = _32693 ^ _32695;
  wire _32697 = _32690 ^ _32696;
  wire _32698 = _32680 ^ _32697;
  wire _32699 = _4155 ^ _4867;
  wire _32700 = _2630 ^ _19613;
  wire _32701 = _32699 ^ _32700;
  wire _32702 = uncoded_block[422] ^ uncoded_block[427];
  wire _32703 = _32702 ^ _4878;
  wire _32704 = uncoded_block[441] ^ uncoded_block[448];
  wire _32705 = _5574 ^ _32704;
  wire _32706 = _32703 ^ _32705;
  wire _32707 = _32701 ^ _32706;
  wire _32708 = uncoded_block[449] ^ uncoded_block[453];
  wire _32709 = uncoded_block[454] ^ uncoded_block[459];
  wire _32710 = _32708 ^ _32709;
  wire _32711 = _15715 ^ _4890;
  wire _32712 = _32710 ^ _32711;
  wire _32713 = _1079 ^ _6906;
  wire _32714 = _5590 ^ _16693;
  wire _32715 = _32713 ^ _32714;
  wire _32716 = _32712 ^ _32715;
  wire _32717 = _32707 ^ _32716;
  wire _32718 = uncoded_block[491] ^ uncoded_block[498];
  wire _32719 = _8111 ^ _32718;
  wire _32720 = _20592 ^ _25167;
  wire _32721 = _32719 ^ _32720;
  wire _32722 = uncoded_block[514] ^ uncoded_block[517];
  wire _32723 = _9295 ^ _32722;
  wire _32724 = _32723 ^ _28124;
  wire _32725 = _32721 ^ _32724;
  wire _32726 = _26514 ^ _4926;
  wire _32727 = _14197 ^ _7540;
  wire _32728 = _32726 ^ _32727;
  wire _32729 = _1908 ^ _1118;
  wire _32730 = _32729 ^ _30180;
  wire _32731 = _32728 ^ _32730;
  wire _32732 = _32725 ^ _32731;
  wire _32733 = _32717 ^ _32732;
  wire _32734 = _32698 ^ _32733;
  wire _32735 = _32668 ^ _32734;
  wire _32736 = uncoded_block[563] ^ uncoded_block[566];
  wire _32737 = _1916 ^ _32736;
  wire _32738 = _6309 ^ _13168;
  wire _32739 = _32737 ^ _32738;
  wire _32740 = _17718 ^ _1933;
  wire _32741 = _32740 ^ _14734;
  wire _32742 = _32739 ^ _32741;
  wire _32743 = _1141 ^ _2700;
  wire _32744 = _32743 ^ _26978;
  wire _32745 = _3488 ^ _16234;
  wire _32746 = _32744 ^ _32745;
  wire _32747 = _32742 ^ _32746;
  wire _32748 = _8744 ^ _4960;
  wire _32749 = _32748 ^ _30196;
  wire _32750 = _1154 ^ _14228;
  wire _32751 = _290 ^ _1163;
  wire _32752 = _32750 ^ _32751;
  wire _32753 = _32749 ^ _32752;
  wire _32754 = _6336 ^ _296;
  wire _32755 = _6341 ^ _304;
  wire _32756 = _32754 ^ _32755;
  wire _32757 = _3513 ^ _2739;
  wire _32758 = _308 ^ _1177;
  wire _32759 = _32757 ^ _32758;
  wire _32760 = _32756 ^ _32759;
  wire _32761 = _32753 ^ _32760;
  wire _32762 = _32747 ^ _32761;
  wire _32763 = _1178 ^ _8760;
  wire _32764 = uncoded_block[681] ^ uncoded_block[686];
  wire _32765 = _8761 ^ _32764;
  wire _32766 = _32763 ^ _32765;
  wire _32767 = uncoded_block[691] ^ uncoded_block[694];
  wire _32768 = _2751 ^ _32767;
  wire _32769 = _32768 ^ _6991;
  wire _32770 = _32766 ^ _32769;
  wire _32771 = _333 ^ _6361;
  wire _32772 = uncoded_block[713] ^ uncoded_block[717];
  wire _32773 = _4996 ^ _32772;
  wire _32774 = _32771 ^ _32773;
  wire _32775 = _1984 ^ _343;
  wire _32776 = _32775 ^ _3545;
  wire _32777 = _32774 ^ _32776;
  wire _32778 = _32770 ^ _32777;
  wire _32779 = uncoded_block[732] ^ uncoded_block[736];
  wire _32780 = _8200 ^ _32779;
  wire _32781 = _350 ^ _352;
  wire _32782 = _32780 ^ _32781;
  wire _32783 = _11576 ^ _5013;
  wire _32784 = _4295 ^ _12663;
  wire _32785 = _32783 ^ _32784;
  wire _32786 = _32782 ^ _32785;
  wire _32787 = _3556 ^ _9914;
  wire _32788 = _2781 ^ _365;
  wire _32789 = _32787 ^ _32788;
  wire _32790 = _1218 ^ _15310;
  wire _32791 = _32790 ^ _13220;
  wire _32792 = _32789 ^ _32791;
  wire _32793 = _32786 ^ _32792;
  wire _32794 = _32778 ^ _32793;
  wire _32795 = _32762 ^ _32794;
  wire _32796 = uncoded_block[793] ^ uncoded_block[802];
  wire _32797 = _2798 ^ _32796;
  wire _32798 = _5716 ^ _32797;
  wire _32799 = uncoded_block[807] ^ uncoded_block[811];
  wire _32800 = _1235 ^ _32799;
  wire _32801 = _32800 ^ _19228;
  wire _32802 = _32798 ^ _32801;
  wire _32803 = _3587 ^ _2812;
  wire _32804 = _11033 ^ _32803;
  wire _32805 = _400 ^ _2035;
  wire _32806 = _32805 ^ _24816;
  wire _32807 = _32804 ^ _32806;
  wire _32808 = _32802 ^ _32807;
  wire _32809 = _21631 ^ _5742;
  wire _32810 = _2045 ^ _32809;
  wire _32811 = _414 ^ _1266;
  wire _32812 = _9950 ^ _32811;
  wire _32813 = _32810 ^ _32812;
  wire _32814 = _6416 ^ _8247;
  wire _32815 = _7653 ^ _32814;
  wire _32816 = uncoded_block[889] ^ uncoded_block[894];
  wire _32817 = _7660 ^ _32816;
  wire _32818 = _32817 ^ _2845;
  wire _32819 = _32815 ^ _32818;
  wire _32820 = _32813 ^ _32819;
  wire _32821 = _32808 ^ _32820;
  wire _32822 = _2065 ^ _2071;
  wire _32823 = _436 ^ _438;
  wire _32824 = _32822 ^ _32823;
  wire _32825 = _16827 ^ _18316;
  wire _32826 = _1294 ^ _32825;
  wire _32827 = _32824 ^ _32826;
  wire _32828 = _453 ^ _455;
  wire _32829 = _28588 ^ _32828;
  wire _32830 = _456 ^ _21191;
  wire _32831 = _32830 ^ _23928;
  wire _32832 = _32829 ^ _32831;
  wire _32833 = _32827 ^ _32832;
  wire _32834 = _10528 ^ _2872;
  wire _32835 = _7682 ^ _3656;
  wire _32836 = _32834 ^ _32835;
  wire _32837 = _15854 ^ _6451;
  wire _32838 = _23938 ^ _1323;
  wire _32839 = _32837 ^ _32838;
  wire _32840 = _32836 ^ _32839;
  wire _32841 = _9449 ^ _20730;
  wire _32842 = _27488 ^ _32841;
  wire _32843 = _11661 ^ _8296;
  wire _32844 = _2118 ^ _2121;
  wire _32845 = _32843 ^ _32844;
  wire _32846 = _32842 ^ _32845;
  wire _32847 = _32840 ^ _32846;
  wire _32848 = _32833 ^ _32847;
  wire _32849 = _32821 ^ _32848;
  wire _32850 = _32795 ^ _32849;
  wire _32851 = _32735 ^ _32850;
  wire _32852 = _13288 ^ _499;
  wire _32853 = _32852 ^ _1347;
  wire _32854 = uncoded_block[1042] ^ uncoded_block[1047];
  wire _32855 = _32854 ^ _1357;
  wire _32856 = _2136 ^ _13295;
  wire _32857 = _32855 ^ _32856;
  wire _32858 = _32853 ^ _32857;
  wire _32859 = _519 ^ _13849;
  wire _32860 = _32859 ^ _14358;
  wire _32861 = _21223 ^ _13307;
  wire _32862 = _32861 ^ _13856;
  wire _32863 = _32860 ^ _32862;
  wire _32864 = _32858 ^ _32863;
  wire _32865 = uncoded_block[1088] ^ uncoded_block[1093];
  wire _32866 = _1373 ^ _32865;
  wire _32867 = _3698 ^ _5843;
  wire _32868 = _32866 ^ _32867;
  wire _32869 = _543 ^ _4444;
  wire _32870 = _20761 ^ _7132;
  wire _32871 = _32869 ^ _32870;
  wire _32872 = _32868 ^ _32871;
  wire _32873 = uncoded_block[1116] ^ uncoded_block[1120];
  wire _32874 = _1386 ^ _32873;
  wire _32875 = _5176 ^ _8343;
  wire _32876 = _32874 ^ _32875;
  wire _32877 = _14380 ^ _8930;
  wire _32878 = uncoded_block[1143] ^ uncoded_block[1147];
  wire _32879 = _32878 ^ _15902;
  wire _32880 = _32877 ^ _32879;
  wire _32881 = _32876 ^ _32880;
  wire _32882 = _32872 ^ _32881;
  wire _32883 = _32864 ^ _32882;
  wire _32884 = uncoded_block[1162] ^ uncoded_block[1166];
  wire _32885 = _8937 ^ _32884;
  wire _32886 = _11160 ^ _9506;
  wire _32887 = _32885 ^ _32886;
  wire _32888 = uncoded_block[1176] ^ uncoded_block[1181];
  wire _32889 = _14901 ^ _32888;
  wire _32890 = _32889 ^ _12253;
  wire _32891 = _32887 ^ _32890;
  wire _32892 = _5203 ^ _4488;
  wire _32893 = _5882 ^ _8370;
  wire _32894 = _32892 ^ _32893;
  wire _32895 = _5885 ^ _7765;
  wire _32896 = _4496 ^ _2219;
  wire _32897 = _32895 ^ _32896;
  wire _32898 = _32894 ^ _32897;
  wire _32899 = _32891 ^ _32898;
  wire _32900 = _7168 ^ _5891;
  wire _32901 = _613 ^ _14921;
  wire _32902 = _32900 ^ _32901;
  wire _32903 = uncoded_block[1242] ^ uncoded_block[1246];
  wire _32904 = _19827 ^ _32903;
  wire _32905 = _1451 ^ _1455;
  wire _32906 = _32904 ^ _32905;
  wire _32907 = _32902 ^ _32906;
  wire _32908 = _5236 ^ _29058;
  wire _32909 = _26718 ^ _3793;
  wire _32910 = _3794 ^ _3797;
  wire _32911 = _32909 ^ _32910;
  wire _32912 = _32908 ^ _32911;
  wire _32913 = _32907 ^ _32912;
  wire _32914 = _32899 ^ _32913;
  wire _32915 = _32883 ^ _32914;
  wire _32916 = _3800 ^ _4531;
  wire _32917 = _17927 ^ _2254;
  wire _32918 = _32916 ^ _32917;
  wire _32919 = uncoded_block[1304] ^ uncoded_block[1308];
  wire _32920 = _32919 ^ _1480;
  wire _32921 = _1486 ^ _3029;
  wire _32922 = _32920 ^ _32921;
  wire _32923 = _32918 ^ _32922;
  wire _32924 = _7201 ^ _2268;
  wire _32925 = _5931 ^ _661;
  wire _32926 = _32924 ^ _32925;
  wire _32927 = _7814 ^ _11215;
  wire _32928 = uncoded_block[1350] ^ uncoded_block[1357];
  wire _32929 = _664 ^ _32928;
  wire _32930 = _32927 ^ _32929;
  wire _32931 = _32926 ^ _32930;
  wire _32932 = _32923 ^ _32931;
  wire _32933 = _5275 ^ _21762;
  wire _32934 = _32933 ^ _28337;
  wire _32935 = uncoded_block[1378] ^ uncoded_block[1383];
  wire _32936 = _32935 ^ _27590;
  wire _32937 = _9574 ^ _32936;
  wire _32938 = _32934 ^ _32937;
  wire _32939 = _6597 ^ _21774;
  wire _32940 = _16458 ^ _3846;
  wire _32941 = _32939 ^ _32940;
  wire _32942 = uncoded_block[1417] ^ uncoded_block[1422];
  wire _32943 = _20347 ^ _32942;
  wire _32944 = _25408 ^ _32943;
  wire _32945 = _32941 ^ _32944;
  wire _32946 = _32938 ^ _32945;
  wire _32947 = _32932 ^ _32946;
  wire _32948 = uncoded_block[1425] ^ uncoded_block[1429];
  wire _32949 = _32948 ^ _1531;
  wire _32950 = _4586 ^ _17470;
  wire _32951 = _32949 ^ _32950;
  wire _32952 = _3861 ^ _6613;
  wire _32953 = _3084 ^ _26763;
  wire _32954 = _32952 ^ _32953;
  wire _32955 = _32951 ^ _32954;
  wire _32956 = _720 ^ _7243;
  wire _32957 = _5314 ^ _18470;
  wire _32958 = _32956 ^ _32957;
  wire _32959 = _1555 ^ _3884;
  wire _32960 = _5990 ^ _12896;
  wire _32961 = _32959 ^ _32960;
  wire _32962 = _32958 ^ _32961;
  wire _32963 = _32955 ^ _32962;
  wire _32964 = uncoded_block[1497] ^ uncoded_block[1503];
  wire _32965 = _3890 ^ _32964;
  wire _32966 = _7874 ^ _750;
  wire _32967 = _32965 ^ _32966;
  wire _32968 = _7264 ^ _754;
  wire _32969 = _9059 ^ _5343;
  wire _32970 = _32968 ^ _32969;
  wire _32971 = _32967 ^ _32970;
  wire _32972 = _8474 ^ _9631;
  wire _32973 = _1586 ^ _12917;
  wire _32974 = _32972 ^ _32973;
  wire _32975 = uncoded_block[1541] ^ uncoded_block[1543];
  wire _32976 = _32975 ^ _4634;
  wire _32977 = _2367 ^ _13472;
  wire _32978 = _32976 ^ _32977;
  wire _32979 = _32974 ^ _32978;
  wire _32980 = _32971 ^ _32979;
  wire _32981 = _32963 ^ _32980;
  wire _32982 = _32947 ^ _32981;
  wire _32983 = _32915 ^ _32982;
  wire _32984 = _767 ^ _15528;
  wire _32985 = uncoded_block[1558] ^ uncoded_block[1563];
  wire _32986 = _32985 ^ _4644;
  wire _32987 = _32984 ^ _32986;
  wire _32988 = _5363 ^ _9080;
  wire _32989 = _782 ^ _12369;
  wire _32990 = _32988 ^ _32989;
  wire _32991 = _32987 ^ _32990;
  wire _32992 = _25008 ^ _20401;
  wire _32993 = _4654 ^ _29550;
  wire _32994 = _32992 ^ _32993;
  wire _32995 = _9088 ^ _5380;
  wire _32996 = _801 ^ _17020;
  wire _32997 = _32995 ^ _32996;
  wire _32998 = _32994 ^ _32997;
  wire _32999 = _32991 ^ _32998;
  wire _33000 = _804 ^ _18023;
  wire _33001 = _2400 ^ _4667;
  wire _33002 = _33000 ^ _33001;
  wire _33003 = uncoded_block[1633] ^ uncoded_block[1638];
  wire _33004 = _5388 ^ _33003;
  wire _33005 = _3948 ^ _3951;
  wire _33006 = _33004 ^ _33005;
  wire _33007 = _33002 ^ _33006;
  wire _33008 = _7312 ^ _819;
  wire _33009 = _18030 ^ _2414;
  wire _33010 = _33008 ^ _33009;
  wire _33011 = _16049 ^ _3180;
  wire _33012 = uncoded_block[1674] ^ uncoded_block[1680];
  wire _33013 = _22763 ^ _33012;
  wire _33014 = _33011 ^ _33013;
  wire _33015 = _33010 ^ _33014;
  wire _33016 = _33007 ^ _33015;
  wire _33017 = _32999 ^ _33016;
  wire _33018 = uncoded_block[1684] ^ uncoded_block[1688];
  wire _33019 = _33018 ^ _7331;
  wire _33020 = _840 ^ _1669;
  wire _33021 = _33019 ^ _33020;
  wire _33022 = _10778 ^ _852;
  wire _33023 = _16550 ^ _33022;
  wire _33024 = _33021 ^ _33023;
  wire _33025 = uncoded_block[1714] ^ uncoded_block[1719];
  wire _33026 = _33025 ^ uncoded_block[1720];
  wire _33027 = _33024 ^ _33026;
  wire _33028 = _33017 ^ _33027;
  wire _33029 = _32983 ^ _33028;
  wire _33030 = _32851 ^ _33029;
  wire _33031 = uncoded_block[11] ^ uncoded_block[16];
  wire _33032 = _4 ^ _33031;
  wire _33033 = _19493 ^ _33032;
  wire _33034 = _4716 ^ _3220;
  wire _33035 = _9694 ^ _9143;
  wire _33036 = _33034 ^ _33035;
  wire _33037 = _33033 ^ _33036;
  wire _33038 = _11 ^ _14047;
  wire _33039 = _12425 ^ _8554;
  wire _33040 = _33038 ^ _33039;
  wire _33041 = uncoded_block[51] ^ uncoded_block[56];
  wire _33042 = _9150 ^ _33041;
  wire _33043 = _33042 ^ _20946;
  wire _33044 = _33040 ^ _33043;
  wire _33045 = _33037 ^ _33044;
  wire _33046 = _34 ^ _5440;
  wire _33047 = _1712 ^ _4735;
  wire _33048 = _33046 ^ _33047;
  wire _33049 = uncoded_block[84] ^ uncoded_block[89];
  wire _33050 = _41 ^ _33049;
  wire _33051 = _903 ^ _30498;
  wire _33052 = _33050 ^ _33051;
  wire _33053 = _33048 ^ _33052;
  wire _33054 = _3249 ^ _6120;
  wire _33055 = _33054 ^ _6764;
  wire _33056 = uncoded_block[116] ^ uncoded_block[118];
  wire _33057 = _10816 ^ _33056;
  wire _33058 = uncoded_block[123] ^ uncoded_block[126];
  wire _33059 = _25070 ^ _33058;
  wire _33060 = _33057 ^ _33059;
  wire _33061 = _33055 ^ _33060;
  wire _33062 = _33053 ^ _33061;
  wire _33063 = _33045 ^ _33062;
  wire _33064 = _1733 ^ _8579;
  wire _33065 = _924 ^ _8581;
  wire _33066 = _33064 ^ _33065;
  wire _33067 = uncoded_block[143] ^ uncoded_block[148];
  wire _33068 = _7999 ^ _33067;
  wire _33069 = uncoded_block[160] ^ uncoded_block[163];
  wire _33070 = _20973 ^ _33069;
  wire _33071 = _33068 ^ _33070;
  wire _33072 = _33066 ^ _33071;
  wire _33073 = _29624 ^ _1752;
  wire _33074 = _938 ^ _20979;
  wire _33075 = _33073 ^ _33074;
  wire _33076 = _5479 ^ _944;
  wire _33077 = uncoded_block[191] ^ uncoded_block[194];
  wire _33078 = _4773 ^ _33077;
  wire _33079 = _33076 ^ _33078;
  wire _33080 = _33075 ^ _33079;
  wire _33081 = _33072 ^ _33080;
  wire _33082 = uncoded_block[205] ^ uncoded_block[209];
  wire _33083 = _33082 ^ _98;
  wire _33084 = _16117 ^ _33083;
  wire _33085 = _16618 ^ _6814;
  wire _33086 = _961 ^ _33085;
  wire _33087 = _33084 ^ _33086;
  wire _33088 = uncoded_block[233] ^ uncoded_block[236];
  wire _33089 = _4081 ^ _33088;
  wire _33090 = _33089 ^ _13049;
  wire _33091 = _113 ^ _5505;
  wire _33092 = _11954 ^ _1785;
  wire _33093 = _33091 ^ _33092;
  wire _33094 = _33090 ^ _33093;
  wire _33095 = _33087 ^ _33094;
  wire _33096 = _33081 ^ _33095;
  wire _33097 = _33063 ^ _33096;
  wire _33098 = _25998 ^ _30977;
  wire _33099 = uncoded_block[268] ^ uncoded_block[270];
  wire _33100 = _33099 ^ _20527;
  wire _33101 = _6837 ^ _2571;
  wire _33102 = _33100 ^ _33101;
  wire _33103 = _33098 ^ _33102;
  wire _33104 = _995 ^ _17142;
  wire _33105 = _17144 ^ _6845;
  wire _33106 = _33104 ^ _33105;
  wire _33107 = _6846 ^ _11439;
  wire _33108 = _6208 ^ _1009;
  wire _33109 = _33107 ^ _33108;
  wire _33110 = _33106 ^ _33109;
  wire _33111 = _33103 ^ _33110;
  wire _33112 = uncoded_block[329] ^ uncoded_block[334];
  wire _33113 = _33112 ^ _8646;
  wire _33114 = _11982 ^ _33113;
  wire _33115 = _159 ^ _1023;
  wire _33116 = _11451 ^ _33115;
  wire _33117 = _33114 ^ _33116;
  wire _33118 = _5541 ^ _24229;
  wire _33119 = uncoded_block[358] ^ uncoded_block[362];
  wire _33120 = _33119 ^ _4851;
  wire _33121 = _33118 ^ _33120;
  wire _33122 = _27738 ^ _25136;
  wire _33123 = _33121 ^ _33122;
  wire _33124 = _33117 ^ _33123;
  wire _33125 = _33111 ^ _33124;
  wire _33126 = _20056 ^ _9799;
  wire _33127 = _33126 ^ _19101;
  wire _33128 = uncoded_block[396] ^ uncoded_block[402];
  wire _33129 = _4152 ^ _33128;
  wire _33130 = _6244 ^ _1052;
  wire _33131 = _33129 ^ _33130;
  wire _33132 = _33127 ^ _33131;
  wire _33133 = _4868 ^ _12548;
  wire _33134 = _4163 ^ _8672;
  wire _33135 = _33133 ^ _33134;
  wire _33136 = uncoded_block[427] ^ uncoded_block[432];
  wire _33137 = _33136 ^ _6255;
  wire _33138 = _16187 ^ _205;
  wire _33139 = _33137 ^ _33138;
  wire _33140 = _33135 ^ _33139;
  wire _33141 = _33132 ^ _33140;
  wire _33142 = _206 ^ _7498;
  wire _33143 = _1866 ^ _17185;
  wire _33144 = _33142 ^ _33143;
  wire _33145 = _10926 ^ _8683;
  wire _33146 = _9283 ^ _6906;
  wire _33147 = _33145 ^ _33146;
  wire _33148 = _33144 ^ _33147;
  wire _33149 = _4895 ^ _15212;
  wire _33150 = _12026 ^ _33149;
  wire _33151 = _5600 ^ _2664;
  wire _33152 = _33151 ^ _1095;
  wire _33153 = _33150 ^ _33152;
  wire _33154 = _33148 ^ _33153;
  wire _33155 = _33141 ^ _33154;
  wire _33156 = _33125 ^ _33155;
  wire _33157 = _33097 ^ _33156;
  wire _33158 = _1887 ^ _5611;
  wire _33159 = _8705 ^ _4208;
  wire _33160 = _33158 ^ _33159;
  wire _33161 = _3444 ^ _1108;
  wire _33162 = uncoded_block[525] ^ uncoded_block[528];
  wire _33163 = _33162 ^ _15230;
  wire _33164 = _33161 ^ _33163;
  wire _33165 = _33160 ^ _33164;
  wire _33166 = _1115 ^ _2684;
  wire _33167 = _2687 ^ _5630;
  wire _33168 = _33166 ^ _33167;
  wire _33169 = uncoded_block[554] ^ uncoded_block[559];
  wire _33170 = _33169 ^ _19153;
  wire _33171 = _4223 ^ _1931;
  wire _33172 = _33170 ^ _33171;
  wire _33173 = _33168 ^ _33172;
  wire _33174 = _33165 ^ _33173;
  wire _33175 = _16225 ^ _28515;
  wire _33176 = _10408 ^ _1145;
  wire _33177 = uncoded_block[606] ^ uncoded_block[611];
  wire _33178 = _33177 ^ _281;
  wire _33179 = _33176 ^ _33178;
  wire _33180 = _33175 ^ _33179;
  wire _33181 = _3495 ^ _1154;
  wire _33182 = _1953 ^ _6330;
  wire _33183 = _33181 ^ _33182;
  wire _33184 = _6331 ^ _11543;
  wire _33185 = _33184 ^ _9878;
  wire _33186 = _33183 ^ _33185;
  wire _33187 = _33180 ^ _33186;
  wire _33188 = _33174 ^ _33187;
  wire _33189 = _1164 ^ _6973;
  wire _33190 = uncoded_block[652] ^ uncoded_block[655];
  wire _33191 = _33190 ^ _3513;
  wire _33192 = _33189 ^ _33191;
  wire _33193 = _2739 ^ _4264;
  wire _33194 = uncoded_block[675] ^ uncoded_block[678];
  wire _33195 = _15775 ^ _33194;
  wire _33196 = _33193 ^ _33195;
  wire _33197 = _33192 ^ _33196;
  wire _33198 = _15280 ^ _325;
  wire _33199 = _33198 ^ _19685;
  wire _33200 = _6992 ^ _6361;
  wire _33201 = _28542 ^ _33200;
  wire _33202 = _33199 ^ _33201;
  wire _33203 = _33197 ^ _33202;
  wire _33204 = uncoded_block[707] ^ uncoded_block[710];
  wire _33205 = uncoded_block[711] ^ uncoded_block[713];
  wire _33206 = _33204 ^ _33205;
  wire _33207 = _4999 ^ _8198;
  wire _33208 = _33206 ^ _33207;
  wire _33209 = _4283 ^ _29765;
  wire _33210 = _15788 ^ _2770;
  wire _33211 = _33209 ^ _33210;
  wire _33212 = _33208 ^ _33211;
  wire _33213 = uncoded_block[741] ^ uncoded_block[746];
  wire _33214 = _33213 ^ _4295;
  wire _33215 = _33214 ^ _26576;
  wire _33216 = _18740 ^ _365;
  wire _33217 = uncoded_block[770] ^ uncoded_block[774];
  wire _33218 = uncoded_block[782] ^ uncoded_block[786];
  wire _33219 = _33217 ^ _33218;
  wire _33220 = _33216 ^ _33219;
  wire _33221 = _33215 ^ _33220;
  wire _33222 = _33212 ^ _33221;
  wire _33223 = _33203 ^ _33222;
  wire _33224 = _33188 ^ _33223;
  wire _33225 = _19709 ^ _14282;
  wire _33226 = _7628 ^ _26589;
  wire _33227 = _33225 ^ _33226;
  wire _33228 = _389 ^ _14287;
  wire _33229 = uncoded_block[812] ^ uncoded_block[816];
  wire _33230 = _33229 ^ _2028;
  wire _33231 = _33228 ^ _33230;
  wire _33232 = _33227 ^ _33231;
  wire _33233 = _27843 ^ _1246;
  wire _33234 = _2032 ^ _3590;
  wire _33235 = _33233 ^ _33234;
  wire _33236 = _7042 ^ _32392;
  wire _33237 = _33235 ^ _33236;
  wire _33238 = _33232 ^ _33237;
  wire _33239 = uncoded_block[846] ^ uncoded_block[850];
  wire _33240 = _4339 ^ _33239;
  wire _33241 = _6406 ^ _7049;
  wire _33242 = _33240 ^ _33241;
  wire _33243 = uncoded_block[868] ^ uncoded_block[873];
  wire _33244 = _33243 ^ _417;
  wire _33245 = _13788 ^ _33244;
  wire _33246 = _33242 ^ _33245;
  wire _33247 = uncoded_block[876] ^ uncoded_block[879];
  wire _33248 = _33247 ^ _2836;
  wire _33249 = uncoded_block[884] ^ uncoded_block[890];
  wire _33250 = uncoded_block[891] ^ uncoded_block[899];
  wire _33251 = _33249 ^ _33250;
  wire _33252 = _33248 ^ _33251;
  wire _33253 = uncoded_block[900] ^ uncoded_block[906];
  wire _33254 = _33253 ^ _1284;
  wire _33255 = _19252 ^ _25731;
  wire _33256 = _33254 ^ _33255;
  wire _33257 = _33252 ^ _33256;
  wire _33258 = _33246 ^ _33257;
  wire _33259 = _33238 ^ _33258;
  wire _33260 = _1295 ^ _16321;
  wire _33261 = _22555 ^ _33260;
  wire _33262 = _2862 ^ _452;
  wire _33263 = _16832 ^ _19747;
  wire _33264 = _33262 ^ _33263;
  wire _33265 = _33261 ^ _33264;
  wire _33266 = _29387 ^ _4382;
  wire _33267 = _1307 ^ _4385;
  wire _33268 = _33266 ^ _33267;
  wire _33269 = _7088 ^ _468;
  wire _33270 = _10532 ^ _33269;
  wire _33271 = _33268 ^ _33270;
  wire _33272 = _33265 ^ _33271;
  wire _33273 = _11091 ^ _11094;
  wire _33274 = uncoded_block[986] ^ uncoded_block[993];
  wire _33275 = _7689 ^ _33274;
  wire _33276 = _33273 ^ _33275;
  wire _33277 = _28985 ^ _2107;
  wire _33278 = _4404 ^ _27077;
  wire _33279 = _33277 ^ _33278;
  wire _33280 = _33276 ^ _33279;
  wire _33281 = _4410 ^ _2117;
  wire _33282 = _33281 ^ _30303;
  wire _33283 = _9998 ^ _8875;
  wire _33284 = _4418 ^ _7707;
  wire _33285 = _33283 ^ _33284;
  wire _33286 = _33282 ^ _33285;
  wire _33287 = _33280 ^ _33286;
  wire _33288 = _33272 ^ _33287;
  wire _33289 = _33259 ^ _33288;
  wire _33290 = _33224 ^ _33289;
  wire _33291 = _33157 ^ _33290;
  wire _33292 = _5810 ^ _6478;
  wire _33293 = _33292 ^ _4428;
  wire _33294 = _4433 ^ _522;
  wire _33295 = _18805 ^ _33294;
  wire _33296 = _33293 ^ _33295;
  wire _33297 = _2142 ^ _3689;
  wire _33298 = _8892 ^ _7722;
  wire _33299 = _33297 ^ _33298;
  wire _33300 = _19301 ^ _2928;
  wire _33301 = _26223 ^ _33300;
  wire _33302 = _33299 ^ _33301;
  wire _33303 = _33296 ^ _33302;
  wire _33304 = _2149 ^ _13857;
  wire _33305 = uncoded_block[1093] ^ uncoded_block[1097];
  wire _33306 = _33305 ^ _18365;
  wire _33307 = _33304 ^ _33306;
  wire _33308 = _13318 ^ _550;
  wire _33309 = _22614 ^ _16376;
  wire _33310 = _33308 ^ _33309;
  wire _33311 = _33307 ^ _33310;
  wire _33312 = uncoded_block[1125] ^ uncoded_block[1127];
  wire _33313 = _33312 ^ _6499;
  wire _33314 = uncoded_block[1132] ^ uncoded_block[1136];
  wire _33315 = _560 ^ _33314;
  wire _33316 = _33313 ^ _33315;
  wire _33317 = _5182 ^ _3724;
  wire _33318 = _4466 ^ _4468;
  wire _33319 = _33317 ^ _33318;
  wire _33320 = _33316 ^ _33319;
  wire _33321 = _33311 ^ _33320;
  wire _33322 = _33303 ^ _33321;
  wire _33323 = _9500 ^ _10043;
  wire _33324 = _6511 ^ _21248;
  wire _33325 = _33323 ^ _33324;
  wire _33326 = _3739 ^ _17396;
  wire _33327 = _33326 ^ _25800;
  wire _33328 = _33325 ^ _33327;
  wire _33329 = uncoded_block[1183] ^ uncoded_block[1188];
  wire _33330 = uncoded_block[1189] ^ uncoded_block[1192];
  wire _33331 = _33329 ^ _33330;
  wire _33332 = _1421 ^ _7163;
  wire _33333 = _33331 ^ _33332;
  wire _33334 = _6530 ^ _5209;
  wire _33335 = _1427 ^ _4496;
  wire _33336 = _33334 ^ _33335;
  wire _33337 = _33333 ^ _33336;
  wire _33338 = _33328 ^ _33337;
  wire _33339 = _1433 ^ _2986;
  wire _33340 = _2221 ^ _33339;
  wire _33341 = _29050 ^ _16408;
  wire _33342 = _29898 ^ _33341;
  wire _33343 = _33340 ^ _33342;
  wire _33344 = _5900 ^ _6549;
  wire _33345 = _16919 ^ _7792;
  wire _33346 = _12837 ^ _24023;
  wire _33347 = _33345 ^ _33346;
  wire _33348 = _33344 ^ _33347;
  wire _33349 = _33343 ^ _33348;
  wire _33350 = _33338 ^ _33349;
  wire _33351 = _33322 ^ _33350;
  wire _33352 = _13381 ^ _32094;
  wire _33353 = _2256 ^ _24938;
  wire _33354 = _33352 ^ _33353;
  wire _33355 = _2261 ^ _12287;
  wire _33356 = _26729 ^ _1494;
  wire _33357 = _33355 ^ _33356;
  wire _33358 = uncoded_block[1337] ^ uncoded_block[1345];
  wire _33359 = _33358 ^ _20327;
  wire _33360 = _11767 ^ _33359;
  wire _33361 = _33357 ^ _33360;
  wire _33362 = _33354 ^ _33361;
  wire _33363 = uncoded_block[1352] ^ uncoded_block[1354];
  wire _33364 = _33363 ^ _23581;
  wire _33365 = _3045 ^ _677;
  wire _33366 = _33364 ^ _33365;
  wire _33367 = _679 ^ _10668;
  wire _33368 = _16449 ^ _15966;
  wire _33369 = _33367 ^ _33368;
  wire _33370 = _33366 ^ _33369;
  wire _33371 = _6600 ^ _26749;
  wire _33372 = _16950 ^ _33371;
  wire _33373 = _2300 ^ _20347;
  wire _33374 = uncoded_block[1415] ^ uncoded_block[1417];
  wire _33375 = uncoded_block[1418] ^ uncoded_block[1423];
  wire _33376 = _33374 ^ _33375;
  wire _33377 = _33373 ^ _33376;
  wire _33378 = _33372 ^ _33377;
  wire _33379 = _33370 ^ _33378;
  wire _33380 = _33362 ^ _33379;
  wire _33381 = _709 ^ _9590;
  wire _33382 = _9591 ^ _2313;
  wire _33383 = _33381 ^ _33382;
  wire _33384 = _17470 ^ _24065;
  wire _33385 = uncoded_block[1445] ^ uncoded_block[1450];
  wire _33386 = _2321 ^ _33385;
  wire _33387 = _33384 ^ _33386;
  wire _33388 = _33383 ^ _33387;
  wire _33389 = _20852 ^ _7241;
  wire _33390 = _33389 ^ _29961;
  wire _33391 = _16977 ^ _12337;
  wire _33392 = _1559 ^ _5321;
  wire _33393 = _33391 ^ _33392;
  wire _33394 = _33390 ^ _33393;
  wire _33395 = _33388 ^ _33394;
  wire _33396 = _1563 ^ _8462;
  wire _33397 = _33396 ^ _27952;
  wire _33398 = _1572 ^ _3894;
  wire _33399 = _5333 ^ _21343;
  wire _33400 = _33398 ^ _33399;
  wire _33401 = _33397 ^ _33400;
  wire _33402 = _6643 ^ _22723;
  wire _33403 = _1582 ^ _5347;
  wire _33404 = _33402 ^ _33403;
  wire _33405 = _20386 ^ _6008;
  wire _33406 = _7274 ^ _14496;
  wire _33407 = _33405 ^ _33406;
  wire _33408 = _33404 ^ _33407;
  wire _33409 = _33401 ^ _33408;
  wire _33410 = _33395 ^ _33409;
  wire _33411 = _33380 ^ _33410;
  wire _33412 = _33351 ^ _33411;
  wire _33413 = _10160 ^ _14498;
  wire _33414 = _5359 ^ _33413;
  wire _33415 = _9081 ^ _15536;
  wire _33416 = _33414 ^ _33415;
  wire _33417 = _15537 ^ _15031;
  wire _33418 = _12934 ^ _11294;
  wire _33419 = _33417 ^ _33418;
  wire _33420 = _797 ^ _3936;
  wire _33421 = _10742 ^ _3154;
  wire _33422 = _33420 ^ _33421;
  wire _33423 = _33419 ^ _33422;
  wire _33424 = _33416 ^ _33423;
  wire _33425 = uncoded_block[1611] ^ uncoded_block[1618];
  wire _33426 = _33425 ^ _7911;
  wire _33427 = _7300 ^ _6685;
  wire _33428 = _33426 ^ _33427;
  wire _33429 = _5388 ^ _18965;
  wire _33430 = _33429 ^ _2409;
  wire _33431 = _33428 ^ _33430;
  wire _33432 = uncoded_block[1645] ^ uncoded_block[1651];
  wire _33433 = _3169 ^ _33432;
  wire _33434 = _10760 ^ _4680;
  wire _33435 = _33433 ^ _33434;
  wire _33436 = _17032 ^ _25476;
  wire _33437 = _33436 ^ _16540;
  wire _33438 = _33435 ^ _33437;
  wire _33439 = _33431 ^ _33438;
  wire _33440 = _33424 ^ _33439;
  wire _33441 = _14019 ^ _21393;
  wire _33442 = _844 ^ _8535;
  wire _33443 = _15063 ^ _27671;
  wire _33444 = _33442 ^ _33443;
  wire _33445 = _33441 ^ _33444;
  wire _33446 = uncoded_block[1711] ^ uncoded_block[1714];
  wire _33447 = _33446 ^ _1677;
  wire _33448 = _33447 ^ _10217;
  wire _33449 = _33445 ^ _33448;
  wire _33450 = _33440 ^ _33449;
  wire _33451 = _33412 ^ _33450;
  wire _33452 = _33291 ^ _33451;
  wire _33453 = _3993 ^ _6083;
  wire _33454 = _25495 ^ _33453;
  wire _33455 = _16564 ^ _4716;
  wire _33456 = _3219 ^ _11890;
  wire _33457 = _33455 ^ _33456;
  wire _33458 = _33454 ^ _33457;
  wire _33459 = _13543 ^ _21871;
  wire _33460 = _4723 ^ _3232;
  wire _33461 = _33459 ^ _33460;
  wire _33462 = _23255 ^ _2471;
  wire _33463 = _33462 ^ _7366;
  wire _33464 = _33461 ^ _33463;
  wire _33465 = _33458 ^ _33464;
  wire _33466 = _9705 ^ _25950;
  wire _33467 = uncoded_block[72] ^ uncoded_block[78];
  wire _33468 = _7976 ^ _33467;
  wire _33469 = _33466 ^ _33468;
  wire _33470 = _9161 ^ _14065;
  wire _33471 = _19515 ^ _14068;
  wire _33472 = _33470 ^ _33471;
  wire _33473 = _33469 ^ _33472;
  wire _33474 = _4028 ^ _7986;
  wire _33475 = _4032 ^ _3253;
  wire _33476 = _33474 ^ _33475;
  wire _33477 = _2502 ^ _13017;
  wire _33478 = _2499 ^ _33477;
  wire _33479 = _33476 ^ _33478;
  wire _33480 = _33473 ^ _33479;
  wire _33481 = _33465 ^ _33480;
  wire _33482 = _4042 ^ _15112;
  wire _33483 = _1736 ^ _5461;
  wire _33484 = _33482 ^ _33483;
  wire _33485 = uncoded_block[145] ^ uncoded_block[150];
  wire _33486 = _6138 ^ _33485;
  wire _33487 = uncoded_block[160] ^ uncoded_block[164];
  wire _33488 = _4049 ^ _33487;
  wire _33489 = _33486 ^ _33488;
  wire _33490 = _33484 ^ _33489;
  wire _33491 = _1751 ^ _6788;
  wire _33492 = _81 ^ _2524;
  wire _33493 = _33491 ^ _33492;
  wire _33494 = uncoded_block[180] ^ uncoded_block[188];
  wire _33495 = _33494 ^ _4773;
  wire _33496 = _6798 ^ _1763;
  wire _33497 = _33495 ^ _33496;
  wire _33498 = _33493 ^ _33497;
  wire _33499 = _33490 ^ _33498;
  wire _33500 = _94 ^ _3289;
  wire _33501 = _28043 ^ _1767;
  wire _33502 = _33500 ^ _33501;
  wire _33503 = _11409 ^ _4076;
  wire _33504 = uncoded_block[225] ^ uncoded_block[229];
  wire _33505 = _33504 ^ _2550;
  wire _33506 = _33503 ^ _33505;
  wire _33507 = _33502 ^ _33506;
  wire _33508 = _5504 ^ _8618;
  wire _33509 = _8034 ^ _9761;
  wire _33510 = uncoded_block[256] ^ uncoded_block[258];
  wire _33511 = _33510 ^ _7438;
  wire _33512 = _33509 ^ _33511;
  wire _33513 = _33508 ^ _33512;
  wire _33514 = _33507 ^ _33513;
  wire _33515 = _33499 ^ _33514;
  wire _33516 = _33481 ^ _33515;
  wire _33517 = uncoded_block[264] ^ uncoded_block[268];
  wire _33518 = _4096 ^ _33517;
  wire _33519 = _2566 ^ _10872;
  wire _33520 = _33518 ^ _33519;
  wire _33521 = _5512 ^ _19071;
  wire _33522 = uncoded_block[282] ^ uncoded_block[285];
  wire _33523 = _33522 ^ _10876;
  wire _33524 = _33521 ^ _33523;
  wire _33525 = _33520 ^ _33524;
  wire _33526 = _15665 ^ _1806;
  wire _33527 = _26012 ^ _4111;
  wire _33528 = _33526 ^ _33527;
  wire _33529 = _12515 ^ _15668;
  wire _33530 = _8056 ^ _11439;
  wire _33531 = _33529 ^ _33530;
  wire _33532 = _33528 ^ _33531;
  wire _33533 = _33525 ^ _33532;
  wire _33534 = uncoded_block[321] ^ uncoded_block[327];
  wire _33535 = _1814 ^ _33534;
  wire _33536 = _2584 ^ _4126;
  wire _33537 = _33535 ^ _33536;
  wire _33538 = _11984 ^ _2595;
  wire _33539 = _4131 ^ _3359;
  wire _33540 = _33538 ^ _33539;
  wire _33541 = _33537 ^ _33540;
  wire _33542 = _1024 ^ _1028;
  wire _33543 = _20554 ^ _21030;
  wire _33544 = _33542 ^ _33543;
  wire _33545 = _8075 ^ _1035;
  wire _33546 = _173 ^ _4143;
  wire _33547 = _33545 ^ _33546;
  wire _33548 = _33544 ^ _33547;
  wire _33549 = _33541 ^ _33548;
  wire _33550 = _33533 ^ _33549;
  wire _33551 = _3377 ^ _13102;
  wire _33552 = _33551 ^ _15695;
  wire _33553 = _2622 ^ _181;
  wire _33554 = _2625 ^ _1051;
  wire _33555 = _33553 ^ _33554;
  wire _33556 = _33552 ^ _33555;
  wire _33557 = uncoded_block[413] ^ uncoded_block[419];
  wire _33558 = _8091 ^ _33557;
  wire _33559 = _28098 ^ _2638;
  wire _33560 = _33558 ^ _33559;
  wire _33561 = _9271 ^ _3405;
  wire _33562 = _33561 ^ _24253;
  wire _33563 = _33560 ^ _33562;
  wire _33564 = _33556 ^ _33563;
  wire _33565 = uncoded_block[449] ^ uncoded_block[454];
  wire _33566 = _33565 ^ _212;
  wire _33567 = _8681 ^ _13662;
  wire _33568 = _33566 ^ _33567;
  wire _33569 = _1874 ^ _1878;
  wire _33570 = uncoded_block[477] ^ uncoded_block[480];
  wire _33571 = _24721 ^ _33570;
  wire _33572 = _33569 ^ _33571;
  wire _33573 = _33568 ^ _33572;
  wire _33574 = _4895 ^ _224;
  wire _33575 = _2664 ^ _7520;
  wire _33576 = _33574 ^ _33575;
  wire _33577 = uncoded_block[503] ^ uncoded_block[507];
  wire _33578 = _19135 ^ _33577;
  wire _33579 = _10376 ^ _3439;
  wire _33580 = _33578 ^ _33579;
  wire _33581 = _33576 ^ _33580;
  wire _33582 = _33573 ^ _33581;
  wire _33583 = _33564 ^ _33582;
  wire _33584 = _33550 ^ _33583;
  wire _33585 = _33516 ^ _33584;
  wire _33586 = _14193 ^ _1900;
  wire _33587 = uncoded_block[528] ^ uncoded_block[533];
  wire _33588 = _33587 ^ _243;
  wire _33589 = _33586 ^ _33588;
  wire _33590 = _14198 ^ _16715;
  wire _33591 = _6300 ^ _31904;
  wire _33592 = _33590 ^ _33591;
  wire _33593 = _33589 ^ _33592;
  wire _33594 = _8721 ^ _1916;
  wire _33595 = _33594 ^ _13695;
  wire _33596 = _6309 ^ _6942;
  wire _33597 = _262 ^ _1931;
  wire _33598 = _33596 ^ _33597;
  wire _33599 = _33595 ^ _33598;
  wire _33600 = _33593 ^ _33599;
  wire _33601 = _10404 ^ _270;
  wire _33602 = _18222 ^ _2700;
  wire _33603 = _33601 ^ _33602;
  wire _33604 = _4952 ^ _2707;
  wire _33605 = _2709 ^ _9870;
  wire _33606 = _33604 ^ _33605;
  wire _33607 = _33603 ^ _33606;
  wire _33608 = _23400 ^ _13713;
  wire _33609 = _4960 ^ _4963;
  wire _33610 = _33608 ^ _33609;
  wire _33611 = _287 ^ _1953;
  wire _33612 = _3501 ^ _31929;
  wire _33613 = _33611 ^ _33612;
  wire _33614 = _33610 ^ _33613;
  wire _33615 = _33607 ^ _33614;
  wire _33616 = _33600 ^ _33615;
  wire _33617 = _6342 ^ _15270;
  wire _33618 = _303 ^ _33617;
  wire _33619 = _15273 ^ _311;
  wire _33620 = _33619 ^ _27810;
  wire _33621 = _33618 ^ _33620;
  wire _33622 = _13731 ^ _1181;
  wire _33623 = _12636 ^ _2751;
  wire _33624 = _33622 ^ _33623;
  wire _33625 = _13735 ^ _4987;
  wire _33626 = uncoded_block[701] ^ uncoded_block[706];
  wire _33627 = _11562 ^ _33626;
  wire _33628 = _33625 ^ _33627;
  wire _33629 = _33624 ^ _33628;
  wire _33630 = _33621 ^ _33629;
  wire _33631 = _2762 ^ _19201;
  wire _33632 = _6367 ^ _7002;
  wire _33633 = _33631 ^ _33632;
  wire _33634 = _1203 ^ _4289;
  wire _33635 = _15301 ^ _2002;
  wire _33636 = _33634 ^ _33635;
  wire _33637 = _33633 ^ _33636;
  wire _33638 = uncoded_block[761] ^ uncoded_block[765];
  wire _33639 = _11012 ^ _33638;
  wire _33640 = _5709 ^ _11019;
  wire _33641 = _33639 ^ _33640;
  wire _33642 = _1221 ^ _9382;
  wire _33643 = uncoded_block[780] ^ uncoded_block[785];
  wire _33644 = _33643 ^ _1224;
  wire _33645 = _33642 ^ _33644;
  wire _33646 = _33641 ^ _33645;
  wire _33647 = _33637 ^ _33646;
  wire _33648 = _33630 ^ _33647;
  wire _33649 = _33616 ^ _33648;
  wire _33650 = _5033 ^ _2799;
  wire _33651 = _33650 ^ _26153;
  wire _33652 = _18286 ^ _2026;
  wire _33653 = _27838 ^ _33652;
  wire _33654 = _33651 ^ _33653;
  wire _33655 = _4324 ^ _1241;
  wire _33656 = uncoded_block[824] ^ uncoded_block[829];
  wire _33657 = _2029 ^ _33656;
  wire _33658 = _33655 ^ _33657;
  wire _33659 = uncoded_block[834] ^ uncoded_block[839];
  wire _33660 = _3590 ^ _33659;
  wire _33661 = _33660 ^ _5059;
  wire _33662 = _33658 ^ _33661;
  wire _33663 = _33654 ^ _33662;
  wire _33664 = _7643 ^ _12146;
  wire _33665 = _5061 ^ _33664;
  wire _33666 = _14300 ^ _5747;
  wire _33667 = _2824 ^ _7650;
  wire _33668 = _33666 ^ _33667;
  wire _33669 = _33665 ^ _33668;
  wire _33670 = _7054 ^ _416;
  wire _33671 = uncoded_block[873] ^ uncoded_block[875];
  wire _33672 = _33671 ^ _5078;
  wire _33673 = _33670 ^ _33672;
  wire _33674 = _3610 ^ _7660;
  wire _33675 = _4354 ^ _5085;
  wire _33676 = _33674 ^ _33675;
  wire _33677 = _33673 ^ _33676;
  wire _33678 = _33669 ^ _33677;
  wire _33679 = _33663 ^ _33678;
  wire _33680 = _5759 ^ _1280;
  wire _33681 = uncoded_block[905] ^ uncoded_block[911];
  wire _33682 = _33681 ^ _1287;
  wire _33683 = _33680 ^ _33682;
  wire _33684 = uncoded_block[922] ^ uncoded_block[927];
  wire _33685 = _33684 ^ _4371;
  wire _33686 = _21645 ^ _33685;
  wire _33687 = _33683 ^ _33686;
  wire _33688 = _448 ^ _2078;
  wire _33689 = _5101 ^ _9971;
  wire _33690 = _33688 ^ _33689;
  wire _33691 = _21187 ^ _21191;
  wire _33692 = _33691 ^ _27061;
  wire _33693 = _33690 ^ _33692;
  wire _33694 = _33687 ^ _33693;
  wire _33695 = _1308 ^ _1310;
  wire _33696 = _5108 ^ _1314;
  wire _33697 = _33695 ^ _33696;
  wire _33698 = _470 ^ _4391;
  wire _33699 = _11094 ^ _13825;
  wire _33700 = _33698 ^ _33699;
  wire _33701 = _33697 ^ _33700;
  wire _33702 = _11099 ^ _7691;
  wire _33703 = _22122 ^ _486;
  wire _33704 = _33702 ^ _33703;
  wire _33705 = _492 ^ _2120;
  wire _33706 = _5132 ^ _33705;
  wire _33707 = _33704 ^ _33706;
  wire _33708 = _33701 ^ _33707;
  wire _33709 = _33694 ^ _33708;
  wire _33710 = _33679 ^ _33709;
  wire _33711 = _33649 ^ _33710;
  wire _33712 = _33585 ^ _33711;
  wire _33713 = _5137 ^ _498;
  wire _33714 = _12756 ^ _1342;
  wire _33715 = _33713 ^ _33714;
  wire _33716 = _2129 ^ _6478;
  wire _33717 = _33716 ^ _13293;
  wire _33718 = _33715 ^ _33717;
  wire _33719 = _13844 ^ _8311;
  wire _33720 = _33719 ^ _19781;
  wire _33721 = uncoded_block[1067] ^ uncoded_block[1075];
  wire _33722 = _33721 ^ _2147;
  wire _33723 = _19301 ^ _4440;
  wire _33724 = _33722 ^ _33723;
  wire _33725 = _33720 ^ _33724;
  wire _33726 = _33718 ^ _33725;
  wire _33727 = _537 ^ _542;
  wire _33728 = _12224 ^ _8914;
  wire _33729 = _33727 ^ _33728;
  wire _33730 = _25323 ^ _10587;
  wire _33731 = _551 ^ _33730;
  wire _33732 = _33729 ^ _33731;
  wire _33733 = _2172 ^ _6499;
  wire _33734 = _564 ^ _1396;
  wire _33735 = _33733 ^ _33734;
  wire _33736 = uncoded_block[1153] ^ uncoded_block[1157];
  wire _33737 = _33736 ^ _578;
  wire _33738 = _17385 ^ _33737;
  wire _33739 = _33735 ^ _33738;
  wire _33740 = _33732 ^ _33739;
  wire _33741 = _33726 ^ _33740;
  wire _33742 = _1408 ^ _589;
  wire _33743 = _10601 ^ _33742;
  wire _33744 = _592 ^ _27116;
  wire _33745 = _12808 ^ _6522;
  wire _33746 = _33744 ^ _33745;
  wire _33747 = _33743 ^ _33746;
  wire _33748 = _8370 ^ _2209;
  wire _33749 = _28294 ^ _33748;
  wire _33750 = uncoded_block[1209] ^ uncoded_block[1213];
  wire _33751 = _33750 ^ _5889;
  wire _33752 = _33751 ^ _28302;
  wire _33753 = _33749 ^ _33752;
  wire _33754 = _33747 ^ _33753;
  wire _33755 = _13355 ^ _2986;
  wire _33756 = _7169 ^ _11732;
  wire _33757 = _33755 ^ _33756;
  wire _33758 = uncoded_block[1244] ^ uncoded_block[1247];
  wire _33759 = _2994 ^ _33758;
  wire _33760 = _33759 ^ _7779;
  wire _33761 = _33757 ^ _33760;
  wire _33762 = _2236 ^ _30361;
  wire _33763 = _627 ^ _3008;
  wire _33764 = _33762 ^ _33763;
  wire _33765 = _631 ^ _29472;
  wire _33766 = _25370 ^ _33765;
  wire _33767 = _33764 ^ _33766;
  wire _33768 = _33761 ^ _33767;
  wire _33769 = _33754 ^ _33768;
  wire _33770 = _33741 ^ _33769;
  wire _33771 = uncoded_block[1289] ^ uncoded_block[1293];
  wire _33772 = _24482 ^ _33771;
  wire _33773 = _22662 ^ _3805;
  wire _33774 = _33772 ^ _33773;
  wire _33775 = uncoded_block[1314] ^ uncoded_block[1320];
  wire _33776 = _33775 ^ _3029;
  wire _33777 = _14941 ^ _33776;
  wire _33778 = _33774 ^ _33777;
  wire _33779 = _4543 ^ _1490;
  wire _33780 = uncoded_block[1335] ^ uncoded_block[1339];
  wire _33781 = _5256 ^ _33780;
  wire _33782 = _33779 ^ _33781;
  wire _33783 = _1497 ^ _29486;
  wire _33784 = _14442 ^ _18436;
  wire _33785 = _33783 ^ _33784;
  wire _33786 = _33782 ^ _33785;
  wire _33787 = _33778 ^ _33786;
  wire _33788 = uncoded_block[1361] ^ uncoded_block[1365];
  wire _33789 = _28679 ^ _33788;
  wire _33790 = _33789 ^ _12865;
  wire _33791 = _22229 ^ _687;
  wire _33792 = _688 ^ _24511;
  wire _33793 = _33791 ^ _33792;
  wire _33794 = _33790 ^ _33793;
  wire _33795 = _23157 ^ _4571;
  wire _33796 = _33795 ^ _28689;
  wire _33797 = _5957 ^ _702;
  wire _33798 = _33797 ^ _29094;
  wire _33799 = _33796 ^ _33798;
  wire _33800 = _33794 ^ _33799;
  wire _33801 = _33787 ^ _33800;
  wire _33802 = _708 ^ _9025;
  wire _33803 = _1534 ^ _17470;
  wire _33804 = _33802 ^ _33803;
  wire _33805 = _24065 ^ _26763;
  wire _33806 = _16474 ^ _23174;
  wire _33807 = _33805 ^ _33806;
  wire _33808 = _33804 ^ _33807;
  wire _33809 = _23176 ^ _7247;
  wire _33810 = uncoded_block[1472] ^ uncoded_block[1477];
  wire _33811 = _33810 ^ _31294;
  wire _33812 = _33809 ^ _33811;
  wire _33813 = _739 ^ _1563;
  wire _33814 = _4610 ^ _6634;
  wire _33815 = _33813 ^ _33814;
  wire _33816 = _33812 ^ _33815;
  wire _33817 = _33808 ^ _33816;
  wire _33818 = uncoded_block[1520] ^ uncoded_block[1524];
  wire _33819 = _16004 ^ _33818;
  wire _33820 = _8466 ^ _33819;
  wire _33821 = _8474 ^ _24994;
  wire _33822 = _5347 ^ _20386;
  wire _33823 = _33821 ^ _33822;
  wire _33824 = _33820 ^ _33823;
  wire _33825 = _20387 ^ _5355;
  wire _33826 = _13471 ^ _17506;
  wire _33827 = _33825 ^ _33826;
  wire _33828 = _15022 ^ _1605;
  wire _33829 = _7285 ^ _9080;
  wire _33830 = _33828 ^ _33829;
  wire _33831 = _33827 ^ _33830;
  wire _33832 = _33824 ^ _33831;
  wire _33833 = _33817 ^ _33832;
  wire _33834 = _33801 ^ _33833;
  wire _33835 = _33770 ^ _33834;
  wire _33836 = _781 ^ _15535;
  wire _33837 = _33836 ^ _22739;
  wire _33838 = _788 ^ _1616;
  wire _33839 = uncoded_block[1596] ^ uncoded_block[1600];
  wire _33840 = _11292 ^ _33839;
  wire _33841 = _33838 ^ _33840;
  wire _33842 = _33837 ^ _33841;
  wire _33843 = _3937 ^ _6042;
  wire _33844 = _8503 ^ _33843;
  wire _33845 = uncoded_block[1617] ^ uncoded_block[1621];
  wire _33846 = _10181 ^ _33845;
  wire _33847 = uncoded_block[1622] ^ uncoded_block[1628];
  wire _33848 = _33847 ^ _15551;
  wire _33849 = _33846 ^ _33848;
  wire _33850 = _33844 ^ _33849;
  wire _33851 = _33842 ^ _33850;
  wire _33852 = uncoded_block[1636] ^ uncoded_block[1638];
  wire _33853 = _1641 ^ _33852;
  wire _33854 = _12383 ^ _13500;
  wire _33855 = _33853 ^ _33854;
  wire _33856 = _5394 ^ _4674;
  wire _33857 = _33856 ^ _4679;
  wire _33858 = _33855 ^ _33857;
  wire _33859 = _10760 ^ _6055;
  wire _33860 = _2419 ^ _7319;
  wire _33861 = _33859 ^ _33860;
  wire _33862 = uncoded_block[1675] ^ uncoded_block[1678];
  wire _33863 = _33862 ^ _17040;
  wire _33864 = _17036 ^ _33863;
  wire _33865 = _33861 ^ _33864;
  wire _33866 = _33858 ^ _33865;
  wire _33867 = _33851 ^ _33866;
  wire _33868 = _3187 ^ _3967;
  wire _33869 = _33868 ^ _21393;
  wire _33870 = _1669 ^ _8533;
  wire _33871 = _33870 ^ _12406;
  wire _33872 = _33869 ^ _33871;
  wire _33873 = _33872 ^ uncoded_block[1715];
  wire _33874 = _33867 ^ _33873;
  wire _33875 = _33835 ^ _33874;
  wire _33876 = _33712 ^ _33875;
  wire _33877 = _18539 ^ _1684;
  wire _33878 = _33877 ^ _15584;
  wire _33879 = _11343 ^ _6728;
  wire _33880 = _16074 ^ _33879;
  wire _33881 = _33878 ^ _33880;
  wire _33882 = _875 ^ _14569;
  wire _33883 = _2466 ^ _15594;
  wire _33884 = _33882 ^ _33883;
  wire _33885 = _1700 ^ _888;
  wire _33886 = uncoded_block[67] ^ uncoded_block[70];
  wire _33887 = _9705 ^ _33886;
  wire _33888 = _33885 ^ _33887;
  wire _33889 = _33884 ^ _33888;
  wire _33890 = _33881 ^ _33889;
  wire _33891 = uncoded_block[77] ^ uncoded_block[82];
  wire _33892 = _33891 ^ _11364;
  wire _33893 = _30494 ^ _33892;
  wire _33894 = uncoded_block[85] ^ uncoded_block[88];
  wire _33895 = _33894 ^ _8566;
  wire _33896 = _8567 ^ _14068;
  wire _33897 = _33895 ^ _33896;
  wire _33898 = _33893 ^ _33897;
  wire _33899 = uncoded_block[101] ^ uncoded_block[105];
  wire _33900 = _9718 ^ _33899;
  wire _33901 = _6126 ^ _13014;
  wire _33902 = _33900 ^ _33901;
  wire _33903 = _2501 ^ _7386;
  wire _33904 = _1733 ^ _20963;
  wire _33905 = _33903 ^ _33904;
  wire _33906 = _33902 ^ _33905;
  wire _33907 = _33898 ^ _33906;
  wire _33908 = _33890 ^ _33907;
  wire _33909 = uncoded_block[143] ^ uncoded_block[147];
  wire _33910 = _20969 ^ _33909;
  wire _33911 = _70 ^ _3269;
  wire _33912 = _33910 ^ _33911;
  wire _33913 = _4048 ^ _73;
  wire _33914 = _33913 ^ _23726;
  wire _33915 = _33912 ^ _33914;
  wire _33916 = _1749 ^ _1751;
  wire _33917 = uncoded_block[168] ^ uncoded_block[174];
  wire _33918 = _33917 ^ _13032;
  wire _33919 = _33916 ^ _33918;
  wire _33920 = _941 ^ _7409;
  wire _33921 = uncoded_block[191] ^ uncoded_block[196];
  wire _33922 = _33921 ^ _4068;
  wire _33923 = _33920 ^ _33922;
  wire _33924 = _33919 ^ _33923;
  wire _33925 = _33915 ^ _33924;
  wire _33926 = _15639 ^ _26879;
  wire _33927 = _6168 ^ _4791;
  wire _33928 = _19055 ^ _33927;
  wire _33929 = _33926 ^ _33928;
  wire _33930 = _2549 ^ _6822;
  wire _33931 = _6824 ^ _4085;
  wire _33932 = _33930 ^ _33931;
  wire _33933 = _14116 ^ _4803;
  wire _33934 = _9761 ^ _1786;
  wire _33935 = _33933 ^ _33934;
  wire _33936 = _33932 ^ _33935;
  wire _33937 = _33929 ^ _33936;
  wire _33938 = _33925 ^ _33937;
  wire _33939 = _33908 ^ _33938;
  wire _33940 = _12501 ^ _4099;
  wire _33941 = _3320 ^ _5512;
  wire _33942 = _33940 ^ _33941;
  wire _33943 = _1803 ^ _5522;
  wire _33944 = _1797 ^ _33943;
  wire _33945 = _33942 ^ _33944;
  wire _33946 = _28817 ^ _13615;
  wire _33947 = _8636 ^ _17144;
  wire _33948 = _33946 ^ _33947;
  wire _33949 = _1000 ^ _20536;
  wire _33950 = _33949 ^ _26456;
  wire _33951 = _33948 ^ _33950;
  wire _33952 = _33945 ^ _33951;
  wire _33953 = _1814 ^ _11441;
  wire _33954 = uncoded_block[327] ^ uncoded_block[332];
  wire _33955 = _152 ^ _33954;
  wire _33956 = _33953 ^ _33955;
  wire _33957 = _4840 ^ _4131;
  wire _33958 = _20048 ^ _33957;
  wire _33959 = _33956 ^ _33958;
  wire _33960 = _9790 ^ _162;
  wire _33961 = _33960 ^ _20054;
  wire _33962 = uncoded_block[377] ^ uncoded_block[385];
  wire _33963 = _6232 ^ _33962;
  wire _33964 = _13636 ^ _33963;
  wire _33965 = _33961 ^ _33964;
  wire _33966 = _33959 ^ _33965;
  wire _33967 = _33952 ^ _33966;
  wire _33968 = _28091 ^ _12541;
  wire _33969 = _12006 ^ _1048;
  wire _33970 = _33968 ^ _33969;
  wire _33971 = uncoded_block[405] ^ uncoded_block[409];
  wire _33972 = _183 ^ _33971;
  wire _33973 = _8091 ^ _1054;
  wire _33974 = _33972 ^ _33973;
  wire _33975 = _33970 ^ _33974;
  wire _33976 = _14160 ^ _8671;
  wire _33977 = _14159 ^ _33976;
  wire _33978 = _9817 ^ _28852;
  wire _33979 = _33977 ^ _33978;
  wire _33980 = _33975 ^ _33979;
  wire _33981 = _3408 ^ _11486;
  wire _33982 = _6900 ^ _6261;
  wire _33983 = _33981 ^ _33982;
  wire _33984 = _7504 ^ _8105;
  wire _33985 = _33984 ^ _26499;
  wire _33986 = _33983 ^ _33985;
  wire _33987 = uncoded_block[480] ^ uncoded_block[483];
  wire _33988 = _2657 ^ _33987;
  wire _33989 = uncoded_block[489] ^ uncoded_block[493];
  wire _33990 = _7515 ^ _33989;
  wire _33991 = _33988 ^ _33990;
  wire _33992 = _1094 ^ _1097;
  wire _33993 = _1887 ^ _1892;
  wire _33994 = _33992 ^ _33993;
  wire _33995 = _33991 ^ _33994;
  wire _33996 = _33986 ^ _33995;
  wire _33997 = _33980 ^ _33996;
  wire _33998 = _33967 ^ _33997;
  wire _33999 = _33939 ^ _33998;
  wire _34000 = _4206 ^ _13151;
  wire _34001 = _20099 ^ _6290;
  wire _34002 = _1114 ^ _4217;
  wire _34003 = _34001 ^ _34002;
  wire _34004 = _34000 ^ _34003;
  wire _34005 = _28882 ^ _6300;
  wire _34006 = _5630 ^ _3464;
  wire _34007 = _34005 ^ _34006;
  wire _34008 = _5635 ^ _25186;
  wire _34009 = _34008 ^ _33597;
  wire _34010 = _34007 ^ _34009;
  wire _34011 = _34004 ^ _34010;
  wire _34012 = _10400 ^ _24289;
  wire _34013 = uncoded_block[590] ^ uncoded_block[593];
  wire _34014 = _270 ^ _34013;
  wire _34015 = _34012 ^ _34014;
  wire _34016 = _2701 ^ _1142;
  wire _34017 = _2710 ^ _4240;
  wire _34018 = _34016 ^ _34017;
  wire _34019 = _34015 ^ _34018;
  wire _34020 = _12609 ^ _13178;
  wire _34021 = _34020 ^ _26541;
  wire _34022 = _10420 ^ _293;
  wire _34023 = _8751 ^ _296;
  wire _34024 = _34022 ^ _34023;
  wire _34025 = _34021 ^ _34024;
  wire _34026 = _34019 ^ _34025;
  wire _34027 = _34011 ^ _34026;
  wire _34028 = uncoded_block[648] ^ uncoded_block[653];
  wire _34029 = _34028 ^ _16249;
  wire _34030 = _18705 ^ _15768;
  wire _34031 = _34029 ^ _34030;
  wire _34032 = _16752 ^ _8177;
  wire _34033 = _15274 ^ _34032;
  wire _34034 = _34031 ^ _34033;
  wire _34035 = _1974 ^ _326;
  wire _34036 = _14245 ^ _34035;
  wire _34037 = _17258 ^ _3533;
  wire _34038 = _330 ^ _34037;
  wire _34039 = _34036 ^ _34038;
  wire _34040 = _34034 ^ _34039;
  wire _34041 = _3535 ^ _31525;
  wire _34042 = _1195 ^ _6367;
  wire _34043 = _34041 ^ _34042;
  wire _34044 = _21129 ^ _7001;
  wire _34045 = _31533 ^ _1203;
  wire _34046 = _34044 ^ _34045;
  wire _34047 = _34043 ^ _34046;
  wire _34048 = uncoded_block[738] ^ uncoded_block[741];
  wire _34049 = uncoded_block[744] ^ uncoded_block[751];
  wire _34050 = _34048 ^ _34049;
  wire _34051 = _34050 ^ _30233;
  wire _34052 = _9917 ^ _13766;
  wire _34053 = _366 ^ _34052;
  wire _34054 = _34051 ^ _34053;
  wire _34055 = _34047 ^ _34054;
  wire _34056 = _34040 ^ _34055;
  wire _34057 = _34027 ^ _34056;
  wire _34058 = _13768 ^ _25694;
  wire _34059 = uncoded_block[789] ^ uncoded_block[793];
  wire _34060 = _34059 ^ _6391;
  wire _34061 = _34058 ^ _34060;
  wire _34062 = uncoded_block[804] ^ uncoded_block[807];
  wire _34063 = _34062 ^ _16793;
  wire _34064 = _4318 ^ _34063;
  wire _34065 = _34061 ^ _34064;
  wire _34066 = _2026 ^ _11030;
  wire _34067 = uncoded_block[827] ^ uncoded_block[832];
  wire _34068 = _28197 ^ _34067;
  wire _34069 = _34066 ^ _34068;
  wire _34070 = _4339 ^ _9943;
  wire _34071 = _15821 ^ _34070;
  wire _34072 = _34069 ^ _34071;
  wire _34073 = _34065 ^ _34072;
  wire _34074 = _8812 ^ _2824;
  wire _34075 = _13243 ^ _34074;
  wire _34076 = _18302 ^ _1269;
  wire _34077 = _34076 ^ _27455;
  wire _34078 = _34075 ^ _34077;
  wire _34079 = uncoded_block[881] ^ uncoded_block[886];
  wire _34080 = _34079 ^ _27046;
  wire _34081 = uncoded_block[897] ^ uncoded_block[901];
  wire _34082 = _2062 ^ _34081;
  wire _34083 = _34080 ^ _34082;
  wire _34084 = _5761 ^ _12708;
  wire _34085 = _17818 ^ _18775;
  wire _34086 = _34084 ^ _34085;
  wire _34087 = _34083 ^ _34086;
  wire _34088 = _34078 ^ _34087;
  wire _34089 = _34073 ^ _34088;
  wire _34090 = _445 ^ _7075;
  wire _34091 = _34090 ^ _5097;
  wire _34092 = _5777 ^ _1303;
  wire _34093 = _27473 ^ _34092;
  wire _34094 = _34091 ^ _34093;
  wire _34095 = _10525 ^ _7680;
  wire _34096 = _4385 ^ _11646;
  wire _34097 = _34095 ^ _34096;
  wire _34098 = _2100 ^ _10537;
  wire _34099 = _28598 ^ _34098;
  wire _34100 = _34097 ^ _34099;
  wire _34101 = _34094 ^ _34100;
  wire _34102 = uncoded_block[984] ^ uncoded_block[991];
  wire _34103 = _34102 ^ _2883;
  wire _34104 = _28241 ^ _22585;
  wire _34105 = _34103 ^ _34104;
  wire _34106 = _4405 ^ _1330;
  wire _34107 = _2117 ^ _2893;
  wire _34108 = _34106 ^ _34107;
  wire _34109 = _34105 ^ _34108;
  wire _34110 = _9454 ^ _19290;
  wire _34111 = _10008 ^ _512;
  wire _34112 = _34110 ^ _34111;
  wire _34113 = _22132 ^ _19295;
  wire _34114 = _2136 ^ _7117;
  wire _34115 = _34113 ^ _34114;
  wire _34116 = _34112 ^ _34115;
  wire _34117 = _34109 ^ _34116;
  wire _34118 = _34101 ^ _34117;
  wire _34119 = _34089 ^ _34118;
  wire _34120 = _34057 ^ _34119;
  wire _34121 = _33999 ^ _34120;
  wire _34122 = uncoded_block[1066] ^ uncoded_block[1070];
  wire _34123 = _34122 ^ _527;
  wire _34124 = _32033 ^ _34123;
  wire _34125 = _3692 ^ _5834;
  wire _34126 = _7724 ^ _20753;
  wire _34127 = _34125 ^ _34126;
  wire _34128 = _34124 ^ _34127;
  wire _34129 = _4441 ^ _5844;
  wire _34130 = _2160 ^ _8336;
  wire _34131 = _29424 ^ _34130;
  wire _34132 = _34129 ^ _34131;
  wire _34133 = _34128 ^ _34132;
  wire _34134 = _5848 ^ _33312;
  wire _34135 = _31619 ^ _34134;
  wire _34136 = _18371 ^ _13866;
  wire _34137 = _34136 ^ _10035;
  wire _34138 = _34135 ^ _34137;
  wire _34139 = _3725 ^ _8354;
  wire _34140 = _10598 ^ _34139;
  wire _34141 = _6510 ^ _32884;
  wire _34142 = _2965 ^ _13339;
  wire _34143 = _34141 ^ _34142;
  wire _34144 = _34140 ^ _34143;
  wire _34145 = _34138 ^ _34144;
  wire _34146 = _34133 ^ _34145;
  wire _34147 = _29887 ^ _3746;
  wire _34148 = _12808 ^ _2971;
  wire _34149 = _34147 ^ _34148;
  wire _34150 = _26250 ^ _7758;
  wire _34151 = _2974 ^ _2217;
  wire _34152 = _34150 ^ _34151;
  wire _34153 = _34149 ^ _34152;
  wire _34154 = _27911 ^ _14914;
  wire _34155 = _5215 ^ _2988;
  wire _34156 = _34154 ^ _34155;
  wire _34157 = _2989 ^ _10067;
  wire _34158 = _1448 ^ _2997;
  wire _34159 = _34157 ^ _34158;
  wire _34160 = _34156 ^ _34159;
  wire _34161 = _34153 ^ _34160;
  wire _34162 = _6543 ^ _11739;
  wire _34163 = uncoded_block[1260] ^ uncoded_block[1264];
  wire _34164 = _5234 ^ _34163;
  wire _34165 = _34162 ^ _34164;
  wire _34166 = _10635 ^ _31239;
  wire _34167 = _34165 ^ _34166;
  wire _34168 = uncoded_block[1288] ^ uncoded_block[1292];
  wire _34169 = _638 ^ _34168;
  wire _34170 = _13376 ^ _34169;
  wire _34171 = _3018 ^ _6571;
  wire _34172 = _14428 ^ _34171;
  wire _34173 = _34170 ^ _34172;
  wire _34174 = _34167 ^ _34173;
  wire _34175 = _34161 ^ _34174;
  wire _34176 = _34146 ^ _34175;
  wire _34177 = _3807 ^ _17435;
  wire _34178 = _9552 ^ _3029;
  wire _34179 = _34177 ^ _34178;
  wire _34180 = _4543 ^ _7201;
  wire _34181 = _1490 ^ _3820;
  wire _34182 = _34180 ^ _34181;
  wire _34183 = _34179 ^ _34182;
  wire _34184 = _2276 ^ _9564;
  wire _34185 = _664 ^ _24499;
  wire _34186 = _34184 ^ _34185;
  wire _34187 = _16942 ^ _23581;
  wire _34188 = _34187 ^ _16945;
  wire _34189 = _34186 ^ _34188;
  wire _34190 = _34183 ^ _34189;
  wire _34191 = _685 ^ _3058;
  wire _34192 = _687 ^ _3061;
  wire _34193 = _34191 ^ _34192;
  wire _34194 = _4571 ^ _2296;
  wire _34195 = _693 ^ _34194;
  wire _34196 = _34193 ^ _34195;
  wire _34197 = _16954 ^ _13947;
  wire _34198 = _13418 ^ _34197;
  wire _34199 = _10683 ^ _2311;
  wire _34200 = _19399 ^ _34199;
  wire _34201 = _34198 ^ _34200;
  wire _34202 = _34196 ^ _34201;
  wire _34203 = _34190 ^ _34202;
  wire _34204 = _5968 ^ _10690;
  wire _34205 = uncoded_block[1438] ^ uncoded_block[1443];
  wire _34206 = _34205 ^ _5305;
  wire _34207 = _34204 ^ _34206;
  wire _34208 = uncoded_block[1446] ^ uncoded_block[1454];
  wire _34209 = _34208 ^ _3868;
  wire _34210 = _34209 ^ _27180;
  wire _34211 = _34207 ^ _34210;
  wire _34212 = _10136 ^ _18919;
  wire _34213 = _4603 ^ _735;
  wire _34214 = _34212 ^ _34213;
  wire _34215 = _12342 ^ _1562;
  wire _34216 = _34215 ^ _15997;
  wire _34217 = _34214 ^ _34216;
  wire _34218 = _34211 ^ _34217;
  wire _34219 = _3109 ^ _4614;
  wire _34220 = _7259 ^ _1574;
  wire _34221 = _34219 ^ _34220;
  wire _34222 = _16488 ^ _9055;
  wire _34223 = _5337 ^ _9058;
  wire _34224 = _34222 ^ _34223;
  wire _34225 = _34221 ^ _34224;
  wire _34226 = _13459 ^ _9631;
  wire _34227 = _29122 ^ _34226;
  wire _34228 = _3906 ^ _3908;
  wire _34229 = _6008 ^ _18492;
  wire _34230 = _34228 ^ _34229;
  wire _34231 = _34227 ^ _34230;
  wire _34232 = _34225 ^ _34231;
  wire _34233 = _34218 ^ _34232;
  wire _34234 = _34203 ^ _34233;
  wire _34235 = _34176 ^ _34234;
  wire _34236 = _6657 ^ _773;
  wire _34237 = uncoded_block[1565] ^ uncoded_block[1569];
  wire _34238 = _34237 ^ _4645;
  wire _34239 = _34236 ^ _34238;
  wire _34240 = uncoded_block[1579] ^ uncoded_block[1585];
  wire _34241 = _24103 ^ _34240;
  wire _34242 = _1615 ^ _3145;
  wire _34243 = _34241 ^ _34242;
  wire _34244 = _34239 ^ _34243;
  wire _34245 = _791 ^ _4654;
  wire _34246 = _13486 ^ _1621;
  wire _34247 = _34245 ^ _34246;
  wire _34248 = _1632 ^ _7911;
  wire _34249 = _20891 ^ _34248;
  wire _34250 = _34247 ^ _34249;
  wire _34251 = _34244 ^ _34250;
  wire _34252 = _3942 ^ _1639;
  wire _34253 = _9655 ^ _34252;
  wire _34254 = _23658 ^ _7306;
  wire _34255 = uncoded_block[1642] ^ uncoded_block[1645];
  wire _34256 = _2407 ^ _34255;
  wire _34257 = _34254 ^ _34256;
  wire _34258 = _34253 ^ _34257;
  wire _34259 = _822 ^ _12960;
  wire _34260 = _23224 ^ _34259;
  wire _34261 = _17537 ^ _7325;
  wire _34262 = _24585 ^ _34261;
  wire _34263 = _34260 ^ _34262;
  wire _34264 = _34258 ^ _34263;
  wire _34265 = _34251 ^ _34264;
  wire _34266 = _3967 ^ _10771;
  wire _34267 = _31764 ^ _34266;
  wire _34268 = _10212 ^ _26832;
  wire _34269 = _848 ^ _7337;
  wire _34270 = _34268 ^ _34269;
  wire _34271 = _34267 ^ _34270;
  wire _34272 = _854 ^ uncoded_block[1717];
  wire _34273 = _34271 ^ _34272;
  wire _34274 = _34265 ^ _34273;
  wire _34275 = _34235 ^ _34274;
  wire _34276 = _34121 ^ _34275;
  wire _34277 = _4711 ^ _33453;
  wire _34278 = _29179 ^ _21865;
  wire _34279 = _34277 ^ _34278;
  wire _34280 = _11344 ^ _31363;
  wire _34281 = _6095 ^ _879;
  wire _34282 = _34280 ^ _34281;
  wire _34283 = _14047 ^ _22;
  wire _34284 = _1699 ^ _5435;
  wire _34285 = _34283 ^ _34284;
  wire _34286 = _34282 ^ _34285;
  wire _34287 = _34279 ^ _34286;
  wire _34288 = _888 ^ _7364;
  wire _34289 = uncoded_block[64] ^ uncoded_block[66];
  wire _34290 = _34289 ^ _35;
  wire _34291 = _34288 ^ _34290;
  wire _34292 = _3241 ^ _900;
  wire _34293 = _6749 ^ _10249;
  wire _34294 = _34292 ^ _34293;
  wire _34295 = _34291 ^ _34294;
  wire _34296 = _14591 ^ _15097;
  wire _34297 = _15101 ^ _6120;
  wire _34298 = _34296 ^ _34297;
  wire _34299 = _9720 ^ _33056;
  wire _34300 = _12451 ^ _917;
  wire _34301 = _34299 ^ _34300;
  wire _34302 = _34298 ^ _34301;
  wire _34303 = _34295 ^ _34302;
  wire _34304 = _34287 ^ _34303;
  wire _34305 = _4754 ^ _2510;
  wire _34306 = _34305 ^ _31391;
  wire _34307 = _1744 ^ _21443;
  wire _34308 = _15118 ^ _12463;
  wire _34309 = _34307 ^ _34308;
  wire _34310 = _34306 ^ _34309;
  wire _34311 = _8589 ^ _2517;
  wire _34312 = uncoded_block[173] ^ uncoded_block[182];
  wire _34313 = _34312 ^ _4772;
  wire _34314 = _34311 ^ _34313;
  wire _34315 = _4773 ^ _3283;
  wire _34316 = _7411 ^ _16116;
  wire _34317 = _34315 ^ _34316;
  wire _34318 = _34314 ^ _34317;
  wire _34319 = _34310 ^ _34318;
  wire _34320 = uncoded_block[210] ^ uncoded_block[213];
  wire _34321 = _3291 ^ _34320;
  wire _34322 = _8019 ^ _34321;
  wire _34323 = _4787 ^ _105;
  wire _34324 = _10287 ^ _2550;
  wire _34325 = _34323 ^ _34324;
  wire _34326 = _34322 ^ _34325;
  wire _34327 = _970 ^ _1780;
  wire _34328 = _4797 ^ _8617;
  wire _34329 = _34327 ^ _34328;
  wire _34330 = _3311 ^ _8041;
  wire _34331 = _17129 ^ _34330;
  wire _34332 = _34329 ^ _34331;
  wire _34333 = _34326 ^ _34332;
  wire _34334 = _34319 ^ _34333;
  wire _34335 = _34304 ^ _34334;
  wire _34336 = _6185 ^ _984;
  wire _34337 = _34336 ^ _28060;
  wire _34338 = _3321 ^ _4103;
  wire _34339 = uncoded_block[286] ^ uncoded_block[290];
  wire _34340 = _4105 ^ _34339;
  wire _34341 = _34338 ^ _34340;
  wire _34342 = _34337 ^ _34341;
  wire _34343 = uncoded_block[304] ^ uncoded_block[308];
  wire _34344 = _4824 ^ _34343;
  wire _34345 = _10313 ^ _34344;
  wire _34346 = _8056 ^ _15671;
  wire _34347 = _4830 ^ _30116;
  wire _34348 = _34346 ^ _34347;
  wire _34349 = _34345 ^ _34348;
  wire _34350 = _34342 ^ _34349;
  wire _34351 = _4123 ^ _5534;
  wire _34352 = uncoded_block[331] ^ uncoded_block[337];
  wire _34353 = _34352 ^ _1825;
  wire _34354 = _34351 ^ _34353;
  wire _34355 = _1021 ^ _4841;
  wire _34356 = _8652 ^ _15179;
  wire _34357 = _34355 ^ _34356;
  wire _34358 = _34354 ^ _34357;
  wire _34359 = _8069 ^ _2606;
  wire _34360 = _3366 ^ _9252;
  wire _34361 = _34359 ^ _34360;
  wire _34362 = _6233 ^ _3377;
  wire _34363 = _31005 ^ _2615;
  wire _34364 = _34362 ^ _34363;
  wire _34365 = _34361 ^ _34364;
  wire _34366 = _34358 ^ _34365;
  wire _34367 = _34350 ^ _34366;
  wire _34368 = _10910 ^ _4865;
  wire _34369 = _3391 ^ _191;
  wire _34370 = _34368 ^ _34369;
  wire _34371 = _1055 ^ _7492;
  wire _34372 = _34371 ^ _31013;
  wire _34373 = _34370 ^ _34372;
  wire _34374 = _14163 ^ _2638;
  wire _34375 = uncoded_block[433] ^ uncoded_block[439];
  wire _34376 = _34375 ^ _5578;
  wire _34377 = _34374 ^ _34376;
  wire _34378 = uncoded_block[445] ^ uncoded_block[449];
  wire _34379 = _34378 ^ _4883;
  wire _34380 = _34379 ^ _4180;
  wire _34381 = _34377 ^ _34380;
  wire _34382 = _34373 ^ _34381;
  wire _34383 = _213 ^ _8105;
  wire _34384 = _1079 ^ _4186;
  wire _34385 = _34383 ^ _34384;
  wire _34386 = _1082 ^ _29702;
  wire _34387 = _5592 ^ _1086;
  wire _34388 = _34386 ^ _34387;
  wire _34389 = _34385 ^ _34388;
  wire _34390 = _4897 ^ _224;
  wire _34391 = _24727 ^ _2667;
  wire _34392 = _34390 ^ _34391;
  wire _34393 = _5611 ^ _8705;
  wire _34394 = _6286 ^ _237;
  wire _34395 = _34393 ^ _34394;
  wire _34396 = _34392 ^ _34395;
  wire _34397 = _34389 ^ _34396;
  wire _34398 = _34382 ^ _34397;
  wire _34399 = _34367 ^ _34398;
  wire _34400 = _34335 ^ _34399;
  wire _34401 = _20603 ^ _1114;
  wire _34402 = _24737 ^ _34401;
  wire _34403 = _14721 ^ _1909;
  wire _34404 = _6300 ^ _3459;
  wire _34405 = _34403 ^ _34404;
  wire _34406 = _34402 ^ _34405;
  wire _34407 = _6304 ^ _4937;
  wire _34408 = _3467 ^ _7551;
  wire _34409 = _34407 ^ _34408;
  wire _34410 = _8731 ^ _6947;
  wire _34411 = _266 ^ _3478;
  wire _34412 = _34410 ^ _34411;
  wire _34413 = _34409 ^ _34412;
  wire _34414 = _34406 ^ _34413;
  wire _34415 = _13705 ^ _6316;
  wire _34416 = _1939 ^ _15252;
  wire _34417 = _34415 ^ _34416;
  wire _34418 = _4240 ^ _8154;
  wire _34419 = _34418 ^ _7565;
  wire _34420 = _34417 ^ _34419;
  wire _34421 = _7567 ^ _6960;
  wire _34422 = _4963 ^ _2720;
  wire _34423 = _34421 ^ _34422;
  wire _34424 = _1953 ^ _290;
  wire _34425 = _34424 ^ _25654;
  wire _34426 = _34423 ^ _34425;
  wire _34427 = _34420 ^ _34426;
  wire _34428 = _34414 ^ _34427;
  wire _34429 = _296 ^ _10427;
  wire _34430 = _28528 ^ _34429;
  wire _34431 = _4262 ^ _11552;
  wire _34432 = _21112 ^ _34431;
  wire _34433 = _34430 ^ _34432;
  wire _34434 = _10442 ^ _6357;
  wire _34435 = _19680 ^ _34434;
  wire _34436 = _4272 ^ _8186;
  wire _34437 = _19195 ^ _6992;
  wire _34438 = _34436 ^ _34437;
  wire _34439 = _34435 ^ _34438;
  wire _34440 = _34433 ^ _34439;
  wire _34441 = _29330 ^ _26564;
  wire _34442 = uncoded_block[725] ^ uncoded_block[729];
  wire _34443 = _5690 ^ _34442;
  wire _34444 = _1991 ^ _3547;
  wire _34445 = _34443 ^ _34444;
  wire _34446 = _34441 ^ _34445;
  wire _34447 = uncoded_block[738] ^ uncoded_block[745];
  wire _34448 = _1995 ^ _34447;
  wire _34449 = _3554 ^ _2002;
  wire _34450 = _34448 ^ _34449;
  wire _34451 = uncoded_block[756] ^ uncoded_block[768];
  wire _34452 = _34451 ^ _7019;
  wire _34453 = _7021 ^ _12673;
  wire _34454 = _34452 ^ _34453;
  wire _34455 = _34450 ^ _34454;
  wire _34456 = _34446 ^ _34455;
  wire _34457 = _34440 ^ _34456;
  wire _34458 = _34428 ^ _34457;
  wire _34459 = _4314 ^ _14282;
  wire _34460 = _9391 ^ _34459;
  wire _34461 = _3576 ^ _4317;
  wire _34462 = uncoded_block[805] ^ uncoded_block[811];
  wire _34463 = _34462 ^ _11030;
  wire _34464 = _34461 ^ _34463;
  wire _34465 = _34460 ^ _34464;
  wire _34466 = _1241 ^ _14290;
  wire _34467 = uncoded_block[832] ^ uncoded_block[836];
  wire _34468 = _33656 ^ _34467;
  wire _34469 = _34466 ^ _34468;
  wire _34470 = uncoded_block[842] ^ uncoded_block[846];
  wire _34471 = _22532 ^ _34470;
  wire _34472 = _25711 ^ _2821;
  wire _34473 = _34471 ^ _34472;
  wire _34474 = _34469 ^ _34473;
  wire _34475 = _34465 ^ _34474;
  wire _34476 = uncoded_block[856] ^ uncoded_block[861];
  wire _34477 = _34476 ^ _29800;
  wire _34478 = _16811 ^ _416;
  wire _34479 = _34477 ^ _34478;
  wire _34480 = _15338 ^ _27044;
  wire _34481 = _34479 ^ _34480;
  wire _34482 = _14829 ^ _6424;
  wire _34483 = _12156 ^ _34482;
  wire _34484 = _9960 ^ _2850;
  wire _34485 = _34484 ^ _18313;
  wire _34486 = _34483 ^ _34485;
  wire _34487 = _34481 ^ _34486;
  wire _34488 = _34475 ^ _34487;
  wire _34489 = _6435 ^ _448;
  wire _34490 = _15351 ^ _34489;
  wire _34491 = _2078 ^ _5101;
  wire _34492 = _7673 ^ _2865;
  wire _34493 = _34491 ^ _34492;
  wire _34494 = _34490 ^ _34493;
  wire _34495 = _2086 ^ _5777;
  wire _34496 = uncoded_block[951] ^ uncoded_block[953];
  wire _34497 = _34496 ^ _461;
  wire _34498 = _34495 ^ _34497;
  wire _34499 = _463 ^ _2872;
  wire _34500 = _15363 ^ _20219;
  wire _34501 = _34499 ^ _34500;
  wire _34502 = _34498 ^ _34501;
  wire _34503 = _34494 ^ _34502;
  wire _34504 = _34098 ^ _19758;
  wire _34505 = _24858 ^ _3666;
  wire _34506 = _8294 ^ _34505;
  wire _34507 = _34504 ^ _34506;
  wire _34508 = _1338 ^ _8874;
  wire _34509 = _19290 ^ _6474;
  wire _34510 = _34508 ^ _34509;
  wire _34511 = _1336 ^ _34510;
  wire _34512 = _34507 ^ _34511;
  wire _34513 = _34503 ^ _34512;
  wire _34514 = _34488 ^ _34513;
  wire _34515 = _34458 ^ _34514;
  wire _34516 = _34400 ^ _34515;
  wire _34517 = _23956 ^ _28257;
  wire _34518 = _1360 ^ _13849;
  wire _34519 = uncoded_block[1063] ^ uncoded_block[1068];
  wire _34520 = _34519 ^ _2143;
  wire _34521 = _34518 ^ _34520;
  wire _34522 = _34517 ^ _34521;
  wire _34523 = uncoded_block[1078] ^ uncoded_block[1082];
  wire _34524 = _14361 ^ _34523;
  wire _34525 = _20253 ^ _22610;
  wire _34526 = _34524 ^ _34525;
  wire _34527 = _1378 ^ _1380;
  wire _34528 = _545 ^ _19794;
  wire _34529 = _34527 ^ _34528;
  wire _34530 = _34526 ^ _34529;
  wire _34531 = _34522 ^ _34530;
  wire _34532 = _14372 ^ _4450;
  wire _34533 = uncoded_block[1114] ^ uncoded_block[1118];
  wire _34534 = _14882 ^ _34533;
  wire _34535 = _34532 ^ _34534;
  wire _34536 = uncoded_block[1125] ^ uncoded_block[1129];
  wire _34537 = _5176 ^ _34536;
  wire _34538 = _8929 ^ _16380;
  wire _34539 = _34537 ^ _34538;
  wire _34540 = _34535 ^ _34539;
  wire _34541 = _2185 ^ _8937;
  wire _34542 = _18379 ^ _34541;
  wire _34543 = _22627 ^ _2965;
  wire _34544 = _5191 ^ _34543;
  wire _34545 = _34542 ^ _34544;
  wire _34546 = _34540 ^ _34545;
  wire _34547 = _34531 ^ _34546;
  wire _34548 = _17890 ^ _6519;
  wire _34549 = _34548 ^ _22176;
  wire _34550 = _19815 ^ _7758;
  wire _34551 = _17897 ^ _34550;
  wire _34552 = _34549 ^ _34551;
  wire _34553 = _5209 ^ _18395;
  wire _34554 = _15433 ^ _34553;
  wire _34555 = _4499 ^ _3766;
  wire _34556 = uncoded_block[1225] ^ uncoded_block[1228];
  wire _34557 = _34556 ^ _2225;
  wire _34558 = _34555 ^ _34557;
  wire _34559 = _34554 ^ _34558;
  wire _34560 = _34552 ^ _34559;
  wire _34561 = _13360 ^ _10067;
  wire _34562 = _34561 ^ _18861;
  wire _34563 = uncoded_block[1261] ^ uncoded_block[1265];
  wire _34564 = _7780 ^ _34563;
  wire _34565 = _3781 ^ _34564;
  wire _34566 = _34562 ^ _34565;
  wire _34567 = uncoded_block[1267] ^ uncoded_block[1272];
  wire _34568 = _34567 ^ _16419;
  wire _34569 = _23123 ^ _6560;
  wire _34570 = _34568 ^ _34569;
  wire _34571 = _4529 ^ _7193;
  wire _34572 = _4531 ^ _646;
  wire _34573 = _34571 ^ _34572;
  wire _34574 = _34570 ^ _34573;
  wire _34575 = _34566 ^ _34574;
  wire _34576 = _34560 ^ _34575;
  wire _34577 = _34547 ^ _34576;
  wire _34578 = _648 ^ _32506;
  wire _34579 = _34578 ^ _28668;
  wire _34580 = _21293 ^ _3029;
  wire _34581 = uncoded_block[1324] ^ uncoded_block[1330];
  wire _34582 = _34581 ^ _8413;
  wire _34583 = _34580 ^ _34582;
  wire _34584 = _34579 ^ _34583;
  wire _34585 = _3034 ^ _3822;
  wire _34586 = _34585 ^ _23578;
  wire _34587 = _12855 ^ _15473;
  wire _34588 = _673 ^ _6588;
  wire _34589 = _34587 ^ _34588;
  wire _34590 = _34586 ^ _34589;
  wire _34591 = _34584 ^ _34590;
  wire _34592 = uncoded_block[1366] ^ uncoded_block[1372];
  wire _34593 = _5275 ^ _34592;
  wire _34594 = _3058 ^ _12307;
  wire _34595 = _34593 ^ _34594;
  wire _34596 = _17953 ^ _13412;
  wire _34597 = _34596 ^ _5953;
  wire _34598 = _34595 ^ _34597;
  wire _34599 = _13939 ^ _14968;
  wire _34600 = _34599 ^ _25408;
  wire _34601 = _5962 ^ _12322;
  wire _34602 = _9588 ^ _7844;
  wire _34603 = _34601 ^ _34602;
  wire _34604 = _34600 ^ _34603;
  wire _34605 = _34598 ^ _34604;
  wire _34606 = _34591 ^ _34605;
  wire _34607 = _6613 ^ _9597;
  wire _34608 = _32950 ^ _34607;
  wire _34609 = uncoded_block[1454] ^ uncoded_block[1457];
  wire _34610 = _34609 ^ _7241;
  wire _34611 = _17474 ^ _34610;
  wire _34612 = _34608 ^ _34611;
  wire _34613 = _726 ^ _1548;
  wire _34614 = _34613 ^ _9039;
  wire _34615 = uncoded_block[1476] ^ uncoded_block[1480];
  wire _34616 = _34615 ^ _12342;
  wire _34617 = _27184 ^ _2350;
  wire _34618 = _34616 ^ _34617;
  wire _34619 = _34614 ^ _34618;
  wire _34620 = _34612 ^ _34619;
  wire _34621 = _18478 ^ _750;
  wire _34622 = _28707 ^ _34621;
  wire _34623 = uncoded_block[1512] ^ uncoded_block[1516];
  wire _34624 = _34623 ^ _9624;
  wire _34625 = _34624 ^ _29122;
  wire _34626 = _34622 ^ _34625;
  wire _34627 = _1582 ^ _6647;
  wire _34628 = _5350 ^ _5355;
  wire _34629 = _34627 ^ _34628;
  wire _34630 = _28378 ^ _11281;
  wire _34631 = _19438 ^ _34630;
  wire _34632 = _34629 ^ _34631;
  wire _34633 = _34626 ^ _34632;
  wire _34634 = _34620 ^ _34633;
  wire _34635 = _34606 ^ _34634;
  wire _34636 = _34577 ^ _34635;
  wire _34637 = _25894 ^ _30870;
  wire _34638 = _2380 ^ _1612;
  wire _34639 = _34637 ^ _34638;
  wire _34640 = _2386 ^ _3145;
  wire _34641 = _14512 ^ _8499;
  wire _34642 = _34640 ^ _34641;
  wire _34643 = _34639 ^ _34642;
  wire _34644 = _6039 ^ _6677;
  wire _34645 = _4662 ^ _20409;
  wire _34646 = _34644 ^ _34645;
  wire _34647 = _9096 ^ _10748;
  wire _34648 = _34646 ^ _34647;
  wire _34649 = _34643 ^ _34648;
  wire _34650 = _1636 ^ _7305;
  wire _34651 = _7308 ^ _1646;
  wire _34652 = _34650 ^ _34651;
  wire _34653 = _1650 ^ _15048;
  wire _34654 = _16049 ^ _25476;
  wire _34655 = _34653 ^ _34654;
  wire _34656 = _34652 ^ _34655;
  wire _34657 = _830 ^ _3962;
  wire _34658 = _20427 ^ _13517;
  wire _34659 = _34657 ^ _34658;
  wire _34660 = _3965 ^ _3189;
  wire _34661 = _3968 ^ _29162;
  wire _34662 = _34660 ^ _34661;
  wire _34663 = _34659 ^ _34662;
  wire _34664 = _34656 ^ _34663;
  wire _34665 = _34649 ^ _34664;
  wire _34666 = _6068 ^ _8535;
  wire _34667 = _34666 ^ _27672;
  wire _34668 = _7944 ^ uncoded_block[1719];
  wire _34669 = _34667 ^ _34668;
  wire _34670 = _34665 ^ _34669;
  wire _34671 = _34636 ^ _34670;
  wire _34672 = _34516 ^ _34671;
  wire _34673 = _1 ^ _3;
  wire _34674 = _2454 ^ _7956;
  wire _34675 = _34673 ^ _34674;
  wire _34676 = uncoded_block[15] ^ uncoded_block[19];
  wire _34677 = _34676 ^ _9694;
  wire _34678 = _11344 ^ _8548;
  wire _34679 = _34677 ^ _34678;
  wire _34680 = _34675 ^ _34679;
  wire _34681 = _30043 ^ _21877;
  wire _34682 = uncoded_block[52] ^ uncoded_block[55];
  wire _34683 = _1699 ^ _34682;
  wire _34684 = _1703 ^ _31;
  wire _34685 = _34683 ^ _34684;
  wire _34686 = _34681 ^ _34685;
  wire _34687 = _34680 ^ _34686;
  wire _34688 = uncoded_block[64] ^ uncoded_block[67];
  wire _34689 = uncoded_block[72] ^ uncoded_block[77];
  wire _34690 = _34688 ^ _34689;
  wire _34691 = _2481 ^ _19019;
  wire _34692 = _34690 ^ _34691;
  wire _34693 = _6754 ^ _9713;
  wire _34694 = uncoded_block[96] ^ uncoded_block[103];
  wire _34695 = _19515 ^ _34694;
  wire _34696 = _34693 ^ _34695;
  wire _34697 = _34692 ^ _34696;
  wire _34698 = uncoded_block[106] ^ uncoded_block[114];
  wire _34699 = _34698 ^ _33056;
  wire _34700 = _34699 ^ _32631;
  wire _34701 = _25523 ^ _33065;
  wire _34702 = _34700 ^ _34701;
  wire _34703 = _34697 ^ _34702;
  wire _34704 = _34687 ^ _34703;
  wire _34705 = _64 ^ _11918;
  wire _34706 = _16600 ^ _9182;
  wire _34707 = _34705 ^ _34706;
  wire _34708 = _70 ^ _7397;
  wire _34709 = uncoded_block[158] ^ uncoded_block[164];
  wire _34710 = _1748 ^ _34709;
  wire _34711 = _34708 ^ _34710;
  wire _34712 = _34707 ^ _34711;
  wire _34713 = _19539 ^ _6149;
  wire _34714 = _33073 ^ _34713;
  wire _34715 = _85 ^ _11395;
  wire _34716 = _16114 ^ _6798;
  wire _34717 = _34715 ^ _34716;
  wire _34718 = _34714 ^ _34717;
  wire _34719 = _34712 ^ _34718;
  wire _34720 = _89 ^ _5485;
  wire _34721 = _95 ^ _29634;
  wire _34722 = _34720 ^ _34721;
  wire _34723 = _8600 ^ _4785;
  wire _34724 = uncoded_block[223] ^ uncoded_block[226];
  wire _34725 = _14105 ^ _34724;
  wire _34726 = _34723 ^ _34725;
  wire _34727 = _34722 ^ _34726;
  wire _34728 = _4791 ^ _2550;
  wire _34729 = _34728 ^ _25552;
  wire _34730 = _11954 ^ _2557;
  wire _34731 = _32662 ^ _34730;
  wire _34732 = _34729 ^ _34731;
  wire _34733 = _34727 ^ _34732;
  wire _34734 = _34719 ^ _34733;
  wire _34735 = _34704 ^ _34734;
  wire _34736 = _9761 ^ _33510;
  wire _34737 = _34736 ^ _19064;
  wire _34738 = _1793 ^ _10300;
  wire _34739 = _26443 ^ _34738;
  wire _34740 = _34737 ^ _34739;
  wire _34741 = _8632 ^ _11429;
  wire _34742 = _11968 ^ _34741;
  wire _34743 = _4819 ^ _138;
  wire _34744 = uncoded_block[301] ^ uncoded_block[306];
  wire _34745 = _34744 ^ _3334;
  wire _34746 = _34743 ^ _34745;
  wire _34747 = _34742 ^ _34746;
  wire _34748 = _34740 ^ _34747;
  wire _34749 = _15670 ^ _9233;
  wire _34750 = _34749 ^ _1010;
  wire _34751 = uncoded_block[330] ^ uncoded_block[335];
  wire _34752 = _30117 ^ _34751;
  wire _34753 = _10323 ^ _32687;
  wire _34754 = _34752 ^ _34753;
  wire _34755 = _34750 ^ _34754;
  wire _34756 = _168 ^ _13094;
  wire _34757 = _22878 ^ _34756;
  wire _34758 = _9798 ^ _6235;
  wire _34759 = _1039 ^ _28091;
  wire _34760 = _34758 ^ _34759;
  wire _34761 = _34757 ^ _34760;
  wire _34762 = _34755 ^ _34761;
  wire _34763 = _34748 ^ _34762;
  wire _34764 = _26042 ^ _4155;
  wire _34765 = _11468 ^ _34764;
  wire _34766 = uncoded_block[409] ^ uncoded_block[412];
  wire _34767 = _184 ^ _34766;
  wire _34768 = _8092 ^ _11477;
  wire _34769 = _34767 ^ _34768;
  wire _34770 = _34765 ^ _34769;
  wire _34771 = uncoded_block[428] ^ uncoded_block[432];
  wire _34772 = _34771 ^ _7497;
  wire _34773 = _3405 ^ _3409;
  wire _34774 = _34772 ^ _34773;
  wire _34775 = _1075 ^ _10926;
  wire _34776 = _4185 ^ _8683;
  wire _34777 = _34775 ^ _34776;
  wire _34778 = _34774 ^ _34777;
  wire _34779 = _34770 ^ _34778;
  wire _34780 = _14175 ^ _29280;
  wire _34781 = _4192 ^ _10368;
  wire _34782 = _34780 ^ _34781;
  wire _34783 = uncoded_block[488] ^ uncoded_block[491];
  wire _34784 = _7515 ^ _34783;
  wire _34785 = uncoded_block[495] ^ uncoded_block[498];
  wire _34786 = _34785 ^ _1097;
  wire _34787 = _34784 ^ _34786;
  wire _34788 = _34782 ^ _34787;
  wire _34789 = uncoded_block[502] ^ uncoded_block[507];
  wire _34790 = _34789 ^ _4205;
  wire _34791 = _15220 ^ _4910;
  wire _34792 = _34790 ^ _34791;
  wire _34793 = _1900 ^ _12039;
  wire _34794 = _28124 ^ _34793;
  wire _34795 = _34792 ^ _34794;
  wire _34796 = _34788 ^ _34795;
  wire _34797 = _34779 ^ _34796;
  wire _34798 = _34763 ^ _34797;
  wire _34799 = _34735 ^ _34798;
  wire _34800 = _24279 ^ _7540;
  wire _34801 = _10959 ^ _1913;
  wire _34802 = _34800 ^ _34801;
  wire _34803 = _1915 ^ _12051;
  wire _34804 = _32736 ^ _8727;
  wire _34805 = _34803 ^ _34804;
  wire _34806 = _34802 ^ _34805;
  wire _34807 = _11526 ^ _2696;
  wire _34808 = _34807 ^ _14734;
  wire _34809 = _6952 ^ _3486;
  wire _34810 = _10406 ^ _34809;
  wire _34811 = _34808 ^ _34810;
  wire _34812 = _34806 ^ _34811;
  wire _34813 = _3487 ^ _8152;
  wire _34814 = _16233 ^ _7563;
  wire _34815 = _34813 ^ _34814;
  wire _34816 = _1149 ^ _4960;
  wire _34817 = _4963 ^ _7570;
  wire _34818 = _34816 ^ _34817;
  wire _34819 = _34815 ^ _34818;
  wire _34820 = _2722 ^ _6330;
  wire _34821 = uncoded_block[635] ^ uncoded_block[639];
  wire _34822 = _34821 ^ _1163;
  wire _34823 = _34820 ^ _34822;
  wire _34824 = _297 ^ _1960;
  wire _34825 = _32754 ^ _34824;
  wire _34826 = _34823 ^ _34825;
  wire _34827 = _34819 ^ _34826;
  wire _34828 = _34812 ^ _34827;
  wire _34829 = uncoded_block[654] ^ uncoded_block[659];
  wire _34830 = _34829 ^ _5670;
  wire _34831 = _5671 ^ _2744;
  wire _34832 = _34830 ^ _34831;
  wire _34833 = _17745 ^ _8177;
  wire _34834 = uncoded_block[684] ^ uncoded_block[688];
  wire _34835 = _1971 ^ _34834;
  wire _34836 = _34833 ^ _34835;
  wire _34837 = _34832 ^ _34836;
  wire _34838 = _11556 ^ _328;
  wire _34839 = _34838 ^ _17256;
  wire _34840 = uncoded_block[701] ^ uncoded_block[704];
  wire _34841 = _34840 ^ _7597;
  wire _34842 = _32772 ^ _1984;
  wire _34843 = _34841 ^ _34842;
  wire _34844 = _34839 ^ _34843;
  wire _34845 = _34837 ^ _34844;
  wire _34846 = _9904 ^ _344;
  wire _34847 = _8200 ^ _23870;
  wire _34848 = _34846 ^ _34847;
  wire _34849 = uncoded_block[748] ^ uncoded_block[751];
  wire _34850 = _34849 ^ _1214;
  wire _34851 = _9373 ^ _34850;
  wire _34852 = _34848 ^ _34851;
  wire _34853 = _29773 ^ _18270;
  wire _34854 = _13762 ^ _1218;
  wire _34855 = uncoded_block[771] ^ uncoded_block[774];
  wire _34856 = _34855 ^ _3562;
  wire _34857 = _34854 ^ _34856;
  wire _34858 = _34853 ^ _34857;
  wire _34859 = _34852 ^ _34858;
  wire _34860 = _34845 ^ _34859;
  wire _34861 = _34828 ^ _34860;
  wire _34862 = uncoded_block[777] ^ uncoded_block[781];
  wire _34863 = _34862 ^ _3570;
  wire _34864 = _5032 ^ _4314;
  wire _34865 = _34863 ^ _34864;
  wire _34866 = _8224 ^ _1235;
  wire _34867 = _15814 ^ _2806;
  wire _34868 = _34866 ^ _34867;
  wire _34869 = _34865 ^ _34868;
  wire _34870 = _22525 ^ _7037;
  wire _34871 = _3587 ^ _1249;
  wire _34872 = _34870 ^ _34871;
  wire _34873 = _34467 ^ _2035;
  wire _34874 = _34873 ^ _24816;
  wire _34875 = _34872 ^ _34874;
  wire _34876 = _34869 ^ _34875;
  wire _34877 = _9945 ^ _23010;
  wire _34878 = _2045 ^ _34877;
  wire _34879 = _14302 ^ _1266;
  wire _34880 = _5072 ^ _1269;
  wire _34881 = _34879 ^ _34880;
  wire _34882 = _34878 ^ _34881;
  wire _34883 = uncoded_block[879] ^ uncoded_block[885];
  wire _34884 = _417 ^ _34883;
  wire _34885 = _11059 ^ _9416;
  wire _34886 = _34884 ^ _34885;
  wire _34887 = _29808 ^ _429;
  wire _34888 = _34887 ^ _17315;
  wire _34889 = _34886 ^ _34888;
  wire _34890 = _34882 ^ _34889;
  wire _34891 = _34876 ^ _34890;
  wire _34892 = _15349 ^ _32823;
  wire _34893 = _16827 ^ _1296;
  wire _34894 = _1294 ^ _34893;
  wire _34895 = _34892 ^ _34894;
  wire _34896 = _5096 ^ _1299;
  wire _34897 = _4377 ^ _8271;
  wire _34898 = _34896 ^ _34897;
  wire _34899 = _456 ^ _13266;
  wire _34900 = _34899 ^ _34497;
  wire _34901 = _34898 ^ _34900;
  wire _34902 = _34895 ^ _34901;
  wire _34903 = _10528 ^ _11086;
  wire _34904 = _11648 ^ _8283;
  wire _34905 = _34903 ^ _34904;
  wire _34906 = uncoded_block[977] ^ uncoded_block[984];
  wire _34907 = _34906 ^ _8856;
  wire _34908 = _8859 ^ _4401;
  wire _34909 = _34907 ^ _34908;
  wire _34910 = _34905 ^ _34909;
  wire _34911 = _2107 ^ _4404;
  wire _34912 = _27488 ^ _34911;
  wire _34913 = uncoded_block[1005] ^ uncoded_block[1010];
  wire _34914 = _34913 ^ _19763;
  wire _34915 = uncoded_block[1018] ^ uncoded_block[1023];
  wire _34916 = _34915 ^ _12752;
  wire _34917 = _34914 ^ _34916;
  wire _34918 = _34912 ^ _34917;
  wire _34919 = _34910 ^ _34918;
  wire _34920 = _34902 ^ _34919;
  wire _34921 = _34891 ^ _34920;
  wire _34922 = _34861 ^ _34921;
  wire _34923 = _34799 ^ _34922;
  wire _34924 = _498 ^ _4417;
  wire _34925 = uncoded_block[1032] ^ uncoded_block[1035];
  wire _34926 = _34925 ^ _1345;
  wire _34927 = _34924 ^ _34926;
  wire _34928 = _1346 ^ _16864;
  wire _34929 = _34928 ^ _1358;
  wire _34930 = _34927 ^ _34929;
  wire _34931 = _5147 ^ _519;
  wire _34932 = _6483 ^ _522;
  wire _34933 = _34931 ^ _34932;
  wire _34934 = uncoded_block[1069] ^ uncoded_block[1074];
  wire _34935 = _34934 ^ _2924;
  wire _34936 = _3690 ^ _34935;
  wire _34937 = _34933 ^ _34936;
  wire _34938 = _34930 ^ _34937;
  wire _34939 = _2925 ^ _8904;
  wire _34940 = _15401 ^ _537;
  wire _34941 = _34939 ^ _34940;
  wire _34942 = _542 ^ _11139;
  wire _34943 = uncoded_block[1104] ^ uncoded_block[1107];
  wire _34944 = _4444 ^ _34943;
  wire _34945 = _34942 ^ _34944;
  wire _34946 = _34941 ^ _34945;
  wire _34947 = _2938 ^ _8920;
  wire _34948 = _4452 ^ _34947;
  wire _34949 = uncoded_block[1123] ^ uncoded_block[1127];
  wire _34950 = _4455 ^ _34949;
  wire _34951 = _8343 ^ _2950;
  wire _34952 = _34950 ^ _34951;
  wire _34953 = _34948 ^ _34952;
  wire _34954 = _34946 ^ _34953;
  wire _34955 = _34938 ^ _34954;
  wire _34956 = _568 ^ _3724;
  wire _34957 = _34956 ^ _34541;
  wire _34958 = _2188 ^ _3736;
  wire _34959 = _34958 ^ _29033;
  wire _34960 = _34957 ^ _34959;
  wire _34961 = uncoded_block[1177] ^ uncoded_block[1181];
  wire _34962 = _585 ^ _34961;
  wire _34963 = _592 ^ _12808;
  wire _34964 = _34962 ^ _34963;
  wire _34965 = _2971 ^ _4488;
  wire _34966 = _13886 ^ _5207;
  wire _34967 = _34965 ^ _34966;
  wire _34968 = _34964 ^ _34967;
  wire _34969 = _34960 ^ _34968;
  wire _34970 = _11171 ^ _26694;
  wire _34971 = _5889 ^ _608;
  wire _34972 = _34970 ^ _34971;
  wire _34973 = _609 ^ _11177;
  wire _34974 = _34973 ^ _32901;
  wire _34975 = _34972 ^ _34974;
  wire _34976 = _29899 ^ _2997;
  wire _34977 = _2998 ^ _11739;
  wire _34978 = _34976 ^ _34977;
  wire _34979 = _24926 ^ _6551;
  wire _34980 = _34978 ^ _34979;
  wire _34981 = _34975 ^ _34980;
  wire _34982 = _34969 ^ _34981;
  wire _34983 = _34955 ^ _34982;
  wire _34984 = _9532 ^ _11746;
  wire _34985 = _630 ^ _3793;
  wire _34986 = _34984 ^ _34985;
  wire _34987 = uncoded_block[1283] ^ uncoded_block[1291];
  wire _34988 = _3794 ^ _34987;
  wire _34989 = _30797 ^ _4531;
  wire _34990 = _34988 ^ _34989;
  wire _34991 = _34986 ^ _34990;
  wire _34992 = uncoded_block[1304] ^ uncoded_block[1309];
  wire _34993 = _6564 ^ _34992;
  wire _34994 = _11759 ^ _21293;
  wire _34995 = _34993 ^ _34994;
  wire _34996 = uncoded_block[1322] ^ uncoded_block[1325];
  wire _34997 = _9555 ^ _34996;
  wire _34998 = _34997 ^ _30806;
  wire _34999 = _34995 ^ _34998;
  wire _35000 = _34991 ^ _34999;
  wire _35001 = _21753 ^ _9563;
  wire _35002 = _16938 ^ _1498;
  wire _35003 = _35001 ^ _35002;
  wire _35004 = _664 ^ _18434;
  wire _35005 = _35004 ^ _14448;
  wire _35006 = _35003 ^ _35005;
  wire _35007 = _21762 ^ _3052;
  wire _35008 = _35007 ^ _8424;
  wire _35009 = uncoded_block[1379] ^ uncoded_block[1383];
  wire _35010 = _3055 ^ _35009;
  wire _35011 = _25399 ^ _24511;
  wire _35012 = _35010 ^ _35011;
  wire _35013 = _35008 ^ _35012;
  wire _35014 = _35006 ^ _35013;
  wire _35015 = _35000 ^ _35014;
  wire _35016 = uncoded_block[1395] ^ uncoded_block[1399];
  wire _35017 = _5952 ^ _35016;
  wire _35018 = _3841 ^ _3846;
  wire _35019 = _35017 ^ _35018;
  wire _35020 = _702 ^ _32942;
  wire _35021 = _9586 ^ _35020;
  wire _35022 = _35019 ^ _35021;
  wire _35023 = _4586 ^ _712;
  wire _35024 = _32949 ^ _35023;
  wire _35025 = _6613 ^ _9033;
  wire _35026 = _26309 ^ _6622;
  wire _35027 = _35025 ^ _35026;
  wire _35028 = _35024 ^ _35027;
  wire _35029 = _35022 ^ _35028;
  wire _35030 = _2329 ^ _3870;
  wire _35031 = _3094 ^ _29519;
  wire _35032 = _35030 ^ _35031;
  wire _35033 = _733 ^ _13446;
  wire _35034 = uncoded_block[1480] ^ uncoded_block[1488];
  wire _35035 = _35034 ^ _15996;
  wire _35036 = _35033 ^ _35035;
  wire _35037 = _35032 ^ _35036;
  wire _35038 = _5333 ^ _7875;
  wire _35039 = _32965 ^ _35038;
  wire _35040 = _11267 ^ _15004;
  wire _35041 = _35040 ^ _32969;
  wire _35042 = _35039 ^ _35041;
  wire _35043 = _35037 ^ _35042;
  wire _35044 = _35029 ^ _35043;
  wire _35045 = _35015 ^ _35044;
  wire _35046 = _34983 ^ _35045;
  wire _35047 = _15009 ^ _5350;
  wire _35048 = _32972 ^ _35047;
  wire _35049 = _2368 ^ _19438;
  wire _35050 = _35048 ^ _35049;
  wire _35051 = _7885 ^ _770;
  wire _35052 = _35051 ^ _21357;
  wire _35053 = _4644 ^ _5363;
  wire _35054 = _9080 ^ _782;
  wire _35055 = _35053 ^ _35054;
  wire _35056 = _35052 ^ _35055;
  wire _35057 = _35050 ^ _35056;
  wire _35058 = _3145 ^ _19448;
  wire _35059 = _13481 ^ _35058;
  wire _35060 = _3934 ^ _9088;
  wire _35061 = _5380 ^ _12940;
  wire _35062 = _35060 ^ _35061;
  wire _35063 = _35059 ^ _35062;
  wire _35064 = uncoded_block[1625] ^ uncoded_block[1629];
  wire _35065 = _3941 ^ _35064;
  wire _35066 = _30879 ^ _35065;
  wire _35067 = _2405 ^ _7308;
  wire _35068 = _1640 ^ _35067;
  wire _35069 = _35066 ^ _35068;
  wire _35070 = _35063 ^ _35069;
  wire _35071 = _35057 ^ _35070;
  wire _35072 = _6689 ^ _5394;
  wire _35073 = uncoded_block[1647] ^ uncoded_block[1652];
  wire _35074 = _35073 ^ _8515;
  wire _35075 = _35072 ^ _35074;
  wire _35076 = uncoded_block[1664] ^ uncoded_block[1669];
  wire _35077 = _20909 ^ _35076;
  wire _35078 = _22763 ^ _31339;
  wire _35079 = _35077 ^ _35078;
  wire _35080 = _35075 ^ _35079;
  wire _35081 = uncoded_block[1680] ^ uncoded_block[1684];
  wire _35082 = _35081 ^ _7331;
  wire _35083 = _840 ^ _25037;
  wire _35084 = _35082 ^ _35083;
  wire _35085 = _24138 ^ _33022;
  wire _35086 = _35084 ^ _35085;
  wire _35087 = _35080 ^ _35086;
  wire _35088 = _7944 ^ _860;
  wire _35089 = _35088 ^ uncoded_block[1722];
  wire _35090 = _35087 ^ _35089;
  wire _35091 = _35071 ^ _35090;
  wire _35092 = _35046 ^ _35091;
  wire _35093 = _34923 ^ _35092;
  wire _35094 = _15073 ^ _1686;
  wire _35095 = _4711 ^ _35094;
  wire _35096 = uncoded_block[23] ^ uncoded_block[27];
  wire _35097 = _19496 ^ _35096;
  wire _35098 = _14041 ^ _35097;
  wire _35099 = _35095 ^ _35098;
  wire _35100 = _874 ^ _15;
  wire _35101 = _16 ^ _15590;
  wire _35102 = _35100 ^ _35101;
  wire _35103 = uncoded_block[44] ^ uncoded_block[50];
  wire _35104 = _20457 ^ _35103;
  wire _35105 = _34682 ^ _23256;
  wire _35106 = _35104 ^ _35105;
  wire _35107 = _35102 ^ _35106;
  wire _35108 = _35099 ^ _35107;
  wire _35109 = _11355 ^ _6744;
  wire _35110 = _35109 ^ _17576;
  wire _35111 = uncoded_block[81] ^ uncoded_block[84];
  wire _35112 = _3243 ^ _35111;
  wire _35113 = uncoded_block[94] ^ uncoded_block[100];
  wire _35114 = _7981 ^ _35113;
  wire _35115 = _35112 ^ _35114;
  wire _35116 = _35110 ^ _35115;
  wire _35117 = uncoded_block[113] ^ uncoded_block[120];
  wire _35118 = _9720 ^ _35117;
  wire _35119 = _34297 ^ _35118;
  wire _35120 = _10256 ^ _917;
  wire _35121 = uncoded_block[136] ^ uncoded_block[140];
  wire _35122 = _4754 ^ _35121;
  wire _35123 = _35120 ^ _35122;
  wire _35124 = _35119 ^ _35123;
  wire _35125 = _35116 ^ _35124;
  wire _35126 = _35108 ^ _35125;
  wire _35127 = _15114 ^ _1744;
  wire _35128 = _21443 ^ _15118;
  wire _35129 = _35127 ^ _35128;
  wire _35130 = uncoded_block[167] ^ uncoded_block[173];
  wire _35131 = _35130 ^ _4772;
  wire _35132 = _28031 ^ _35131;
  wire _35133 = _35129 ^ _35132;
  wire _35134 = uncoded_block[206] ^ uncoded_block[213];
  wire _35135 = _12479 ^ _35134;
  wire _35136 = uncoded_block[219] ^ uncoded_block[223];
  wire _35137 = _8606 ^ _35136;
  wire _35138 = _35135 ^ _35137;
  wire _35139 = _30081 ^ _35138;
  wire _35140 = _35133 ^ _35139;
  wire _35141 = uncoded_block[234] ^ uncoded_block[237];
  wire _35142 = _29225 ^ _35141;
  wire _35143 = _19057 ^ _35142;
  wire _35144 = _5500 ^ _10860;
  wire _35145 = uncoded_block[244] ^ uncoded_block[247];
  wire _35146 = _35145 ^ _2556;
  wire _35147 = _35144 ^ _35146;
  wire _35148 = _35143 ^ _35147;
  wire _35149 = _4803 ^ _9761;
  wire _35150 = _35149 ^ _6828;
  wire _35151 = _21932 ^ _985;
  wire _35152 = _35151 ^ _25116;
  wire _35153 = _35150 ^ _35152;
  wire _35154 = _35148 ^ _35153;
  wire _35155 = _35140 ^ _35154;
  wire _35156 = _35126 ^ _35155;
  wire _35157 = uncoded_block[284] ^ uncoded_block[290];
  wire _35158 = _1796 ^ _35157;
  wire _35159 = uncoded_block[291] ^ uncoded_block[297];
  wire _35160 = _35159 ^ _2577;
  wire _35161 = _35158 ^ _35160;
  wire _35162 = _34343 ^ _8056;
  wire _35163 = _35162 ^ _30987;
  wire _35164 = _35161 ^ _35163;
  wire _35165 = uncoded_block[322] ^ uncoded_block[330];
  wire _35166 = _4832 ^ _35165;
  wire _35167 = _24685 ^ _4840;
  wire _35168 = _35166 ^ _35167;
  wire _35169 = _3355 ^ _4845;
  wire _35170 = uncoded_block[359] ^ uncoded_block[362];
  wire _35171 = _13089 ^ _35170;
  wire _35172 = _35169 ^ _35171;
  wire _35173 = _35168 ^ _35172;
  wire _35174 = _35164 ^ _35173;
  wire _35175 = uncoded_block[364] ^ uncoded_block[375];
  wire _35176 = _35175 ^ _6233;
  wire _35177 = _35176 ^ _10337;
  wire _35178 = _176 ^ _14678;
  wire _35179 = _1849 ^ _8088;
  wire _35180 = _35178 ^ _35179;
  wire _35181 = _35177 ^ _35180;
  wire _35182 = _1052 ^ _9266;
  wire _35183 = _5565 ^ _14160;
  wire _35184 = _35182 ^ _35183;
  wire _35185 = _1060 ^ _1062;
  wire _35186 = _35185 ^ _23792;
  wire _35187 = _35184 ^ _35186;
  wire _35188 = _35181 ^ _35187;
  wire _35189 = _35174 ^ _35188;
  wire _35190 = _201 ^ _19115;
  wire _35191 = _206 ^ _34378;
  wire _35192 = _35190 ^ _35191;
  wire _35193 = _4883 ^ _1075;
  wire _35194 = _35193 ^ _214;
  wire _35195 = _35192 ^ _35194;
  wire _35196 = _1873 ^ _8683;
  wire _35197 = _35196 ^ _4892;
  wire _35198 = _29702 ^ _8693;
  wire _35199 = _15212 ^ _1090;
  wire _35200 = _35198 ^ _35199;
  wire _35201 = _35197 ^ _35200;
  wire _35202 = _35195 ^ _35201;
  wire _35203 = _5600 ^ _4903;
  wire _35204 = _35203 ^ _34790;
  wire _35205 = _9298 ^ _19638;
  wire _35206 = _13152 ^ _4921;
  wire _35207 = _35205 ^ _35206;
  wire _35208 = _35204 ^ _35207;
  wire _35209 = _9310 ^ _16714;
  wire _35210 = _14725 ^ _8721;
  wire _35211 = _5629 ^ _35210;
  wire _35212 = _35209 ^ _35211;
  wire _35213 = _35208 ^ _35212;
  wire _35214 = _35202 ^ _35213;
  wire _35215 = _35189 ^ _35214;
  wire _35216 = _35156 ^ _35215;
  wire _35217 = _12051 ^ _3467;
  wire _35218 = _3472 ^ _10967;
  wire _35219 = _35217 ^ _35218;
  wire _35220 = uncoded_block[585] ^ uncoded_block[588];
  wire _35221 = _5641 ^ _35220;
  wire _35222 = uncoded_block[591] ^ uncoded_block[594];
  wire _35223 = _35222 ^ _1939;
  wire _35224 = _35221 ^ _35223;
  wire _35225 = _35219 ^ _35224;
  wire _35226 = _15252 ^ _4240;
  wire _35227 = _35226 ^ _16237;
  wire _35228 = uncoded_block[623] ^ uncoded_block[627];
  wire _35229 = _7568 ^ _35228;
  wire _35230 = _12070 ^ _35229;
  wire _35231 = _35227 ^ _35230;
  wire _35232 = _35225 ^ _35231;
  wire _35233 = _34424 ^ _24304;
  wire _35234 = _19177 ^ _304;
  wire _35235 = _14749 ^ _35234;
  wire _35236 = _35233 ^ _35235;
  wire _35237 = _308 ^ _11552;
  wire _35238 = _3515 ^ _35237;
  wire _35239 = _6353 ^ _10442;
  wire _35240 = _6357 ^ _9895;
  wire _35241 = _35239 ^ _35240;
  wire _35242 = _35238 ^ _35241;
  wire _35243 = _35236 ^ _35242;
  wire _35244 = _35232 ^ _35243;
  wire _35245 = _20654 ^ _19688;
  wire _35246 = _16760 ^ _35245;
  wire _35247 = uncoded_block[716] ^ uncoded_block[719];
  wire _35248 = _337 ^ _35247;
  wire _35249 = _18259 ^ _7603;
  wire _35250 = _35248 ^ _35249;
  wire _35251 = _35246 ^ _35250;
  wire _35252 = _1996 ^ _3554;
  wire _35253 = _25681 ^ _35252;
  wire _35254 = uncoded_block[751] ^ uncoded_block[756];
  wire _35255 = uncoded_block[757] ^ uncoded_block[768];
  wire _35256 = _35254 ^ _35255;
  wire _35257 = uncoded_block[772] ^ uncoded_block[778];
  wire _35258 = _35257 ^ _3568;
  wire _35259 = _35256 ^ _35258;
  wire _35260 = _35253 ^ _35259;
  wire _35261 = _35251 ^ _35260;
  wire _35262 = _3570 ^ _1224;
  wire _35263 = _35262 ^ _5722;
  wire _35264 = _2799 ^ _3576;
  wire _35265 = _4317 ^ _389;
  wire _35266 = _35264 ^ _35265;
  wire _35267 = _35263 ^ _35266;
  wire _35268 = uncoded_block[806] ^ uncoded_block[811];
  wire _35269 = _35268 ^ _5046;
  wire _35270 = _12131 ^ _14290;
  wire _35271 = _35269 ^ _35270;
  wire _35272 = _22532 ^ _10495;
  wire _35273 = _34468 ^ _35272;
  wire _35274 = _35271 ^ _35273;
  wire _35275 = _35267 ^ _35274;
  wire _35276 = _35261 ^ _35275;
  wire _35277 = _35244 ^ _35276;
  wire _35278 = _13238 ^ _6406;
  wire _35279 = _35278 ^ _32809;
  wire _35280 = _9948 ^ _2827;
  wire _35281 = uncoded_block[870] ^ uncoded_block[872];
  wire _35282 = _35281 ^ _2831;
  wire _35283 = _35280 ^ _35282;
  wire _35284 = _35279 ^ _35283;
  wire _35285 = _420 ^ _2054;
  wire _35286 = _35285 ^ _2060;
  wire _35287 = uncoded_block[890] ^ uncoded_block[895];
  wire _35288 = _35287 ^ _1278;
  wire _35289 = uncoded_block[904] ^ uncoded_block[909];
  wire _35290 = _10508 ^ _35289;
  wire _35291 = _35288 ^ _35290;
  wire _35292 = _35286 ^ _35291;
  wire _35293 = _35284 ^ _35292;
  wire _35294 = _7665 ^ _436;
  wire _35295 = _35294 ^ _22555;
  wire _35296 = uncoded_block[923] ^ uncoded_block[930];
  wire _35297 = _35296 ^ _5096;
  wire _35298 = _25736 ^ _7080;
  wire _35299 = _35297 ^ _35298;
  wire _35300 = _35295 ^ _35299;
  wire _35301 = _1300 ^ _2086;
  wire _35302 = _5777 ^ _8275;
  wire _35303 = _35301 ^ _35302;
  wire _35304 = _4384 ^ _10531;
  wire _35305 = _8847 ^ _3657;
  wire _35306 = _35304 ^ _35305;
  wire _35307 = _35303 ^ _35306;
  wire _35308 = _35300 ^ _35307;
  wire _35309 = _35293 ^ _35308;
  wire _35310 = _7689 ^ _8856;
  wire _35311 = _4396 ^ _35310;
  wire _35312 = _10543 ^ _11101;
  wire _35313 = _2107 ^ _20730;
  wire _35314 = _35312 ^ _35313;
  wire _35315 = _35311 ^ _35314;
  wire _35316 = _4409 ^ _491;
  wire _35317 = _11663 ^ _2120;
  wire _35318 = _35316 ^ _35317;
  wire _35319 = _5137 ^ _12752;
  wire _35320 = uncoded_block[1029] ^ uncoded_block[1033];
  wire _35321 = _498 ^ _35320;
  wire _35322 = _35319 ^ _35321;
  wire _35323 = _35318 ^ _35322;
  wire _35324 = _35315 ^ _35323;
  wire _35325 = _6474 ^ _512;
  wire _35326 = _35325 ^ _13293;
  wire _35327 = _518 ^ _1359;
  wire _35328 = _35327 ^ _34518;
  wire _35329 = _35326 ^ _35328;
  wire _35330 = _34519 ^ _15396;
  wire _35331 = _34523 ^ _13311;
  wire _35332 = _35330 ^ _35331;
  wire _35333 = _10021 ^ _537;
  wire _35334 = _35333 ^ _12225;
  wire _35335 = _35332 ^ _35334;
  wire _35336 = _35329 ^ _35335;
  wire _35337 = _35324 ^ _35336;
  wire _35338 = _35309 ^ _35337;
  wire _35339 = _35277 ^ _35338;
  wire _35340 = _35216 ^ _35339;
  wire _35341 = _5175 ^ _2172;
  wire _35342 = _21236 ^ _35341;
  wire _35343 = uncoded_block[1137] ^ uncoded_block[1140];
  wire _35344 = _6501 ^ _35343;
  wire _35345 = _24439 ^ _4465;
  wire _35346 = _35344 ^ _35345;
  wire _35347 = _35342 ^ _35346;
  wire _35348 = _33318 ^ _5191;
  wire _35349 = _22627 ^ _7151;
  wire _35350 = _35349 ^ _26685;
  wire _35351 = _35348 ^ _35350;
  wire _35352 = _35347 ^ _35351;
  wire _35353 = _5872 ^ _6519;
  wire _35354 = uncoded_block[1183] ^ uncoded_block[1186];
  wire _35355 = _590 ^ _35354;
  wire _35356 = _35353 ^ _35355;
  wire _35357 = _12808 ^ _19815;
  wire _35358 = _35357 ^ _16906;
  wire _35359 = _35356 ^ _35358;
  wire _35360 = uncoded_block[1213] ^ uncoded_block[1218];
  wire _35361 = _26694 ^ _35360;
  wire _35362 = _26693 ^ _35361;
  wire _35363 = _5215 ^ _8958;
  wire _35364 = uncoded_block[1228] ^ uncoded_block[1232];
  wire _35365 = _35364 ^ _5219;
  wire _35366 = _35363 ^ _35365;
  wire _35367 = _35362 ^ _35366;
  wire _35368 = _35359 ^ _35367;
  wire _35369 = _35352 ^ _35368;
  wire _35370 = _10067 ^ _18860;
  wire _35371 = _1449 ^ _3779;
  wire _35372 = _35370 ^ _35371;
  wire _35373 = _32082 ^ _5234;
  wire _35374 = _6550 ^ _34567;
  wire _35375 = _35373 ^ _35374;
  wire _35376 = _35372 ^ _35375;
  wire _35377 = _16419 ^ _7183;
  wire _35378 = _35377 ^ _33346;
  wire _35379 = _13380 ^ _9545;
  wire _35380 = uncoded_block[1296] ^ uncoded_block[1300];
  wire _35381 = _7193 ^ _35380;
  wire _35382 = _35379 ^ _35381;
  wire _35383 = _35378 ^ _35382;
  wire _35384 = _35376 ^ _35383;
  wire _35385 = _20812 ^ _8991;
  wire _35386 = _17435 ^ _14430;
  wire _35387 = _35385 ^ _35386;
  wire _35388 = _21748 ^ _21293;
  wire _35389 = uncoded_block[1324] ^ uncoded_block[1333];
  wire _35390 = _3029 ^ _35389;
  wire _35391 = _35388 ^ _35390;
  wire _35392 = _35387 ^ _35391;
  wire _35393 = _5932 ^ _12292;
  wire _35394 = _35393 ^ _23143;
  wire _35395 = _3041 ^ _16942;
  wire _35396 = _5273 ^ _3045;
  wire _35397 = _35395 ^ _35396;
  wire _35398 = _35394 ^ _35397;
  wire _35399 = _35392 ^ _35398;
  wire _35400 = _35384 ^ _35399;
  wire _35401 = _35369 ^ _35400;
  wire _35402 = uncoded_block[1362] ^ uncoded_block[1366];
  wire _35403 = _35402 ^ _1509;
  wire _35404 = _22229 ^ _16451;
  wire _35405 = _35403 ^ _35404;
  wire _35406 = _3061 ^ _3838;
  wire _35407 = _2293 ^ _21774;
  wire _35408 = _35406 ^ _35407;
  wire _35409 = _35405 ^ _35408;
  wire _35410 = _13939 ^ _1519;
  wire _35411 = _35410 ^ _5958;
  wire _35412 = _34601 ^ _24059;
  wire _35413 = _35411 ^ _35412;
  wire _35414 = _35409 ^ _35413;
  wire _35415 = _5299 ^ _2313;
  wire _35416 = uncoded_block[1438] ^ uncoded_block[1442];
  wire _35417 = _35416 ^ _716;
  wire _35418 = _35415 ^ _35417;
  wire _35419 = _719 ^ _34609;
  wire _35420 = _21790 ^ _35419;
  wire _35421 = _35418 ^ _35420;
  wire _35422 = _3089 ^ _3870;
  wire _35423 = uncoded_block[1468] ^ uncoded_block[1473];
  wire _35424 = _24070 ^ _35423;
  wire _35425 = _35422 ^ _35424;
  wire _35426 = _5316 ^ _1558;
  wire _35427 = uncoded_block[1487] ^ uncoded_block[1493];
  wire _35428 = _5320 ^ _35427;
  wire _35429 = _35426 ^ _35428;
  wire _35430 = _35425 ^ _35429;
  wire _35431 = _35421 ^ _35430;
  wire _35432 = _35414 ^ _35431;
  wire _35433 = _1572 ^ _750;
  wire _35434 = _9047 ^ _35433;
  wire _35435 = _35434 ^ _34625;
  wire _35436 = uncoded_block[1533] ^ uncoded_block[1541];
  wire _35437 = _35436 ^ _4634;
  wire _35438 = _34627 ^ _35437;
  wire _35439 = uncoded_block[1546] ^ uncoded_block[1548];
  wire _35440 = _35439 ^ _13472;
  wire _35441 = _15020 ^ _3914;
  wire _35442 = _35440 ^ _35441;
  wire _35443 = _35438 ^ _35442;
  wire _35444 = _35435 ^ _35443;
  wire _35445 = _2380 ^ _18952;
  wire _35446 = _34637 ^ _35445;
  wire _35447 = _4653 ^ _24565;
  wire _35448 = _33417 ^ _35447;
  wire _35449 = _35446 ^ _35448;
  wire _35450 = uncoded_block[1598] ^ uncoded_block[1602];
  wire _35451 = _35450 ^ _8502;
  wire _35452 = _1625 ^ _3154;
  wire _35453 = _35451 ^ _35452;
  wire _35454 = _12940 ^ _9094;
  wire _35455 = _35454 ^ _13495;
  wire _35456 = _35453 ^ _35455;
  wire _35457 = _35449 ^ _35456;
  wire _35458 = _35444 ^ _35457;
  wire _35459 = _35432 ^ _35458;
  wire _35460 = _35401 ^ _35459;
  wire _35461 = _14525 ^ _2404;
  wire _35462 = _6049 ^ _3948;
  wire _35463 = _35461 ^ _35462;
  wire _35464 = _27651 ^ _17529;
  wire _35465 = _12957 ^ _823;
  wire _35466 = _35464 ^ _35465;
  wire _35467 = _35463 ^ _35466;
  wire _35468 = _19466 ^ _2422;
  wire _35469 = _6059 ^ _5401;
  wire _35470 = _35468 ^ _35469;
  wire _35471 = uncoded_block[1688] ^ uncoded_block[1692];
  wire _35472 = _19475 ^ _35471;
  wire _35473 = _34658 ^ _35472;
  wire _35474 = _35470 ^ _35473;
  wire _35475 = _35467 ^ _35474;
  wire _35476 = _840 ^ _3973;
  wire _35477 = uncoded_block[1701] ^ uncoded_block[1705];
  wire _35478 = _35477 ^ _9126;
  wire _35479 = _35476 ^ _35478;
  wire _35480 = _855 ^ uncoded_block[1719];
  wire _35481 = _35479 ^ _35480;
  wire _35482 = _35475 ^ _35481;
  wire _35483 = _35460 ^ _35482;
  wire _35484 = _35340 ^ _35483;
  wire _35485 = _19959 ^ _1686;
  wire _35486 = _3998 ^ _30036;
  wire _35487 = _35485 ^ _35486;
  wire _35488 = _7353 ^ _24150;
  wire _35489 = _11 ^ _15080;
  wire _35490 = _35488 ^ _35489;
  wire _35491 = _35487 ^ _35490;
  wire _35492 = _8549 ^ _882;
  wire _35493 = _4009 ^ _1699;
  wire _35494 = _35492 ^ _35493;
  wire _35495 = _886 ^ _16572;
  wire _35496 = _20465 ^ _2474;
  wire _35497 = _35495 ^ _35496;
  wire _35498 = _35494 ^ _35497;
  wire _35499 = _35491 ^ _35498;
  wire _35500 = _12435 ^ _11357;
  wire _35501 = _35500 ^ _17576;
  wire _35502 = _6750 ^ _11364;
  wire _35503 = _14061 ^ _35502;
  wire _35504 = _35501 ^ _35503;
  wire _35505 = _4738 ^ _7374;
  wire _35506 = _14068 ^ _11909;
  wire _35507 = _35505 ^ _35506;
  wire _35508 = _33899 ^ _13011;
  wire _35509 = _35508 ^ _4035;
  wire _35510 = _35507 ^ _35509;
  wire _35511 = _35504 ^ _35510;
  wire _35512 = _35499 ^ _35511;
  wire _35513 = _2497 ^ _2501;
  wire _35514 = _2502 ^ _923;
  wire _35515 = _35513 ^ _35514;
  wire _35516 = _20963 ^ _64;
  wire _35517 = _35516 ^ _32234;
  wire _35518 = _35515 ^ _35517;
  wire _35519 = _14082 ^ _32236;
  wire _35520 = _10834 ^ _33069;
  wire _35521 = _35519 ^ _35520;
  wire _35522 = uncoded_block[171] ^ uncoded_block[176];
  wire _35523 = _35522 ^ _18110;
  wire _35524 = _18578 ^ _35523;
  wire _35525 = _35521 ^ _35524;
  wire _35526 = _35518 ^ _35525;
  wire _35527 = _17106 ^ _945;
  wire _35528 = _35527 ^ _20006;
  wire _35529 = _3284 ^ _10849;
  wire _35530 = _12479 ^ _2540;
  wire _35531 = _35529 ^ _35530;
  wire _35532 = _35528 ^ _35531;
  wire _35533 = _5492 ^ _5497;
  wire _35534 = _6171 ^ _15144;
  wire _35535 = _35533 ^ _35534;
  wire _35536 = _16129 ^ _13053;
  wire _35537 = _14117 ^ _8041;
  wire _35538 = _35536 ^ _35537;
  wire _35539 = _35535 ^ _35538;
  wire _35540 = _35532 ^ _35539;
  wire _35541 = _35526 ^ _35540;
  wire _35542 = _35512 ^ _35541;
  wire _35543 = _28808 ^ _30549;
  wire _35544 = uncoded_block[281] ^ uncoded_block[286];
  wire _35545 = _35544 ^ _5522;
  wire _35546 = _3328 ^ _4820;
  wire _35547 = _35545 ^ _35546;
  wire _35548 = _35543 ^ _35547;
  wire _35549 = _34343 ^ _3337;
  wire _35550 = _20535 ^ _35549;
  wire _35551 = _11441 ^ _152;
  wire _35552 = _15169 ^ _35551;
  wire _35553 = _35550 ^ _35552;
  wire _35554 = _35548 ^ _35553;
  wire _35555 = _11444 ^ _9235;
  wire _35556 = _3352 ^ _6857;
  wire _35557 = _35555 ^ _35556;
  wire _35558 = uncoded_block[347] ^ uncoded_block[352];
  wire _35559 = _35558 ^ _3361;
  wire _35560 = _21026 ^ _35559;
  wire _35561 = _35557 ^ _35560;
  wire _35562 = _1029 ^ _2608;
  wire _35563 = uncoded_block[376] ^ uncoded_block[380];
  wire _35564 = _35563 ^ _1038;
  wire _35565 = _35562 ^ _35564;
  wire _35566 = uncoded_block[385] ^ uncoded_block[390];
  wire _35567 = _35566 ^ _3383;
  wire _35568 = _35567 ^ _6882;
  wire _35569 = _35565 ^ _35568;
  wire _35570 = _35561 ^ _35569;
  wire _35571 = _35554 ^ _35570;
  wire _35572 = _3389 ^ _190;
  wire _35573 = uncoded_block[412] ^ uncoded_block[422];
  wire _35574 = _8091 ^ _35573;
  wire _35575 = _35572 ^ _35574;
  wire _35576 = uncoded_block[426] ^ uncoded_block[431];
  wire _35577 = _1060 ^ _35576;
  wire _35578 = _28103 ^ _21974;
  wire _35579 = _35577 ^ _35578;
  wire _35580 = _35575 ^ _35579;
  wire _35581 = _7498 ^ _3411;
  wire _35582 = uncoded_block[451] ^ uncoded_block[456];
  wire _35583 = uncoded_block[457] ^ uncoded_block[462];
  wire _35584 = _35582 ^ _35583;
  wire _35585 = _35581 ^ _35584;
  wire _35586 = _1874 ^ _21523;
  wire _35587 = uncoded_block[475] ^ uncoded_block[479];
  wire _35588 = _1083 ^ _35587;
  wire _35589 = _35586 ^ _35588;
  wire _35590 = _35585 ^ _35589;
  wire _35591 = _35580 ^ _35590;
  wire _35592 = uncoded_block[490] ^ uncoded_block[494];
  wire _35593 = _4194 ^ _35592;
  wire _35594 = _19627 ^ _35593;
  wire _35595 = uncoded_block[507] ^ uncoded_block[514];
  wire _35596 = _2668 ^ _35595;
  wire _35597 = _19635 ^ _35596;
  wire _35598 = _35594 ^ _35597;
  wire _35599 = _28503 ^ _1108;
  wire _35600 = _20099 ^ _4925;
  wire _35601 = _35599 ^ _35600;
  wire _35602 = uncoded_block[532] ^ uncoded_block[536];
  wire _35603 = _35602 ^ _4217;
  wire _35604 = uncoded_block[545] ^ uncoded_block[553];
  wire _35605 = _8132 ^ _35604;
  wire _35606 = _35603 ^ _35605;
  wire _35607 = _35601 ^ _35606;
  wire _35608 = _35598 ^ _35607;
  wire _35609 = _35591 ^ _35608;
  wire _35610 = _35571 ^ _35609;
  wire _35611 = _35542 ^ _35610;
  wire _35612 = _4937 ^ _258;
  wire _35613 = _4223 ^ _3472;
  wire _35614 = _35612 ^ _35613;
  wire _35615 = _28136 ^ _15747;
  wire _35616 = _35615 ^ _21562;
  wire _35617 = _35614 ^ _35616;
  wire _35618 = _2700 ^ _17228;
  wire _35619 = _16229 ^ _35618;
  wire _35620 = _11535 ^ _17232;
  wire _35621 = _7564 ^ _4960;
  wire _35622 = _35620 ^ _35621;
  wire _35623 = _35619 ^ _35622;
  wire _35624 = _35617 ^ _35623;
  wire _35625 = _12618 ^ _1154;
  wire _35626 = _35625 ^ _28149;
  wire _35627 = _31506 ^ _4255;
  wire _35628 = _35627 ^ _17737;
  wire _35629 = _35626 ^ _35628;
  wire _35630 = uncoded_block[649] ^ uncoded_block[653];
  wire _35631 = _10425 ^ _35630;
  wire _35632 = _8755 ^ _15270;
  wire _35633 = _35631 ^ _35632;
  wire _35634 = _13726 ^ _1177;
  wire _35635 = uncoded_block[680] ^ uncoded_block[685];
  wire _35636 = _6349 ^ _35635;
  wire _35637 = _35634 ^ _35636;
  wire _35638 = _35633 ^ _35637;
  wire _35639 = _35629 ^ _35638;
  wire _35640 = _35624 ^ _35639;
  wire _35641 = _322 ^ _29756;
  wire _35642 = _19195 ^ _4990;
  wire _35643 = _35641 ^ _35642;
  wire _35644 = _14255 ^ _22499;
  wire _35645 = _17266 ^ _341;
  wire _35646 = _35644 ^ _35645;
  wire _35647 = _35643 ^ _35646;
  wire _35648 = _1989 ^ _29766;
  wire _35649 = _14264 ^ _5013;
  wire _35650 = _32781 ^ _35649;
  wire _35651 = _35648 ^ _35650;
  wire _35652 = _35647 ^ _35651;
  wire _35653 = _2777 ^ _7013;
  wire _35654 = uncoded_block[755] ^ uncoded_block[764];
  wire _35655 = _35654 ^ _367;
  wire _35656 = _35653 ^ _35655;
  wire _35657 = _27017 ^ _16786;
  wire _35658 = _35657 ^ _27835;
  wire _35659 = _35656 ^ _35658;
  wire _35660 = _2801 ^ _22071;
  wire _35661 = _28190 ^ _35660;
  wire _35662 = _35661 ^ _25246;
  wire _35663 = _35659 ^ _35662;
  wire _35664 = _35652 ^ _35663;
  wire _35665 = _35640 ^ _35664;
  wire _35666 = uncoded_block[824] ^ uncoded_block[830];
  wire _35667 = _14290 ^ _35666;
  wire _35668 = uncoded_block[836] ^ uncoded_block[840];
  wire _35669 = _35668 ^ _5058;
  wire _35670 = _35667 ^ _35669;
  wire _35671 = _5064 ^ _5742;
  wire _35672 = _5061 ^ _35671;
  wire _35673 = _35670 ^ _35672;
  wire _35674 = _17803 ^ _5071;
  wire _35675 = _2828 ^ _2830;
  wire _35676 = _35674 ^ _35675;
  wire _35677 = _18304 ^ _8820;
  wire _35678 = uncoded_block[886] ^ uncoded_block[889];
  wire _35679 = _35678 ^ _2061;
  wire _35680 = _35677 ^ _35679;
  wire _35681 = _35676 ^ _35680;
  wire _35682 = _35673 ^ _35681;
  wire _35683 = _12706 ^ _1282;
  wire _35684 = _2070 ^ _7665;
  wire _35685 = _3628 ^ _16315;
  wire _35686 = _35684 ^ _35685;
  wire _35687 = _35683 ^ _35686;
  wire _35688 = uncoded_block[935] ^ uncoded_block[938];
  wire _35689 = _1296 ^ _35688;
  wire _35690 = _35689 ^ _6440;
  wire _35691 = _2865 ^ _27476;
  wire _35692 = uncoded_block[955] ^ uncoded_block[961];
  wire _35693 = _5779 ^ _35692;
  wire _35694 = _35691 ^ _35693;
  wire _35695 = _35690 ^ _35694;
  wire _35696 = _35687 ^ _35695;
  wire _35697 = _35682 ^ _35696;
  wire _35698 = _11649 ^ _32425;
  wire _35699 = _23931 ^ _35698;
  wire _35700 = _471 ^ _29832;
  wire _35701 = _2102 ^ _480;
  wire _35702 = _35700 ^ _35701;
  wire _35703 = _35699 ^ _35702;
  wire _35704 = uncoded_block[999] ^ uncoded_block[1002];
  wire _35705 = _35704 ^ _11104;
  wire _35706 = _1331 ^ _5134;
  wire _35707 = _35705 ^ _35706;
  wire _35708 = uncoded_block[1018] ^ uncoded_block[1021];
  wire _35709 = _35708 ^ _5137;
  wire _35710 = uncoded_block[1026] ^ uncoded_block[1032];
  wire _35711 = _8301 ^ _35710;
  wire _35712 = _35709 ^ _35711;
  wire _35713 = _35707 ^ _35712;
  wire _35714 = _35703 ^ _35713;
  wire _35715 = _19768 ^ _512;
  wire _35716 = _22132 ^ _2134;
  wire _35717 = _35715 ^ _35716;
  wire _35718 = _13295 ^ _519;
  wire _35719 = uncoded_block[1059] ^ uncoded_block[1063];
  wire _35720 = _35719 ^ _8888;
  wire _35721 = _35718 ^ _35720;
  wire _35722 = _35717 ^ _35721;
  wire _35723 = uncoded_block[1067] ^ uncoded_block[1073];
  wire _35724 = _35723 ^ _5832;
  wire _35725 = _12219 ^ _30740;
  wire _35726 = _35724 ^ _35725;
  wire _35727 = _16880 ^ _3711;
  wire _35728 = _34527 ^ _35727;
  wire _35729 = _35726 ^ _35728;
  wire _35730 = _35722 ^ _35729;
  wire _35731 = _35714 ^ _35730;
  wire _35732 = _35697 ^ _35731;
  wire _35733 = _35665 ^ _35732;
  wire _35734 = _35611 ^ _35733;
  wire _35735 = _4451 ^ _25323;
  wire _35736 = _35735 ^ _12790;
  wire _35737 = _33312 ^ _9494;
  wire _35738 = _5181 ^ _20269;
  wire _35739 = _35737 ^ _35738;
  wire _35740 = _35736 ^ _35739;
  wire _35741 = _32468 ^ _2185;
  wire _35742 = _35741 ^ _3729;
  wire _35743 = _578 ^ _2964;
  wire _35744 = _15907 ^ _27537;
  wire _35745 = _35743 ^ _35744;
  wire _35746 = _35742 ^ _35745;
  wire _35747 = _35740 ^ _35746;
  wire _35748 = _27902 ^ _31637;
  wire _35749 = uncoded_block[1188] ^ uncoded_block[1192];
  wire _35750 = _4486 ^ _35749;
  wire _35751 = _35748 ^ _35750;
  wire _35752 = _8367 ^ _11170;
  wire _35753 = _35751 ^ _35752;
  wire _35754 = _18395 ^ _11726;
  wire _35755 = _2218 ^ _35754;
  wire _35756 = _608 ^ _8958;
  wire _35757 = _35756 ^ _18405;
  wire _35758 = _35755 ^ _35757;
  wire _35759 = _35753 ^ _35758;
  wire _35760 = _35747 ^ _35759;
  wire _35761 = _3772 ^ _6536;
  wire _35762 = _4509 ^ _1449;
  wire _35763 = _35761 ^ _35762;
  wire _35764 = _4511 ^ _5231;
  wire _35765 = _24471 ^ _3003;
  wire _35766 = _35764 ^ _35765;
  wire _35767 = _35763 ^ _35766;
  wire _35768 = _6554 ^ _7792;
  wire _35769 = _11744 ^ _35768;
  wire _35770 = _3793 ^ _9541;
  wire _35771 = _20808 ^ _33771;
  wire _35772 = _35770 ^ _35771;
  wire _35773 = _35769 ^ _35772;
  wire _35774 = _35767 ^ _35773;
  wire _35775 = _18870 ^ _2259;
  wire _35776 = _17435 ^ _9552;
  wire _35777 = _35775 ^ _35776;
  wire _35778 = _1494 ^ _4550;
  wire _35779 = _24492 ^ _35778;
  wire _35780 = _35777 ^ _35779;
  wire _35781 = _3034 ^ _9563;
  wire _35782 = _2277 ^ _11218;
  wire _35783 = _35781 ^ _35782;
  wire _35784 = _33363 ^ _10097;
  wire _35785 = _5275 ^ _15962;
  wire _35786 = _35784 ^ _35785;
  wire _35787 = _35783 ^ _35786;
  wire _35788 = _35780 ^ _35787;
  wire _35789 = _35774 ^ _35788;
  wire _35790 = _35760 ^ _35789;
  wire _35791 = _22224 ^ _15966;
  wire _35792 = uncoded_block[1384] ^ uncoded_block[1392];
  wire _35793 = _3834 ^ _35792;
  wire _35794 = _35791 ^ _35793;
  wire _35795 = _694 ^ _10676;
  wire _35796 = _35795 ^ _13418;
  wire _35797 = _35794 ^ _35796;
  wire _35798 = uncoded_block[1405] ^ uncoded_block[1417];
  wire _35799 = _35798 ^ _3072;
  wire _35800 = _32948 ^ _2313;
  wire _35801 = _35799 ^ _35800;
  wire _35802 = _1540 ^ _4590;
  wire _35803 = _35802 ^ _35025;
  wire _35804 = _35801 ^ _35803;
  wire _35805 = _35797 ^ _35804;
  wire _35806 = _26309 ^ _18465;
  wire _35807 = _35806 ^ _29102;
  wire _35808 = _8455 ^ _1550;
  wire _35809 = _1555 ^ _4607;
  wire _35810 = _35808 ^ _35809;
  wire _35811 = _35807 ^ _35810;
  wire _35812 = uncoded_block[1495] ^ uncoded_block[1501];
  wire _35813 = _9614 ^ _35812;
  wire _35814 = _26777 ^ _35813;
  wire _35815 = uncoded_block[1503] ^ uncoded_block[1510];
  wire _35816 = _35815 ^ _7875;
  wire _35817 = uncoded_block[1516] ^ uncoded_block[1519];
  wire _35818 = _9055 ^ _35817;
  wire _35819 = _35816 ^ _35818;
  wire _35820 = _35814 ^ _35819;
  wire _35821 = _35811 ^ _35820;
  wire _35822 = _35805 ^ _35821;
  wire _35823 = _26784 ^ _9631;
  wire _35824 = _10717 ^ _35823;
  wire _35825 = _1589 ^ _35439;
  wire _35826 = _15010 ^ _35825;
  wire _35827 = _35824 ^ _35826;
  wire _35828 = uncoded_block[1555] ^ uncoded_block[1561];
  wire _35829 = _15020 ^ _35828;
  wire _35830 = _11283 ^ _4645;
  wire _35831 = _35829 ^ _35830;
  wire _35832 = _1608 ^ _13479;
  wire _35833 = _11838 ^ _16515;
  wire _35834 = _35832 ^ _35833;
  wire _35835 = _35831 ^ _35834;
  wire _35836 = _35827 ^ _35835;
  wire _35837 = uncoded_block[1595] ^ uncoded_block[1599];
  wire _35838 = _11292 ^ _35837;
  wire _35839 = _6039 ^ _14000;
  wire _35840 = _35838 ^ _35839;
  wire _35841 = _24115 ^ _22292;
  wire _35842 = _14525 ^ _13496;
  wire _35843 = _35841 ^ _35842;
  wire _35844 = _35840 ^ _35843;
  wire _35845 = _2405 ^ _6689;
  wire _35846 = _17527 ^ _1649;
  wire _35847 = _35845 ^ _35846;
  wire _35848 = _1654 ^ _4687;
  wire _35849 = _15049 ^ _35848;
  wire _35850 = _35847 ^ _35849;
  wire _35851 = _35844 ^ _35850;
  wire _35852 = _35836 ^ _35851;
  wire _35853 = _35822 ^ _35852;
  wire _35854 = _35790 ^ _35853;
  wire _35855 = uncoded_block[1678] ^ uncoded_block[1682];
  wire _35856 = _6059 ^ _35855;
  wire _35857 = _35856 ^ _25922;
  wire _35858 = _14025 ^ _2435;
  wire _35859 = _841 ^ _35858;
  wire _35860 = _35857 ^ _35859;
  wire _35861 = _3200 ^ uncoded_block[1715];
  wire _35862 = _35860 ^ _35861;
  wire _35863 = _35854 ^ _35862;
  wire _35864 = _35734 ^ _35863;
  wire _35865 = uncoded_block[7] ^ uncoded_block[13];
  wire _35866 = _21407 ^ _35865;
  wire _35867 = _871 ^ _10791;
  wire _35868 = _35866 ^ _35867;
  wire _35869 = _4001 ^ _9143;
  wire _35870 = _35869 ^ _17;
  wire _35871 = _35868 ^ _35870;
  wire _35872 = _24610 ^ _28005;
  wire _35873 = _10238 ^ _6742;
  wire _35874 = _16577 ^ _897;
  wire _35875 = _35873 ^ _35874;
  wire _35876 = _35872 ^ _35875;
  wire _35877 = _35871 ^ _35876;
  wire _35878 = _6109 ^ _4735;
  wire _35879 = _35878 ^ _13559;
  wire _35880 = uncoded_block[98] ^ uncoded_block[103];
  wire _35881 = _6758 ^ _35880;
  wire _35882 = _17580 ^ _35881;
  wire _35883 = _35879 ^ _35882;
  wire _35884 = uncoded_block[119] ^ uncoded_block[127];
  wire _35885 = _13014 ^ _35884;
  wire _35886 = _31383 ^ _35885;
  wire _35887 = _9180 ^ _6138;
  wire _35888 = _6775 ^ _35887;
  wire _35889 = _35886 ^ _35888;
  wire _35890 = _35883 ^ _35889;
  wire _35891 = _35877 ^ _35890;
  wire _35892 = _9182 ^ _1744;
  wire _35893 = _1745 ^ _5469;
  wire _35894 = _35892 ^ _35893;
  wire _35895 = _3271 ^ _24182;
  wire _35896 = _12463 ^ _1751;
  wire _35897 = _35895 ^ _35896;
  wire _35898 = _35894 ^ _35897;
  wire _35899 = _7399 ^ _1756;
  wire _35900 = _940 ^ _13034;
  wire _35901 = _35899 ^ _35900;
  wire _35902 = _2528 ^ _4062;
  wire _35903 = _7409 ^ _4776;
  wire _35904 = _35902 ^ _35903;
  wire _35905 = _35901 ^ _35904;
  wire _35906 = _35898 ^ _35905;
  wire _35907 = _6800 ^ _8018;
  wire _35908 = uncoded_block[203] ^ uncoded_block[205];
  wire _35909 = uncoded_block[208] ^ uncoded_block[214];
  wire _35910 = _35908 ^ _35909;
  wire _35911 = _35907 ^ _35910;
  wire _35912 = uncoded_block[221] ^ uncoded_block[225];
  wire _35913 = _6811 ^ _35912;
  wire _35914 = _4791 ^ _8029;
  wire _35915 = _35913 ^ _35914;
  wire _35916 = _35911 ^ _35915;
  wire _35917 = _6824 ^ _10860;
  wire _35918 = _16129 ^ _14116;
  wire _35919 = _35917 ^ _35918;
  wire _35920 = _6185 ^ _6188;
  wire _35921 = _19564 ^ _35920;
  wire _35922 = _35919 ^ _35921;
  wire _35923 = _35916 ^ _35922;
  wire _35924 = _35906 ^ _35923;
  wire _35925 = _35891 ^ _35924;
  wire _35926 = _33099 ^ _10872;
  wire _35927 = _35926 ^ _25563;
  wire _35928 = _24212 ^ _9772;
  wire _35929 = uncoded_block[292] ^ uncoded_block[297];
  wire _35930 = _10876 ^ _35929;
  wire _35931 = _35928 ^ _35930;
  wire _35932 = _35927 ^ _35931;
  wire _35933 = uncoded_block[301] ^ uncoded_block[304];
  wire _35934 = _8636 ^ _35933;
  wire _35935 = _28067 ^ _23764;
  wire _35936 = _35934 ^ _35935;
  wire _35937 = _15677 ^ _9240;
  wire _35938 = _15676 ^ _35937;
  wire _35939 = _35936 ^ _35938;
  wire _35940 = _35932 ^ _35939;
  wire _35941 = _5536 ^ _2593;
  wire _35942 = _35941 ^ _9788;
  wire _35943 = _19090 ^ _25582;
  wire _35944 = _35942 ^ _35943;
  wire _35945 = uncoded_block[360] ^ uncoded_block[365];
  wire _35946 = _35945 ^ _3369;
  wire _35947 = _10334 ^ _8079;
  wire _35948 = _35946 ^ _35947;
  wire _35949 = _4854 ^ _12538;
  wire _35950 = _1842 ^ _3381;
  wire _35951 = _35949 ^ _35950;
  wire _35952 = _35948 ^ _35951;
  wire _35953 = _35944 ^ _35952;
  wire _35954 = _35940 ^ _35953;
  wire _35955 = _2615 ^ _177;
  wire _35956 = uncoded_block[398] ^ uncoded_block[404];
  wire _35957 = _10910 ^ _35956;
  wire _35958 = _35955 ^ _35957;
  wire _35959 = _33971 ^ _191;
  wire _35960 = _3396 ^ _8665;
  wire _35961 = _35959 ^ _35960;
  wire _35962 = _35958 ^ _35961;
  wire _35963 = _9816 ^ _13115;
  wire _35964 = _8673 ^ _35963;
  wire _35965 = _5574 ^ _21049;
  wire _35966 = _206 ^ _9275;
  wire _35967 = _35965 ^ _35966;
  wire _35968 = _35964 ^ _35967;
  wire _35969 = _35962 ^ _35968;
  wire _35970 = _11486 ^ _1070;
  wire _35971 = _1867 ^ _26495;
  wire _35972 = _35970 ^ _35971;
  wire _35973 = _8681 ^ _15715;
  wire _35974 = _4890 ^ _1079;
  wire _35975 = _35973 ^ _35974;
  wire _35976 = _35972 ^ _35975;
  wire _35977 = uncoded_block[473] ^ uncoded_block[478];
  wire _35978 = _1082 ^ _35977;
  wire _35979 = _35978 ^ _12570;
  wire _35980 = _2660 ^ _2665;
  wire _35981 = _5604 ^ _228;
  wire _35982 = _35980 ^ _35981;
  wire _35983 = _35979 ^ _35982;
  wire _35984 = _35976 ^ _35983;
  wire _35985 = _35969 ^ _35984;
  wire _35986 = _35954 ^ _35985;
  wire _35987 = _35925 ^ _35986;
  wire _35988 = _7521 ^ _2671;
  wire _35989 = _5611 ^ _7531;
  wire _35990 = _35988 ^ _35989;
  wire _35991 = _8122 ^ _236;
  wire _35992 = uncoded_block[520] ^ uncoded_block[527];
  wire _35993 = _35992 ^ _20603;
  wire _35994 = _35991 ^ _35993;
  wire _35995 = _35990 ^ _35994;
  wire _35996 = uncoded_block[545] ^ uncoded_block[555];
  wire _35997 = _1908 ^ _35996;
  wire _35998 = _6294 ^ _35997;
  wire _35999 = _31490 ^ _13165;
  wire _36000 = _3462 ^ _35999;
  wire _36001 = _35998 ^ _36000;
  wire _36002 = _35995 ^ _36001;
  wire _36003 = _13698 ^ _28136;
  wire _36004 = _36003 ^ _25190;
  wire _36005 = _19656 ^ _4236;
  wire _36006 = _4952 ^ _9868;
  wire _36007 = _36005 ^ _36006;
  wire _36008 = _36004 ^ _36007;
  wire _36009 = _16233 ^ _4242;
  wire _36010 = _6959 ^ _1946;
  wire _36011 = _36009 ^ _36010;
  wire _36012 = _14224 ^ _4964;
  wire _36013 = _36012 ^ _21103;
  wire _36014 = _36011 ^ _36013;
  wire _36015 = _36008 ^ _36014;
  wire _36016 = _36002 ^ _36015;
  wire _36017 = uncoded_block[644] ^ uncoded_block[647];
  wire _36018 = _6336 ^ _36017;
  wire _36019 = _28527 ^ _36018;
  wire _36020 = _19177 ^ _28908;
  wire _36021 = _304 ^ _3513;
  wire _36022 = _36020 ^ _36021;
  wire _36023 = _36019 ^ _36022;
  wire _36024 = _309 ^ _1174;
  wire _36025 = _7583 ^ _36024;
  wire _36026 = _1971 ^ _3526;
  wire _36027 = _32349 ^ _36026;
  wire _36028 = _36025 ^ _36027;
  wire _36029 = _36023 ^ _36028;
  wire _36030 = _11556 ^ _4987;
  wire _36031 = _22491 ^ _36030;
  wire _36032 = _5685 ^ _336;
  wire _36033 = _28542 ^ _36032;
  wire _36034 = _36031 ^ _36033;
  wire _36035 = _4996 ^ _3536;
  wire _36036 = uncoded_block[715] ^ uncoded_block[721];
  wire _36037 = _36036 ^ _5691;
  wire _36038 = _36035 ^ _36037;
  wire _36039 = _344 ^ _2768;
  wire _36040 = uncoded_block[739] ^ uncoded_block[743];
  wire _36041 = _7605 ^ _36040;
  wire _36042 = _36039 ^ _36041;
  wire _36043 = _36038 ^ _36042;
  wire _36044 = _36034 ^ _36043;
  wire _36045 = _36029 ^ _36044;
  wire _36046 = _36016 ^ _36045;
  wire _36047 = _25229 ^ _22060;
  wire _36048 = _10470 ^ _1218;
  wire _36049 = _27014 ^ _36048;
  wire _36050 = _36047 ^ _36049;
  wire _36051 = _15799 ^ _14278;
  wire _36052 = _2015 ^ _5032;
  wire _36053 = _36051 ^ _36052;
  wire _36054 = _19223 ^ _385;
  wire _36055 = _18753 ^ _36054;
  wire _36056 = _36053 ^ _36055;
  wire _36057 = _36050 ^ _36056;
  wire _36058 = uncoded_block[802] ^ uncoded_block[812];
  wire _36059 = _36058 ^ _5045;
  wire _36060 = _36059 ^ _1243;
  wire _36061 = _14290 ^ _23450;
  wire _36062 = _6401 ^ _17797;
  wire _36063 = _36061 ^ _36062;
  wire _36064 = _36060 ^ _36063;
  wire _36065 = _1254 ^ _11609;
  wire _36066 = _12689 ^ _36065;
  wire _36067 = _14815 ^ _18764;
  wire _36068 = _36066 ^ _36067;
  wire _36069 = _36064 ^ _36068;
  wire _36070 = _36057 ^ _36069;
  wire _36071 = _30258 ^ _34879;
  wire _36072 = _5072 ^ _9953;
  wire _36073 = _36072 ^ _3609;
  wire _36074 = _36071 ^ _36073;
  wire _36075 = _17811 ^ _8250;
  wire _36076 = _25259 ^ _36075;
  wire _36077 = _5089 ^ _22096;
  wire _36078 = _6428 ^ _6430;
  wire _36079 = _36077 ^ _36078;
  wire _36080 = _36076 ^ _36079;
  wire _36081 = _36074 ^ _36080;
  wire _36082 = _2852 ^ _8259;
  wire _36083 = _31141 ^ _7075;
  wire _36084 = _36082 ^ _36083;
  wire _36085 = _12717 ^ _2862;
  wire _36086 = _36085 ^ _6440;
  wire _36087 = _36084 ^ _36086;
  wire _36088 = _9433 ^ _5779;
  wire _36089 = _461 ^ _10528;
  wire _36090 = _36088 ^ _36089;
  wire _36091 = _1310 ^ _2093;
  wire _36092 = _8847 ^ _13272;
  wire _36093 = _36091 ^ _36092;
  wire _36094 = _36090 ^ _36093;
  wire _36095 = _36087 ^ _36094;
  wire _36096 = _36081 ^ _36095;
  wire _36097 = _36070 ^ _36096;
  wire _36098 = _36046 ^ _36097;
  wire _36099 = _35987 ^ _36098;
  wire _36100 = _8856 ^ _1323;
  wire _36101 = _27485 ^ _36100;
  wire _36102 = _10543 ^ _480;
  wire _36103 = _2107 ^ _22585;
  wire _36104 = _36102 ^ _36103;
  wire _36105 = _36101 ^ _36104;
  wire _36106 = _4405 ^ _487;
  wire _36107 = _8296 ^ _2891;
  wire _36108 = _36106 ^ _36107;
  wire _36109 = _16853 ^ _8872;
  wire _36110 = _11666 ^ _499;
  wire _36111 = _36109 ^ _36110;
  wire _36112 = _36108 ^ _36111;
  wire _36113 = _36105 ^ _36112;
  wire _36114 = _2908 ^ _511;
  wire _36115 = _12208 ^ _17855;
  wire _36116 = _36114 ^ _36115;
  wire _36117 = _12762 ^ _8311;
  wire _36118 = _4431 ^ _20247;
  wire _36119 = _36117 ^ _36118;
  wire _36120 = _36116 ^ _36119;
  wire _36121 = _8889 ^ _13851;
  wire _36122 = _2146 ^ _6486;
  wire _36123 = _36121 ^ _36122;
  wire _36124 = _7724 ^ _1373;
  wire _36125 = _1374 ^ _31189;
  wire _36126 = _36124 ^ _36125;
  wire _36127 = _36123 ^ _36126;
  wire _36128 = _36120 ^ _36127;
  wire _36129 = _36113 ^ _36128;
  wire _36130 = _8330 ^ _545;
  wire _36131 = _8914 ^ _4450;
  wire _36132 = _36130 ^ _36131;
  wire _36133 = _4451 ^ _1388;
  wire _36134 = uncoded_block[1121] ^ uncoded_block[1125];
  wire _36135 = _3714 ^ _36134;
  wire _36136 = _36133 ^ _36135;
  wire _36137 = _36132 ^ _36136;
  wire _36138 = _23523 ^ _5856;
  wire _36139 = uncoded_block[1140] ^ uncoded_block[1142];
  wire _36140 = uncoded_block[1143] ^ uncoded_block[1151];
  wire _36141 = _36139 ^ _36140;
  wire _36142 = _36138 ^ _36141;
  wire _36143 = _5190 ^ _2188;
  wire _36144 = _20276 ^ _36143;
  wire _36145 = _36142 ^ _36144;
  wire _36146 = _36137 ^ _36145;
  wire _36147 = _13335 ^ _11160;
  wire _36148 = _584 ^ _4481;
  wire _36149 = _36147 ^ _36148;
  wire _36150 = _10612 ^ _11719;
  wire _36151 = _30764 ^ _36150;
  wire _36152 = _36149 ^ _36151;
  wire _36153 = _3755 ^ _1427;
  wire _36154 = _33748 ^ _36153;
  wire _36155 = uncoded_block[1221] ^ uncoded_block[1230];
  wire _36156 = _4499 ^ _36155;
  wire _36157 = _17905 ^ _36156;
  wire _36158 = _36154 ^ _36157;
  wire _36159 = _36152 ^ _36158;
  wire _36160 = _36146 ^ _36159;
  wire _36161 = _36129 ^ _36160;
  wire _36162 = _1440 ^ _2226;
  wire _36163 = _8962 ^ _4509;
  wire _36164 = _36162 ^ _36163;
  wire _36165 = _621 ^ _5231;
  wire _36166 = _15445 ^ _36165;
  wire _36167 = _36164 ^ _36166;
  wire _36168 = _11739 ^ _624;
  wire _36169 = _3003 ^ _2244;
  wire _36170 = _36168 ^ _36169;
  wire _36171 = _9538 ^ _16419;
  wire _36172 = _36171 ^ _3795;
  wire _36173 = _36170 ^ _36172;
  wire _36174 = _36167 ^ _36173;
  wire _36175 = _6557 ^ _5913;
  wire _36176 = _3801 ^ _22662;
  wire _36177 = _36175 ^ _36176;
  wire _36178 = _1480 ^ _20816;
  wire _36179 = _31246 ^ _36178;
  wire _36180 = _36177 ^ _36179;
  wire _36181 = _23134 ^ _3029;
  wire _36182 = _36181 ^ _5929;
  wire _36183 = _4551 ^ _9563;
  wire _36184 = _4553 ^ _13927;
  wire _36185 = _36183 ^ _36184;
  wire _36186 = _36182 ^ _36185;
  wire _36187 = _36180 ^ _36186;
  wire _36188 = _36174 ^ _36187;
  wire _36189 = _15473 ^ _6587;
  wire _36190 = _10096 ^ _36189;
  wire _36191 = _4559 ^ _5275;
  wire _36192 = _677 ^ _10665;
  wire _36193 = _36191 ^ _36192;
  wire _36194 = _36190 ^ _36193;
  wire _36195 = _6594 ^ _12305;
  wire _36196 = _4564 ^ _12311;
  wire _36197 = _36195 ^ _36196;
  wire _36198 = _5950 ^ _6597;
  wire _36199 = _4569 ^ _5955;
  wire _36200 = _36198 ^ _36199;
  wire _36201 = _36197 ^ _36200;
  wire _36202 = _36194 ^ _36201;
  wire _36203 = _3841 ^ _3847;
  wire _36204 = _13422 ^ _3850;
  wire _36205 = _36203 ^ _36204;
  wire _36206 = _7842 ^ _3074;
  wire _36207 = _36206 ^ _10691;
  wire _36208 = _36205 ^ _36207;
  wire _36209 = _14469 ^ _5305;
  wire _36210 = uncoded_block[1447] ^ uncoded_block[1455];
  wire _36211 = _36210 ^ _3088;
  wire _36212 = _36209 ^ _36211;
  wire _36213 = uncoded_block[1458] ^ uncoded_block[1462];
  wire _36214 = _36213 ^ _8455;
  wire _36215 = _36214 ^ _11256;
  wire _36216 = _36212 ^ _36215;
  wire _36217 = _36208 ^ _36216;
  wire _36218 = _36202 ^ _36217;
  wire _36219 = _36188 ^ _36218;
  wire _36220 = _36161 ^ _36219;
  wire _36221 = _735 ^ _1556;
  wire _36222 = _15994 ^ _5988;
  wire _36223 = _36221 ^ _36222;
  wire _36224 = _5329 ^ _6631;
  wire _36225 = _13451 ^ _36224;
  wire _36226 = _36223 ^ _36225;
  wire _36227 = _15515 ^ _3112;
  wire _36228 = _7865 ^ _36227;
  wire _36229 = _15002 ^ _1575;
  wire _36230 = uncoded_block[1519] ^ uncoded_block[1528];
  wire _36231 = _36230 ^ _6002;
  wire _36232 = _36229 ^ _36231;
  wire _36233 = _36228 ^ _36232;
  wire _36234 = _36226 ^ _36233;
  wire _36235 = _6005 ^ _5347;
  wire _36236 = _3906 ^ _16010;
  wire _36237 = _36235 ^ _36236;
  wire _36238 = uncoded_block[1547] ^ uncoded_block[1554];
  wire _36239 = _7274 ^ _36238;
  wire _36240 = uncoded_block[1557] ^ uncoded_block[1562];
  wire _36241 = _22731 ^ _36240;
  wire _36242 = _36239 ^ _36241;
  wire _36243 = _36237 ^ _36242;
  wire _36244 = _2376 ^ _777;
  wire _36245 = _30870 ^ _4651;
  wire _36246 = _36244 ^ _36245;
  wire _36247 = _788 ^ _12934;
  wire _36248 = _27640 ^ _36247;
  wire _36249 = _36246 ^ _36248;
  wire _36250 = _36243 ^ _36249;
  wire _36251 = _36234 ^ _36250;
  wire _36252 = _15541 ^ _11295;
  wire _36253 = _11847 ^ _798;
  wire _36254 = _36252 ^ _36253;
  wire _36255 = _10742 ^ _6040;
  wire _36256 = uncoded_block[1610] ^ uncoded_block[1617];
  wire _36257 = _36256 ^ _9095;
  wire _36258 = _36255 ^ _36257;
  wire _36259 = _36254 ^ _36258;
  wire _36260 = _7300 ^ _807;
  wire _36261 = _8509 ^ _16529;
  wire _36262 = _36260 ^ _36261;
  wire _36263 = uncoded_block[1640] ^ uncoded_block[1647];
  wire _36264 = _7308 ^ _36263;
  wire _36265 = _36264 ^ _14012;
  wire _36266 = _36262 ^ _36265;
  wire _36267 = _36259 ^ _36266;
  wire _36268 = _17534 ^ _31757;
  wire _36269 = uncoded_block[1672] ^ uncoded_block[1675];
  wire _36270 = _36269 ^ _17538;
  wire _36271 = uncoded_block[1684] ^ uncoded_block[1690];
  wire _36272 = _17040 ^ _36271;
  wire _36273 = _36270 ^ _36272;
  wire _36274 = _36268 ^ _36273;
  wire _36275 = _11874 ^ _24137;
  wire _36276 = _22314 ^ _8536;
  wire _36277 = _36275 ^ _36276;
  wire _36278 = _11879 ^ _30027;
  wire _36279 = _2443 ^ uncoded_block[1720];
  wire _36280 = _36278 ^ _36279;
  wire _36281 = _36277 ^ _36280;
  wire _36282 = _36274 ^ _36281;
  wire _36283 = _36267 ^ _36282;
  wire _36284 = _36251 ^ _36283;
  wire _36285 = _36220 ^ _36284;
  wire _36286 = _36099 ^ _36285;
  wire _36287 = _18539 ^ _6082;
  wire _36288 = _36287 ^ _10789;
  wire _36289 = _7956 ^ _5423;
  wire _36290 = _10226 ^ _3220;
  wire _36291 = _36289 ^ _36290;
  wire _36292 = _36288 ^ _36291;
  wire _36293 = uncoded_block[30] ^ uncoded_block[34];
  wire _36294 = _11344 ^ _36293;
  wire _36295 = uncoded_block[35] ^ uncoded_block[39];
  wire _36296 = _36295 ^ _882;
  wire _36297 = _36294 ^ _36296;
  wire _36298 = _22 ^ _12428;
  wire _36299 = _36298 ^ _29597;
  wire _36300 = _36297 ^ _36299;
  wire _36301 = _36292 ^ _36300;
  wire _36302 = _23698 ^ _35;
  wire _36303 = _36302 ^ _10245;
  wire _36304 = _14060 ^ _28438;
  wire _36305 = _18077 ^ _1718;
  wire _36306 = _36304 ^ _36305;
  wire _36307 = _36303 ^ _36306;
  wire _36308 = _1719 ^ _15101;
  wire _36309 = _17584 ^ _1722;
  wire _36310 = _36308 ^ _36309;
  wire _36311 = _19520 ^ _6763;
  wire _36312 = _915 ^ _12451;
  wire _36313 = _36311 ^ _36312;
  wire _36314 = _36310 ^ _36313;
  wire _36315 = _36307 ^ _36314;
  wire _36316 = _36301 ^ _36315;
  wire _36317 = _4751 ^ _9175;
  wire _36318 = _32634 ^ _9177;
  wire _36319 = _36317 ^ _36318;
  wire _36320 = _2510 ^ _5461;
  wire _36321 = _17097 ^ _15622;
  wire _36322 = _36320 ^ _36321;
  wire _36323 = _36319 ^ _36322;
  wire _36324 = _1745 ^ _7397;
  wire _36325 = _1748 ^ _4049;
  wire _36326 = _36324 ^ _36325;
  wire _36327 = _1749 ^ _7399;
  wire _36328 = _35522 ^ _11933;
  wire _36329 = _36327 ^ _36328;
  wire _36330 = _36326 ^ _36329;
  wire _36331 = _36323 ^ _36330;
  wire _36332 = _944 ^ _4062;
  wire _36333 = _13588 ^ _4776;
  wire _36334 = _36332 ^ _36333;
  wire _36335 = _9745 ^ _6805;
  wire _36336 = _3291 ^ _30963;
  wire _36337 = _36335 ^ _36336;
  wire _36338 = _36334 ^ _36337;
  wire _36339 = _27295 ^ _1772;
  wire _36340 = _36339 ^ _35533;
  wire _36341 = _967 ^ _7423;
  wire _36342 = _10288 ^ _36341;
  wire _36343 = _36340 ^ _36342;
  wire _36344 = _36338 ^ _36343;
  wire _36345 = _36331 ^ _36344;
  wire _36346 = _36316 ^ _36345;
  wire _36347 = _10292 ^ _971;
  wire _36348 = uncoded_block[248] ^ uncoded_block[251];
  wire _36349 = _36348 ^ _4803;
  wire _36350 = _36347 ^ _36349;
  wire _36351 = uncoded_block[258] ^ uncoded_block[262];
  wire _36352 = _3311 ^ _36351;
  wire _36353 = _36352 ^ _6189;
  wire _36354 = _36350 ^ _36353;
  wire _36355 = _14642 ^ _3320;
  wire _36356 = _36355 ^ _15661;
  wire _36357 = _11428 ^ _5522;
  wire _36358 = _17635 ^ _14133;
  wire _36359 = _36357 ^ _36358;
  wire _36360 = _36356 ^ _36359;
  wire _36361 = _36354 ^ _36360;
  wire _36362 = _3337 ^ _15671;
  wire _36363 = _10314 ^ _36362;
  wire _36364 = _3341 ^ _13625;
  wire _36365 = _21947 ^ _1821;
  wire _36366 = _36364 ^ _36365;
  wire _36367 = _36363 ^ _36366;
  wire _36368 = _18621 ^ _11454;
  wire _36369 = _28829 ^ _36368;
  wire _36370 = uncoded_block[356] ^ uncoded_block[364];
  wire _36371 = _11455 ^ _36370;
  wire _36372 = _36371 ^ _26917;
  wire _36373 = _36369 ^ _36372;
  wire _36374 = _36367 ^ _36373;
  wire _36375 = _36361 ^ _36374;
  wire _36376 = _1036 ^ _14671;
  wire _36377 = _30128 ^ _36376;
  wire _36378 = _1841 ^ _11999;
  wire _36379 = _6879 ^ _1847;
  wire _36380 = _36378 ^ _36379;
  wire _36381 = _36377 ^ _36380;
  wire _36382 = _34764 ^ _20565;
  wire _36383 = _8091 ^ _24245;
  wire _36384 = _4164 ^ _24248;
  wire _36385 = _36383 ^ _36384;
  wire _36386 = _36382 ^ _36385;
  wire _36387 = _36381 ^ _36386;
  wire _36388 = _23348 ^ _2641;
  wire _36389 = _3408 ^ _12559;
  wire _36390 = _36388 ^ _36389;
  wire _36391 = _3411 ^ _12562;
  wire _36392 = _2650 ^ _213;
  wire _36393 = _36391 ^ _36392;
  wire _36394 = _36390 ^ _36393;
  wire _36395 = _2654 ^ _1878;
  wire _36396 = _33567 ^ _36395;
  wire _36397 = _6266 ^ _12025;
  wire _36398 = _5592 ^ _4895;
  wire _36399 = _36397 ^ _36398;
  wire _36400 = _36396 ^ _36399;
  wire _36401 = _36394 ^ _36400;
  wire _36402 = _36387 ^ _36401;
  wire _36403 = _36375 ^ _36402;
  wire _36404 = _36346 ^ _36403;
  wire _36405 = _6276 ^ _5603;
  wire _36406 = _35199 ^ _36405;
  wire _36407 = _2667 ^ _6921;
  wire _36408 = _36407 ^ _24268;
  wire _36409 = _36406 ^ _36408;
  wire _36410 = _13676 ^ _18665;
  wire _36411 = _16709 ^ _20602;
  wire _36412 = _36410 ^ _36411;
  wire _36413 = _10385 ^ _9854;
  wire _36414 = _31896 ^ _36413;
  wire _36415 = _36412 ^ _36414;
  wire _36416 = _36409 ^ _36415;
  wire _36417 = _25630 ^ _25182;
  wire _36418 = _4937 ^ _9319;
  wire _36419 = _36417 ^ _36418;
  wire _36420 = _5635 ^ _13165;
  wire _36421 = _13698 ^ _1931;
  wire _36422 = _36420 ^ _36421;
  wire _36423 = _36419 ^ _36422;
  wire _36424 = uncoded_block[579] ^ uncoded_block[586];
  wire _36425 = _36424 ^ _4950;
  wire _36426 = _36425 ^ _26100;
  wire _36427 = _4952 ^ _5646;
  wire _36428 = _36427 ^ _34017;
  wire _36429 = _36426 ^ _36428;
  wire _36430 = _36423 ^ _36429;
  wire _36431 = _36416 ^ _36430;
  wire _36432 = _16734 ^ _6325;
  wire _36433 = _13713 ^ _6328;
  wire _36434 = _36432 ^ _36433;
  wire _36435 = uncoded_block[632] ^ uncoded_block[640];
  wire _36436 = _36435 ^ _8751;
  wire _36437 = _30197 ^ _36436;
  wire _36438 = _36434 ^ _36437;
  wire _36439 = _1957 ^ _1960;
  wire _36440 = _4975 ^ _2738;
  wire _36441 = _36439 ^ _36440;
  wire _36442 = uncoded_block[674] ^ uncoded_block[679];
  wire _36443 = _4265 ^ _36442;
  wire _36444 = uncoded_block[690] ^ uncoded_block[699];
  wire _36445 = _15281 ^ _36444;
  wire _36446 = _36443 ^ _36445;
  wire _36447 = _36441 ^ _36446;
  wire _36448 = _36438 ^ _36447;
  wire _36449 = _6992 ^ _17757;
  wire _36450 = _3535 ^ _10452;
  wire _36451 = _36449 ^ _36450;
  wire _36452 = _8193 ^ _2765;
  wire _36453 = _9905 ^ _1991;
  wire _36454 = _36452 ^ _36453;
  wire _36455 = _36451 ^ _36454;
  wire _36456 = _23870 ^ _11576;
  wire _36457 = _12104 ^ _36456;
  wire _36458 = _2775 ^ _31537;
  wire _36459 = _7013 ^ _3556;
  wire _36460 = _36458 ^ _36459;
  wire _36461 = _36457 ^ _36460;
  wire _36462 = _36455 ^ _36461;
  wire _36463 = _36448 ^ _36462;
  wire _36464 = _36431 ^ _36463;
  wire _36465 = _4299 ^ _2781;
  wire _36466 = uncoded_block[766] ^ uncoded_block[770];
  wire _36467 = _2783 ^ _36466;
  wire _36468 = _36465 ^ _36467;
  wire _36469 = uncoded_block[774] ^ uncoded_block[779];
  wire _36470 = _12114 ^ _36469;
  wire _36471 = _3568 ^ _19218;
  wire _36472 = _36470 ^ _36471;
  wire _36473 = _36468 ^ _36472;
  wire _36474 = _2799 ^ _1233;
  wire _36475 = _5722 ^ _36474;
  wire _36476 = _16790 ^ _389;
  wire _36477 = uncoded_block[809] ^ uncoded_block[813];
  wire _36478 = _16791 ^ _36477;
  wire _36479 = _36476 ^ _36478;
  wire _36480 = _36475 ^ _36479;
  wire _36481 = _36473 ^ _36480;
  wire _36482 = _2808 ^ _28197;
  wire _36483 = _23450 ^ _5052;
  wire _36484 = _36482 ^ _36483;
  wire _36485 = _400 ^ _1253;
  wire _36486 = _36485 ^ _19722;
  wire _36487 = _36484 ^ _36486;
  wire _36488 = _5060 ^ _19725;
  wire _36489 = _14814 ^ _2821;
  wire _36490 = _36488 ^ _36489;
  wire _36491 = _3600 ^ _5069;
  wire _36492 = _12150 ^ _33671;
  wire _36493 = _36491 ^ _36492;
  wire _36494 = _36490 ^ _36493;
  wire _36495 = _36487 ^ _36494;
  wire _36496 = _36481 ^ _36495;
  wire _36497 = uncoded_block[883] ^ uncoded_block[885];
  wire _36498 = _5078 ^ _36497;
  wire _36499 = _36498 ^ _25724;
  wire _36500 = _8254 ^ _3623;
  wire _36501 = _17311 ^ _36500;
  wire _36502 = _36499 ^ _36501;
  wire _36503 = _2071 ^ _16313;
  wire _36504 = _36503 ^ _5765;
  wire _36505 = _446 ^ _5096;
  wire _36506 = _15353 ^ _36505;
  wire _36507 = _36504 ^ _36506;
  wire _36508 = _36502 ^ _36507;
  wire _36509 = _10517 ^ _7080;
  wire _36510 = _2084 ^ _23926;
  wire _36511 = _36509 ^ _36510;
  wire _36512 = _10525 ^ _1308;
  wire _36513 = _4383 ^ _36512;
  wire _36514 = _36511 ^ _36513;
  wire _36515 = uncoded_block[968] ^ uncoded_block[971];
  wire _36516 = _36515 ^ _2877;
  wire _36517 = _9982 ^ _36516;
  wire _36518 = uncoded_block[978] ^ uncoded_block[981];
  wire _36519 = _28233 ^ _36518;
  wire _36520 = _23038 ^ _1317;
  wire _36521 = _36519 ^ _36520;
  wire _36522 = _36517 ^ _36521;
  wire _36523 = _36514 ^ _36522;
  wire _36524 = _36508 ^ _36523;
  wire _36525 = _36496 ^ _36524;
  wire _36526 = _36464 ^ _36525;
  wire _36527 = _36404 ^ _36526;
  wire _36528 = _23938 ^ _13277;
  wire _36529 = _5798 ^ _9449;
  wire _36530 = _36528 ^ _36529;
  wire _36531 = _20730 ^ _4405;
  wire _36532 = uncoded_block[1012] ^ uncoded_block[1017];
  wire _36533 = _487 ^ _36532;
  wire _36534 = _36531 ^ _36533;
  wire _36535 = _36530 ^ _36534;
  wire _36536 = _2121 ^ _4417;
  wire _36537 = _22127 ^ _36536;
  wire _36538 = _11668 ^ _2908;
  wire _36539 = _36538 ^ _25766;
  wire _36540 = _36537 ^ _36539;
  wire _36541 = _36535 ^ _36540;
  wire _36542 = _2130 ^ _2913;
  wire _36543 = uncoded_block[1060] ^ uncoded_block[1066];
  wire _36544 = _2136 ^ _36543;
  wire _36545 = _36542 ^ _36544;
  wire _36546 = _3689 ^ _527;
  wire _36547 = _36546 ^ _24422;
  wire _36548 = _36545 ^ _36547;
  wire _36549 = _5834 ^ _534;
  wire _36550 = _4440 ^ _22610;
  wire _36551 = _36549 ^ _36550;
  wire _36552 = _3704 ^ _5169;
  wire _36553 = _36552 ^ _23074;
  wire _36554 = _36551 ^ _36553;
  wire _36555 = _36548 ^ _36554;
  wire _36556 = _36541 ^ _36555;
  wire _36557 = _14882 ^ _2167;
  wire _36558 = _1389 ^ _12791;
  wire _36559 = _36557 ^ _36558;
  wire _36560 = _13866 ^ _564;
  wire _36561 = uncoded_block[1141] ^ uncoded_block[1146];
  wire _36562 = _4462 ^ _36561;
  wire _36563 = _36560 ^ _36562;
  wire _36564 = _36559 ^ _36563;
  wire _36565 = _2186 ^ _29878;
  wire _36566 = _29877 ^ _36565;
  wire _36567 = uncoded_block[1159] ^ uncoded_block[1163];
  wire _36568 = _36567 ^ _6513;
  wire _36569 = _36568 ^ _16388;
  wire _36570 = _36566 ^ _36569;
  wire _36571 = _36564 ^ _36570;
  wire _36572 = _1411 ^ _590;
  wire _36573 = uncoded_block[1184] ^ uncoded_block[1189];
  wire _36574 = _592 ^ _36573;
  wire _36575 = _36572 ^ _36574;
  wire _36576 = _2971 ^ _24910;
  wire _36577 = uncoded_block[1201] ^ uncoded_block[1206];
  wire _36578 = _7758 ^ _36577;
  wire _36579 = _36576 ^ _36578;
  wire _36580 = _36575 ^ _36579;
  wire _36581 = uncoded_block[1208] ^ uncoded_block[1213];
  wire _36582 = _36581 ^ _605;
  wire _36583 = _606 ^ _34556;
  wire _36584 = _36582 ^ _36583;
  wire _36585 = _3772 ^ _17910;
  wire _36586 = _2227 ^ _36585;
  wire _36587 = _36584 ^ _36586;
  wire _36588 = _36580 ^ _36587;
  wire _36589 = _36571 ^ _36588;
  wire _36590 = _36556 ^ _36589;
  wire _36591 = _27131 ^ _18862;
  wire _36592 = uncoded_block[1266] ^ uncoded_block[1269];
  wire _36593 = _9530 ^ _36592;
  wire _36594 = _23557 ^ _36593;
  wire _36595 = _36591 ^ _36594;
  wire _36596 = _27134 ^ _6558;
  wire _36597 = _7193 ^ _645;
  wire _36598 = _24024 ^ _36597;
  wire _36599 = _36596 ^ _36598;
  wire _36600 = _36595 ^ _36599;
  wire _36601 = _2255 ^ _7802;
  wire _36602 = _11199 ^ _36601;
  wire _36603 = _14430 ^ _4540;
  wire _36604 = uncoded_block[1323] ^ uncoded_block[1329];
  wire _36605 = _9555 ^ _36604;
  wire _36606 = _36603 ^ _36605;
  wire _36607 = _36602 ^ _36606;
  wire _36608 = _1494 ^ _18431;
  wire _36609 = _13399 ^ _5262;
  wire _36610 = _36608 ^ _36609;
  wire _36611 = _17938 ^ _670;
  wire _36612 = _36611 ^ _18437;
  wire _36613 = _36610 ^ _36612;
  wire _36614 = _36607 ^ _36613;
  wire _36615 = _36600 ^ _36614;
  wire _36616 = _23581 ^ _3045;
  wire _36617 = _36616 ^ _36192;
  wire _36618 = _12302 ^ _2289;
  wire _36619 = _5285 ^ _6596;
  wire _36620 = _36618 ^ _36619;
  wire _36621 = _36617 ^ _36620;
  wire _36622 = _4569 ^ _35016;
  wire _36623 = _36198 ^ _36622;
  wire _36624 = _9016 ^ _3847;
  wire _36625 = _36624 ^ _9586;
  wire _36626 = _36623 ^ _36625;
  wire _36627 = _36621 ^ _36626;
  wire _36628 = _10118 ^ _16463;
  wire _36629 = _27938 ^ _36628;
  wire _36630 = _15494 ^ _5299;
  wire _36631 = _2313 ^ _3857;
  wire _36632 = _36630 ^ _36631;
  wire _36633 = _36629 ^ _36632;
  wire _36634 = _2318 ^ _6613;
  wire _36635 = uncoded_block[1450] ^ uncoded_block[1455];
  wire _36636 = _8450 ^ _36635;
  wire _36637 = _36634 ^ _36636;
  wire _36638 = _3089 ^ _3879;
  wire _36639 = _14989 ^ _13446;
  wire _36640 = _36638 ^ _36639;
  wire _36641 = _36637 ^ _36640;
  wire _36642 = _36633 ^ _36641;
  wire _36643 = _36627 ^ _36642;
  wire _36644 = _36615 ^ _36643;
  wire _36645 = _36590 ^ _36644;
  wire _36646 = _1558 ^ _17980;
  wire _36647 = _25426 ^ _1565;
  wire _36648 = _36646 ^ _36647;
  wire _36649 = _6631 ^ _6634;
  wire _36650 = _1571 ^ _4614;
  wire _36651 = _36649 ^ _36650;
  wire _36652 = _36648 ^ _36651;
  wire _36653 = uncoded_block[1511] ^ uncoded_block[1517];
  wire _36654 = _24539 ^ _36653;
  wire _36655 = uncoded_block[1519] ^ uncoded_block[1523];
  wire _36656 = uncoded_block[1528] ^ uncoded_block[1534];
  wire _36657 = _36655 ^ _36656;
  wire _36658 = _36654 ^ _36657;
  wire _36659 = _3909 ^ _4634;
  wire _36660 = _34228 ^ _36659;
  wire _36661 = _36658 ^ _36660;
  wire _36662 = _36652 ^ _36661;
  wire _36663 = _2367 ^ _2370;
  wire _36664 = uncoded_block[1553] ^ uncoded_block[1558];
  wire _36665 = _36664 ^ _7888;
  wire _36666 = _36663 ^ _36665;
  wire _36667 = _11283 ^ _7891;
  wire _36668 = _36667 ^ _29133;
  wire _36669 = _36666 ^ _36668;
  wire _36670 = uncoded_block[1578] ^ uncoded_block[1585];
  wire _36671 = _782 ^ _36670;
  wire _36672 = _36671 ^ _34242;
  wire _36673 = _3146 ^ _11294;
  wire _36674 = _36673 ^ _27645;
  wire _36675 = _36672 ^ _36674;
  wire _36676 = _36669 ^ _36675;
  wire _36677 = _36662 ^ _36676;
  wire _36678 = _3153 ^ _7906;
  wire _36679 = _7908 ^ _12376;
  wire _36680 = _36678 ^ _36679;
  wire _36681 = _16528 ^ _30885;
  wire _36682 = _36680 ^ _36681;
  wire _36683 = _7309 ^ _3169;
  wire _36684 = uncoded_block[1646] ^ uncoded_block[1648];
  wire _36685 = _36684 ^ _7314;
  wire _36686 = _36683 ^ _36685;
  wire _36687 = uncoded_block[1657] ^ uncoded_block[1661];
  wire _36688 = _36687 ^ _3179;
  wire _36689 = _36688 ^ _14537;
  wire _36690 = _36686 ^ _36689;
  wire _36691 = _36682 ^ _36690;
  wire _36692 = _7323 ^ _16541;
  wire _36693 = uncoded_block[1686] ^ uncoded_block[1692];
  wire _36694 = _18982 ^ _36693;
  wire _36695 = _36692 ^ _36694;
  wire _36696 = _3972 ^ _5409;
  wire _36697 = _22314 ^ _2437;
  wire _36698 = _36696 ^ _36697;
  wire _36699 = _36695 ^ _36698;
  wire _36700 = _3980 ^ _2441;
  wire _36701 = _36700 ^ uncoded_block[1720];
  wire _36702 = _36699 ^ _36701;
  wire _36703 = _36691 ^ _36702;
  wire _36704 = _36677 ^ _36703;
  wire _36705 = _36645 ^ _36704;
  wire _36706 = _36527 ^ _36705;
  wire _36707 = uncoded_block[4] ^ uncoded_block[13];
  wire _36708 = _36707 ^ _868;
  wire _36709 = _3211 ^ _36708;
  wire _36710 = _6087 ^ _1690;
  wire _36711 = _4000 ^ _9694;
  wire _36712 = _36710 ^ _36711;
  wire _36713 = _36709 ^ _36712;
  wire _36714 = _11344 ^ _11890;
  wire _36715 = _875 ^ _6095;
  wire _36716 = _36714 ^ _36715;
  wire _36717 = _879 ^ _4723;
  wire _36718 = _36717 ^ _34284;
  wire _36719 = _36716 ^ _36718;
  wire _36720 = _36713 ^ _36719;
  wire _36721 = _25 ^ _6106;
  wire _36722 = _36721 ^ _35500;
  wire _36723 = uncoded_block[71] ^ uncoded_block[78];
  wire _36724 = _7367 ^ _36723;
  wire _36725 = _28438 ^ _14586;
  wire _36726 = _36724 ^ _36725;
  wire _36727 = _36722 ^ _36726;
  wire _36728 = uncoded_block[96] ^ uncoded_block[100];
  wire _36729 = _6115 ^ _36728;
  wire _36730 = _16583 ^ _36729;
  wire _36731 = _4028 ^ _4031;
  wire _36732 = _1722 ^ _915;
  wire _36733 = _36731 ^ _36732;
  wire _36734 = _36730 ^ _36733;
  wire _36735 = _36727 ^ _36734;
  wire _36736 = _36720 ^ _36735;
  wire _36737 = _4750 ^ _10256;
  wire _36738 = _11374 ^ _32634;
  wire _36739 = _36737 ^ _36738;
  wire _36740 = _9180 ^ _18100;
  wire _36741 = _73 ^ _21906;
  wire _36742 = _36740 ^ _36741;
  wire _36743 = _36739 ^ _36742;
  wire _36744 = _6788 ^ _81;
  wire _36745 = _15122 ^ _36744;
  wire _36746 = _19539 ^ _5477;
  wire _36747 = uncoded_block[181] ^ uncoded_block[186];
  wire _36748 = _36747 ^ _18113;
  wire _36749 = _36746 ^ _36748;
  wire _36750 = _36745 ^ _36749;
  wire _36751 = _36743 ^ _36750;
  wire _36752 = uncoded_block[194] ^ uncoded_block[201];
  wire _36753 = _36752 ^ _10278;
  wire _36754 = _1764 ^ _956;
  wire _36755 = _36753 ^ _36754;
  wire _36756 = _4787 ^ _7419;
  wire _36757 = _36756 ^ _27299;
  wire _36758 = _36755 ^ _36757;
  wire _36759 = _33088 ^ _5500;
  wire _36760 = _8032 ^ _13053;
  wire _36761 = _36759 ^ _36760;
  wire _36762 = _9762 ^ _19064;
  wire _36763 = _36761 ^ _36762;
  wire _36764 = _36758 ^ _36763;
  wire _36765 = _36751 ^ _36764;
  wire _36766 = _36736 ^ _36765;
  wire _36767 = _15154 ^ _17134;
  wire _36768 = uncoded_block[277] ^ uncoded_block[282];
  wire _36769 = _36768 ^ _19072;
  wire _36770 = _36767 ^ _36769;
  wire _36771 = _34339 ^ _137;
  wire _36772 = _1810 ^ _143;
  wire _36773 = _36771 ^ _36772;
  wire _36774 = _36770 ^ _36773;
  wire _36775 = _26016 ^ _3340;
  wire _36776 = _15677 ^ _11444;
  wire _36777 = _36775 ^ _36776;
  wire _36778 = _9241 ^ _30120;
  wire _36779 = _36777 ^ _36778;
  wire _36780 = _36774 ^ _36779;
  wire _36781 = _4841 ^ _16161;
  wire _36782 = uncoded_block[351] ^ uncoded_block[354];
  wire _36783 = _36782 ^ _21497;
  wire _36784 = _36781 ^ _36783;
  wire _36785 = _5548 ^ _1838;
  wire _36786 = _36785 ^ _19596;
  wire _36787 = _36784 ^ _36786;
  wire _36788 = _10899 ^ _1841;
  wire _36789 = _17661 ^ _10907;
  wire _36790 = _36788 ^ _36789;
  wire _36791 = _5554 ^ _9806;
  wire _36792 = _36791 ^ _31450;
  wire _36793 = _36790 ^ _36792;
  wire _36794 = _36787 ^ _36793;
  wire _36795 = _36780 ^ _36794;
  wire _36796 = uncoded_block[405] ^ uncoded_block[411];
  wire _36797 = _36796 ^ _1055;
  wire _36798 = _36797 ^ _3398;
  wire _36799 = _1063 ^ _2640;
  wire _36800 = _6890 ^ _36799;
  wire _36801 = _36798 ^ _36800;
  wire _36802 = _3405 ^ _5578;
  wire _36803 = _36802 ^ _25156;
  wire _36804 = _17185 ^ _1871;
  wire _36805 = _13662 ^ _2654;
  wire _36806 = _36804 ^ _36805;
  wire _36807 = _36803 ^ _36806;
  wire _36808 = _36801 ^ _36807;
  wire _36809 = _1878 ^ _3418;
  wire _36810 = _221 ^ _21526;
  wire _36811 = _36809 ^ _36810;
  wire _36812 = _5593 ^ _21528;
  wire _36813 = _7516 ^ _3424;
  wire _36814 = _36812 ^ _36813;
  wire _36815 = _36811 ^ _36814;
  wire _36816 = _7520 ^ _2668;
  wire _36817 = _6922 ^ _4208;
  wire _36818 = _36816 ^ _36817;
  wire _36819 = _13152 ^ _1900;
  wire _36820 = _20603 ^ _16215;
  wire _36821 = _36819 ^ _36820;
  wire _36822 = _36818 ^ _36821;
  wire _36823 = _36815 ^ _36822;
  wire _36824 = _36808 ^ _36823;
  wire _36825 = _36795 ^ _36824;
  wire _36826 = _36766 ^ _36825;
  wire _36827 = _7541 ^ _12592;
  wire _36828 = _247 ^ _1915;
  wire _36829 = _36827 ^ _36828;
  wire _36830 = _1123 ^ _8139;
  wire _36831 = _29726 ^ _4223;
  wire _36832 = _36830 ^ _36831;
  wire _36833 = _36829 ^ _36832;
  wire _36834 = _3472 ^ _11527;
  wire _36835 = _8733 ^ _18222;
  wire _36836 = _36834 ^ _36835;
  wire _36837 = _1938 ^ _2701;
  wire _36838 = _2706 ^ _3487;
  wire _36839 = _36837 ^ _36838;
  wire _36840 = _36836 ^ _36839;
  wire _36841 = _36833 ^ _36840;
  wire _36842 = uncoded_block[606] ^ uncoded_block[612];
  wire _36843 = _8738 ^ _36842;
  wire _36844 = _7564 ^ _7567;
  wire _36845 = _36843 ^ _36844;
  wire _36846 = _29313 ^ _1154;
  wire _36847 = uncoded_block[629] ^ uncoded_block[633];
  wire _36848 = _36847 ^ _5661;
  wire _36849 = _36846 ^ _36848;
  wire _36850 = _36845 ^ _36849;
  wire _36851 = _3505 ^ _6973;
  wire _36852 = _7579 ^ _36851;
  wire _36853 = uncoded_block[652] ^ uncoded_block[658];
  wire _36854 = _36853 ^ _8172;
  wire _36855 = _4262 ^ _10990;
  wire _36856 = _36854 ^ _36855;
  wire _36857 = _36852 ^ _36856;
  wire _36858 = _36850 ^ _36857;
  wire _36859 = _36841 ^ _36858;
  wire _36860 = _8177 ^ _6352;
  wire _36861 = _15276 ^ _36860;
  wire _36862 = _18247 ^ _15281;
  wire _36863 = _36862 ^ _13736;
  wire _36864 = _36861 ^ _36863;
  wire _36865 = _6361 ^ _10448;
  wire _36866 = _28542 ^ _36865;
  wire _36867 = _12097 ^ _16767;
  wire _36868 = _36866 ^ _36867;
  wire _36869 = _36864 ^ _36868;
  wire _36870 = _5693 ^ _2768;
  wire _36871 = _349 ^ _1206;
  wire _36872 = _36870 ^ _36871;
  wire _36873 = uncoded_block[746] ^ uncoded_block[750];
  wire _36874 = _36873 ^ _7013;
  wire _36875 = _22977 ^ _36874;
  wire _36876 = _36872 ^ _36875;
  wire _36877 = _24796 ^ _4301;
  wire _36878 = uncoded_block[772] ^ uncoded_block[780];
  wire _36879 = _11019 ^ _36878;
  wire _36880 = _36877 ^ _36879;
  wire _36881 = _1225 ^ _3574;
  wire _36882 = _20172 ^ _36881;
  wire _36883 = _36880 ^ _36882;
  wire _36884 = _36876 ^ _36883;
  wire _36885 = _36869 ^ _36884;
  wire _36886 = _36859 ^ _36885;
  wire _36887 = _8224 ^ _3577;
  wire _36888 = _36887 ^ _30245;
  wire _36889 = _22525 ^ _15320;
  wire _36890 = _1250 ^ _401;
  wire _36891 = _36889 ^ _36890;
  wire _36892 = _36888 ^ _36891;
  wire _36893 = _9938 ^ _5057;
  wire _36894 = _36893 ^ _32395;
  wire _36895 = _3599 ^ _7643;
  wire _36896 = _6406 ^ _3600;
  wire _36897 = _36895 ^ _36896;
  wire _36898 = _36894 ^ _36897;
  wire _36899 = _36892 ^ _36898;
  wire _36900 = _2047 ^ _9948;
  wire _36901 = _36900 ^ _10500;
  wire _36902 = _6415 ^ _33671;
  wire _36903 = uncoded_block[881] ^ uncoded_block[883];
  wire _36904 = _16304 ^ _36903;
  wire _36905 = _36902 ^ _36904;
  wire _36906 = _36901 ^ _36905;
  wire _36907 = _14827 ^ _5083;
  wire _36908 = _20700 ^ _36907;
  wire _36909 = _2843 ^ _6425;
  wire _36910 = _5086 ^ _36909;
  wire _36911 = _36908 ^ _36910;
  wire _36912 = _36906 ^ _36911;
  wire _36913 = _36899 ^ _36912;
  wire _36914 = _9421 ^ _2071;
  wire _36915 = uncoded_block[917] ^ uncoded_block[927];
  wire _36916 = _3628 ^ _36915;
  wire _36917 = _36914 ^ _36916;
  wire _36918 = _4371 ^ _3637;
  wire _36919 = _15848 ^ _10523;
  wire _36920 = _36918 ^ _36919;
  wire _36921 = _36917 ^ _36920;
  wire _36922 = _1302 ^ _14326;
  wire _36923 = _36922 ^ _23928;
  wire _36924 = _7680 ^ _464;
  wire _36925 = _4388 ^ _32009;
  wire _36926 = _36924 ^ _36925;
  wire _36927 = _36923 ^ _36926;
  wire _36928 = _36921 ^ _36927;
  wire _36929 = _5789 ^ _13822;
  wire _36930 = _12186 ^ _7094;
  wire _36931 = _36929 ^ _36930;
  wire _36932 = _4402 ^ _23945;
  wire _36933 = _36932 ^ _25757;
  wire _36934 = _36931 ^ _36933;
  wire _36935 = _486 ^ _4409;
  wire _36936 = _36935 ^ _33281;
  wire _36937 = _9996 ^ _35708;
  wire _36938 = uncoded_block[1027] ^ uncoded_block[1030];
  wire _36939 = _12752 ^ _36938;
  wire _36940 = _36937 ^ _36939;
  wire _36941 = _36936 ^ _36940;
  wire _36942 = _36934 ^ _36941;
  wire _36943 = _36928 ^ _36942;
  wire _36944 = _36913 ^ _36943;
  wire _36945 = _36886 ^ _36944;
  wire _36946 = _36826 ^ _36945;
  wire _36947 = _22131 ^ _17855;
  wire _36948 = _33284 ^ _36947;
  wire _36949 = uncoded_block[1056] ^ uncoded_block[1063];
  wire _36950 = _1359 ^ _36949;
  wire _36951 = _3689 ^ _3691;
  wire _36952 = _36950 ^ _36951;
  wire _36953 = _36948 ^ _36952;
  wire _36954 = _3692 ^ _3696;
  wire _36955 = uncoded_block[1091] ^ uncoded_block[1096];
  wire _36956 = _36955 ^ _5169;
  wire _36957 = _36954 ^ _36956;
  wire _36958 = _4450 ^ _8917;
  wire _36959 = _21690 ^ _36958;
  wire _36960 = _36957 ^ _36959;
  wire _36961 = _36953 ^ _36960;
  wire _36962 = _34533 ^ _1389;
  wire _36963 = _1392 ^ _19322;
  wire _36964 = _36962 ^ _36963;
  wire _36965 = _12794 ^ _20770;
  wire _36966 = _36964 ^ _36965;
  wire _36967 = _6505 ^ _2185;
  wire _36968 = uncoded_block[1153] ^ uncoded_block[1159];
  wire _36969 = _36968 ^ _2964;
  wire _36970 = _36967 ^ _36969;
  wire _36971 = _3736 ^ _11160;
  wire _36972 = _36971 ^ _22630;
  wire _36973 = _36970 ^ _36972;
  wire _36974 = _36966 ^ _36973;
  wire _36975 = _36961 ^ _36974;
  wire _36976 = _2967 ^ _3740;
  wire _36977 = _590 ^ _13882;
  wire _36978 = _36976 ^ _36977;
  wire _36979 = _593 ^ _24910;
  wire _36980 = _7160 ^ _5207;
  wire _36981 = _36979 ^ _36980;
  wire _36982 = _36978 ^ _36981;
  wire _36983 = _2216 ^ _26694;
  wire _36984 = _5889 ^ _2220;
  wire _36985 = _36983 ^ _36984;
  wire _36986 = uncoded_block[1232] ^ uncoded_block[1241];
  wire _36987 = _13357 ^ _36986;
  wire _36988 = _10062 ^ _36987;
  wire _36989 = _36985 ^ _36988;
  wire _36990 = _36982 ^ _36989;
  wire _36991 = _2995 ^ _3777;
  wire _36992 = _1451 ^ _5231;
  wire _36993 = _36991 ^ _36992;
  wire _36994 = _2236 ^ _3784;
  wire _36995 = _36994 ^ _21276;
  wire _36996 = _36993 ^ _36995;
  wire _36997 = _2247 ^ _631;
  wire _36998 = _12271 ^ _36997;
  wire _36999 = _4525 ^ _6560;
  wire _37000 = _639 ^ _4529;
  wire _37001 = _36999 ^ _37000;
  wire _37002 = _36998 ^ _37001;
  wire _37003 = _36996 ^ _37002;
  wire _37004 = _36990 ^ _37003;
  wire _37005 = _36975 ^ _37004;
  wire _37006 = _642 ^ _645;
  wire _37007 = _16424 ^ _3805;
  wire _37008 = _37006 ^ _37007;
  wire _37009 = _2261 ^ _21748;
  wire _37010 = _650 ^ _37009;
  wire _37011 = _37008 ^ _37010;
  wire _37012 = _21293 ^ _5254;
  wire _37013 = _4543 ^ _32513;
  wire _37014 = _37012 ^ _37013;
  wire _37015 = _6583 ^ _5268;
  wire _37016 = _5260 ^ _37015;
  wire _37017 = _37014 ^ _37016;
  wire _37018 = _37011 ^ _37017;
  wire _37019 = _5269 ^ _18436;
  wire _37020 = _5273 ^ _5275;
  wire _37021 = _37019 ^ _37020;
  wire _37022 = _13407 ^ _11776;
  wire _37023 = uncoded_block[1376] ^ uncoded_block[1380];
  wire _37024 = _10103 ^ _37023;
  wire _37025 = _37022 ^ _37024;
  wire _37026 = _37021 ^ _37025;
  wire _37027 = _22687 ^ _17953;
  wire _37028 = _37027 ^ _4570;
  wire _37029 = _5955 ^ _2297;
  wire _37030 = _15489 ^ _4580;
  wire _37031 = _37029 ^ _37030;
  wire _37032 = _37028 ^ _37031;
  wire _37033 = _37026 ^ _37032;
  wire _37034 = _37018 ^ _37033;
  wire _37035 = _1526 ^ _14466;
  wire _37036 = _706 ^ _37035;
  wire _37037 = _15980 ^ _10124;
  wire _37038 = _3857 ^ _2318;
  wire _37039 = _37037 ^ _37038;
  wire _37040 = _37036 ^ _37039;
  wire _37041 = _4590 ^ _3864;
  wire _37042 = _11246 ^ _2328;
  wire _37043 = _37041 ^ _37042;
  wire _37044 = _5309 ^ _12335;
  wire _37045 = _7243 ^ _10136;
  wire _37046 = _37044 ^ _37045;
  wire _37047 = _37043 ^ _37046;
  wire _37048 = _37040 ^ _37047;
  wire _37049 = _17976 ^ _4603;
  wire _37050 = uncoded_block[1481] ^ uncoded_block[1487];
  wire _37051 = _3881 ^ _37050;
  wire _37052 = _37049 ^ _37051;
  wire _37053 = _12899 ^ _4614;
  wire _37054 = _7253 ^ _37053;
  wire _37055 = _37052 ^ _37054;
  wire _37056 = _15002 ^ _31302;
  wire _37057 = uncoded_block[1522] ^ uncoded_block[1528];
  wire _37058 = _12352 ^ _37057;
  wire _37059 = _37056 ^ _37058;
  wire _37060 = _6002 ^ _12915;
  wire _37061 = _12917 ^ _16499;
  wire _37062 = _37060 ^ _37061;
  wire _37063 = _37059 ^ _37062;
  wire _37064 = _37055 ^ _37063;
  wire _37065 = _37048 ^ _37064;
  wire _37066 = _37034 ^ _37065;
  wire _37067 = _37005 ^ _37066;
  wire _37068 = _14496 ^ _769;
  wire _37069 = _24094 ^ _3139;
  wire _37070 = _37068 ^ _37069;
  wire _37071 = _17007 ^ _32567;
  wire _37072 = _36244 ^ _37071;
  wire _37073 = _37070 ^ _37072;
  wire _37074 = _5368 ^ _20401;
  wire _37075 = _6673 ^ _13996;
  wire _37076 = _37074 ^ _37075;
  wire _37077 = _12937 ^ _1625;
  wire _37078 = _37077 ^ _17018;
  wire _37079 = _37076 ^ _37078;
  wire _37080 = _37073 ^ _37079;
  wire _37081 = _10181 ^ _24115;
  wire _37082 = _7912 ^ _12947;
  wire _37083 = _37081 ^ _37082;
  wire _37084 = _1636 ^ _3166;
  wire _37085 = _7306 ^ _7309;
  wire _37086 = _37084 ^ _37085;
  wire _37087 = _37083 ^ _37086;
  wire _37088 = _33008 ^ _29567;
  wire _37089 = _3179 ^ _19470;
  wire _37090 = _3176 ^ _37089;
  wire _37091 = _37088 ^ _37090;
  wire _37092 = _37087 ^ _37091;
  wire _37093 = _37080 ^ _37092;
  wire _37094 = uncoded_block[1672] ^ uncoded_block[1677];
  wire _37095 = _37094 ^ _11321;
  wire _37096 = _10766 ^ _2427;
  wire _37097 = _37095 ^ _37096;
  wire _37098 = _837 ^ _1666;
  wire _37099 = _21394 ^ _25037;
  wire _37100 = _37098 ^ _37099;
  wire _37101 = _37097 ^ _37100;
  wire _37102 = _10215 ^ _7338;
  wire _37103 = _1677 ^ _3988;
  wire _37104 = _37103 ^ uncoded_block[1720];
  wire _37105 = _37102 ^ _37104;
  wire _37106 = _37101 ^ _37105;
  wire _37107 = _37093 ^ _37106;
  wire _37108 = _37067 ^ _37107;
  wire _37109 = _36946 ^ _37108;
  wire _37110 = _1 ^ _3212;
  wire _37111 = _37110 ^ _18059;
  wire _37112 = _8545 ^ _13537;
  wire _37113 = _7353 ^ _7959;
  wire _37114 = _37112 ^ _37113;
  wire _37115 = _37111 ^ _37114;
  wire _37116 = uncoded_block[31] ^ uncoded_block[35];
  wire _37117 = _11890 ^ _37116;
  wire _37118 = _8549 ^ _14571;
  wire _37119 = _37117 ^ _37118;
  wire _37120 = _7965 ^ _23;
  wire _37121 = _6099 ^ _21417;
  wire _37122 = _37120 ^ _37121;
  wire _37123 = _37119 ^ _37122;
  wire _37124 = _37115 ^ _37123;
  wire _37125 = _12996 ^ _1705;
  wire _37126 = _37125 ^ _25510;
  wire _37127 = uncoded_block[69] ^ uncoded_block[75];
  wire _37128 = _37127 ^ _3243;
  wire _37129 = uncoded_block[83] ^ uncoded_block[91];
  wire _37130 = _37129 ^ _22345;
  wire _37131 = _37128 ^ _37130;
  wire _37132 = _37126 ^ _37131;
  wire _37133 = _910 ^ _3250;
  wire _37134 = _37133 ^ _22350;
  wire _37135 = uncoded_block[113] ^ uncoded_block[117];
  wire _37136 = _37135 ^ _9721;
  wire _37137 = _37136 ^ _11375;
  wire _37138 = _37134 ^ _37137;
  wire _37139 = _37132 ^ _37138;
  wire _37140 = _37124 ^ _37139;
  wire _37141 = uncoded_block[131] ^ uncoded_block[136];
  wire _37142 = _37141 ^ _11918;
  wire _37143 = _11381 ^ _29204;
  wire _37144 = _37142 ^ _37143;
  wire _37145 = _1748 ^ _4053;
  wire _37146 = _8589 ^ _6788;
  wire _37147 = _37145 ^ _37146;
  wire _37148 = _37144 ^ _37147;
  wire _37149 = _21448 ^ _7403;
  wire _37150 = uncoded_block[182] ^ uncoded_block[189];
  wire _37151 = _37150 ^ _6798;
  wire _37152 = _37149 ^ _37151;
  wire _37153 = _9744 ^ _4068;
  wire _37154 = _12479 ^ _11405;
  wire _37155 = _37153 ^ _37154;
  wire _37156 = _37152 ^ _37155;
  wire _37157 = _37148 ^ _37156;
  wire _37158 = _34320 ^ _960;
  wire _37159 = _3298 ^ _4076;
  wire _37160 = _37158 ^ _37159;
  wire _37161 = _6168 ^ _6821;
  wire _37162 = _967 ^ _20994;
  wire _37163 = _37161 ^ _37162;
  wire _37164 = _37160 ^ _37163;
  wire _37165 = _5503 ^ _6179;
  wire _37166 = _974 ^ _11419;
  wire _37167 = _37165 ^ _37166;
  wire _37168 = uncoded_block[255] ^ uncoded_block[260];
  wire _37169 = _37168 ^ _6185;
  wire _37170 = _6187 ^ _985;
  wire _37171 = _37169 ^ _37170;
  wire _37172 = _37167 ^ _37171;
  wire _37173 = _37164 ^ _37172;
  wire _37174 = _37157 ^ _37173;
  wire _37175 = _37140 ^ _37174;
  wire _37176 = _26447 ^ _4105;
  wire _37177 = _991 ^ _13069;
  wire _37178 = _37176 ^ _37177;
  wire _37179 = _20038 ^ _29241;
  wire _37180 = _3334 ^ _6846;
  wire _37181 = _37179 ^ _37180;
  wire _37182 = _37178 ^ _37181;
  wire _37183 = _3346 ^ _8642;
  wire _37184 = _18146 ^ _37183;
  wire _37185 = _12521 ^ _4125;
  wire _37186 = uncoded_block[339] ^ uncoded_block[344];
  wire _37187 = _4126 ^ _37186;
  wire _37188 = _37185 ^ _37187;
  wire _37189 = _37184 ^ _37188;
  wire _37190 = _37182 ^ _37189;
  wire _37191 = _20050 ^ _8069;
  wire _37192 = _3362 ^ _3365;
  wire _37193 = _37191 ^ _37192;
  wire _37194 = _5548 ^ _17163;
  wire _37195 = _3369 ^ _13094;
  wire _37196 = _37194 ^ _37195;
  wire _37197 = _37193 ^ _37196;
  wire _37198 = _1841 ^ _3380;
  wire _37199 = _10900 ^ _37198;
  wire _37200 = _7483 ^ _19604;
  wire _37201 = _37200 ^ _23782;
  wire _37202 = _37199 ^ _37201;
  wire _37203 = _37197 ^ _37202;
  wire _37204 = _37190 ^ _37203;
  wire _37205 = uncoded_block[406] ^ uncoded_block[409];
  wire _37206 = _181 ^ _37205;
  wire _37207 = _11473 ^ _19612;
  wire _37208 = _37206 ^ _37207;
  wire _37209 = uncoded_block[424] ^ uncoded_block[432];
  wire _37210 = _37209 ^ _4169;
  wire _37211 = _15198 ^ _37210;
  wire _37212 = _37208 ^ _37211;
  wire _37213 = uncoded_block[443] ^ uncoded_block[448];
  wire _37214 = _5577 ^ _37213;
  wire _37215 = _37214 ^ _14171;
  wire _37216 = _212 ^ _3415;
  wire _37217 = _37216 ^ _35974;
  wire _37218 = _37215 ^ _37217;
  wire _37219 = _37212 ^ _37218;
  wire _37220 = _21523 ^ _4188;
  wire _37221 = _4189 ^ _3421;
  wire _37222 = _37220 ^ _37221;
  wire _37223 = _16693 ^ _6276;
  wire _37224 = _10370 ^ _8117;
  wire _37225 = _37223 ^ _37224;
  wire _37226 = _37222 ^ _37225;
  wire _37227 = _2668 ^ _2671;
  wire _37228 = _35981 ^ _37227;
  wire _37229 = _9294 ^ _10945;
  wire _37230 = uncoded_block[519] ^ uncoded_block[524];
  wire _37231 = _4910 ^ _37230;
  wire _37232 = _37229 ^ _37231;
  wire _37233 = _37228 ^ _37232;
  wire _37234 = _37226 ^ _37233;
  wire _37235 = _37219 ^ _37234;
  wire _37236 = _37204 ^ _37235;
  wire _37237 = _37175 ^ _37236;
  wire _37238 = _33162 ^ _4214;
  wire _37239 = _3451 ^ _7540;
  wire _37240 = _37238 ^ _37239;
  wire _37241 = _24282 ^ _8134;
  wire _37242 = _6940 ^ _3464;
  wire _37243 = _37241 ^ _37242;
  wire _37244 = _37240 ^ _37243;
  wire _37245 = _8731 ^ _1133;
  wire _37246 = _13699 ^ _37245;
  wire _37247 = uncoded_block[584] ^ uncoded_block[587];
  wire _37248 = _1138 ^ _37247;
  wire _37249 = _18222 ^ _6316;
  wire _37250 = _37248 ^ _37249;
  wire _37251 = _37246 ^ _37250;
  wire _37252 = _37244 ^ _37251;
  wire _37253 = uncoded_block[595] ^ uncoded_block[598];
  wire _37254 = _37253 ^ _4953;
  wire _37255 = _37254 ^ _10410;
  wire _37256 = _14218 ^ _14739;
  wire _37257 = _17232 ^ _7567;
  wire _37258 = _37256 ^ _37257;
  wire _37259 = _37255 ^ _37258;
  wire _37260 = _10980 ^ _7577;
  wire _37261 = _4965 ^ _37260;
  wire _37262 = _11543 ^ _1163;
  wire _37263 = _4972 ^ _19177;
  wire _37264 = _37262 ^ _37263;
  wire _37265 = _37261 ^ _37264;
  wire _37266 = _37259 ^ _37265;
  wire _37267 = _37252 ^ _37266;
  wire _37268 = _33190 ^ _16747;
  wire _37269 = _2739 ^ _12081;
  wire _37270 = _37268 ^ _37269;
  wire _37271 = _4265 ^ _3519;
  wire _37272 = _1968 ^ _319;
  wire _37273 = _37271 ^ _37272;
  wire _37274 = _37270 ^ _37273;
  wire _37275 = _13194 ^ _325;
  wire _37276 = _37275 ^ _6986;
  wire _37277 = _28542 ^ _9364;
  wire _37278 = _37276 ^ _37277;
  wire _37279 = _37274 ^ _37278;
  wire _37280 = _7597 ^ _5002;
  wire _37281 = _6367 ^ _18259;
  wire _37282 = _37280 ^ _37281;
  wire _37283 = uncoded_block[731] ^ uncoded_block[735];
  wire _37284 = _37283 ^ _13208;
  wire _37285 = _12652 ^ _37284;
  wire _37286 = _37282 ^ _37285;
  wire _37287 = uncoded_block[748] ^ uncoded_block[756];
  wire _37288 = _37287 ^ _13761;
  wire _37289 = _5703 ^ _37288;
  wire _37290 = _6382 ^ _12117;
  wire _37291 = _28181 ^ _37290;
  wire _37292 = _37289 ^ _37291;
  wire _37293 = _37286 ^ _37292;
  wire _37294 = _37279 ^ _37293;
  wire _37295 = _37267 ^ _37294;
  wire _37296 = _16786 ^ _5032;
  wire _37297 = _7022 ^ _37296;
  wire _37298 = _2019 ^ _3574;
  wire _37299 = _37298 ^ _16286;
  wire _37300 = _37297 ^ _37299;
  wire _37301 = _22071 ^ _16791;
  wire _37302 = _9396 ^ _2808;
  wire _37303 = _37301 ^ _37302;
  wire _37304 = _28197 ^ _1246;
  wire _37305 = _37304 ^ _36062;
  wire _37306 = _37303 ^ _37305;
  wire _37307 = _37300 ^ _37306;
  wire _37308 = _16293 ^ _5737;
  wire _37309 = _11609 ^ _3599;
  wire _37310 = _37308 ^ _37309;
  wire _37311 = _25711 ^ _21631;
  wire _37312 = _37311 ^ _14818;
  wire _37313 = _37310 ^ _37312;
  wire _37314 = _413 ^ _2828;
  wire _37315 = _35281 ^ _6416;
  wire _37316 = _37314 ^ _37315;
  wire _37317 = _11620 ^ _16815;
  wire _37318 = _20696 ^ _2838;
  wire _37319 = _37317 ^ _37318;
  wire _37320 = _37316 ^ _37319;
  wire _37321 = _37313 ^ _37320;
  wire _37322 = _37307 ^ _37321;
  wire _37323 = _4354 ^ _18307;
  wire _37324 = _25261 ^ _37323;
  wire _37325 = _4358 ^ _1281;
  wire _37326 = _1284 ^ _2071;
  wire _37327 = _37325 ^ _37326;
  wire _37328 = _37324 ^ _37327;
  wire _37329 = _7665 ^ _2852;
  wire _37330 = _37329 ^ _29818;
  wire _37331 = _4368 ^ _1295;
  wire _37332 = _37331 ^ _25270;
  wire _37333 = _37330 ^ _37332;
  wire _37334 = _37328 ^ _37333;
  wire _37335 = _453 ^ _23926;
  wire _37336 = _36509 ^ _37335;
  wire _37337 = uncoded_block[956] ^ uncoded_block[962];
  wire _37338 = _37337 ^ _10531;
  wire _37339 = _4383 ^ _37338;
  wire _37340 = _37336 ^ _37339;
  wire _37341 = uncoded_block[970] ^ uncoded_block[974];
  wire _37342 = _2093 ^ _37341;
  wire _37343 = _471 ^ _5790;
  wire _37344 = _37342 ^ _37343;
  wire _37345 = _8287 ^ _7094;
  wire _37346 = _8860 ^ _13277;
  wire _37347 = _37345 ^ _37346;
  wire _37348 = _37344 ^ _37347;
  wire _37349 = _37340 ^ _37348;
  wire _37350 = _37334 ^ _37349;
  wire _37351 = _37322 ^ _37350;
  wire _37352 = _37295 ^ _37351;
  wire _37353 = _37237 ^ _37352;
  wire _37354 = _5798 ^ _16343;
  wire _37355 = _4405 ^ _13283;
  wire _37356 = _37354 ^ _37355;
  wire _37357 = _1331 ^ _492;
  wire _37358 = _2894 ^ _11666;
  wire _37359 = _37357 ^ _37358;
  wire _37360 = _37356 ^ _37359;
  wire _37361 = _5806 ^ _5810;
  wire _37362 = _1346 ^ _2133;
  wire _37363 = _37361 ^ _37362;
  wire _37364 = _1360 ^ _4433;
  wire _37365 = _5148 ^ _37364;
  wire _37366 = _37363 ^ _37365;
  wire _37367 = _37360 ^ _37366;
  wire _37368 = _522 ^ _8889;
  wire _37369 = _1366 ^ _3692;
  wire _37370 = _37368 ^ _37369;
  wire _37371 = _5162 ^ _10575;
  wire _37372 = _37371 ^ _10020;
  wire _37373 = _37370 ^ _37372;
  wire _37374 = _5840 ^ _1378;
  wire _37375 = _37374 ^ _11694;
  wire _37376 = _7133 ^ _30326;
  wire _37377 = _2166 ^ _37376;
  wire _37378 = _37375 ^ _37377;
  wire _37379 = _37373 ^ _37378;
  wire _37380 = _37367 ^ _37379;
  wire _37381 = _2172 ^ _15894;
  wire _37382 = _13866 ^ _2177;
  wire _37383 = _37381 ^ _37382;
  wire _37384 = _567 ^ _1400;
  wire _37385 = _10597 ^ _8351;
  wire _37386 = _37384 ^ _37385;
  wire _37387 = _37383 ^ _37386;
  wire _37388 = uncoded_block[1165] ^ uncoded_block[1169];
  wire _37389 = _3734 ^ _37388;
  wire _37390 = _33323 ^ _37389;
  wire _37391 = _9506 ^ _13339;
  wire _37392 = _4481 ^ _590;
  wire _37393 = _37391 ^ _37392;
  wire _37394 = _37390 ^ _37393;
  wire _37395 = _37387 ^ _37394;
  wire _37396 = _5200 ^ _33330;
  wire _37397 = _37396 ^ _29891;
  wire _37398 = _12259 ^ _606;
  wire _37399 = _29892 ^ _37398;
  wire _37400 = _37397 ^ _37399;
  wire _37401 = _5215 ^ _609;
  wire _37402 = _34556 ^ _5218;
  wire _37403 = _37401 ^ _37402;
  wire _37404 = _15927 ^ _8382;
  wire _37405 = _11734 ^ _2997;
  wire _37406 = _37404 ^ _37405;
  wire _37407 = _37403 ^ _37406;
  wire _37408 = _37400 ^ _37407;
  wire _37409 = _37395 ^ _37408;
  wire _37410 = _37380 ^ _37409;
  wire _37411 = _3783 ^ _6550;
  wire _37412 = _25363 ^ _37411;
  wire _37413 = uncoded_block[1275] ^ uncoded_block[1282];
  wire _37414 = _37413 ^ _638;
  wire _37415 = _4524 ^ _37414;
  wire _37416 = _37412 ^ _37415;
  wire _37417 = _24023 ^ _641;
  wire _37418 = _37417 ^ _11198;
  wire _37419 = _6564 ^ _1479;
  wire _37420 = _8407 ^ _6574;
  wire _37421 = _37419 ^ _37420;
  wire _37422 = _37418 ^ _37421;
  wire _37423 = _37416 ^ _37422;
  wire _37424 = _12287 ^ _4543;
  wire _37425 = _21752 ^ _14437;
  wire _37426 = _37424 ^ _37425;
  wire _37427 = uncoded_block[1347] ^ uncoded_block[1351];
  wire _37428 = _11215 ^ _37427;
  wire _37429 = _19852 ^ _37428;
  wire _37430 = _37426 ^ _37429;
  wire _37431 = uncoded_block[1353] ^ uncoded_block[1360];
  wire _37432 = _37431 ^ _5275;
  wire _37433 = _2283 ^ _12302;
  wire _37434 = _37432 ^ _37433;
  wire _37435 = _17945 ^ _12305;
  wire _37436 = _11781 ^ _3061;
  wire _37437 = _37435 ^ _37436;
  wire _37438 = _37434 ^ _37437;
  wire _37439 = _37430 ^ _37438;
  wire _37440 = _37423 ^ _37439;
  wire _37441 = _29498 ^ _694;
  wire _37442 = _4572 ^ _26749;
  wire _37443 = _37441 ^ _37442;
  wire _37444 = _10681 ^ _26301;
  wire _37445 = _17959 ^ _37444;
  wire _37446 = _37443 ^ _37445;
  wire _37447 = _24969 ^ _27172;
  wire _37448 = _10124 ^ _24521;
  wire _37449 = _10130 ^ _8450;
  wire _37450 = _37448 ^ _37449;
  wire _37451 = _37447 ^ _37450;
  wire _37452 = _37446 ^ _37451;
  wire _37453 = _6620 ^ _19408;
  wire _37454 = _723 ^ _2335;
  wire _37455 = _37453 ^ _37454;
  wire _37456 = _3871 ^ _18919;
  wire _37457 = _11255 ^ _5316;
  wire _37458 = _37456 ^ _37457;
  wire _37459 = _37455 ^ _37458;
  wire _37460 = _5988 ^ _2349;
  wire _37461 = _1563 ^ _9614;
  wire _37462 = _37460 ^ _37461;
  wire _37463 = _24084 ^ _4616;
  wire _37464 = _16983 ^ _37463;
  wire _37465 = _37462 ^ _37464;
  wire _37466 = _37459 ^ _37465;
  wire _37467 = _37452 ^ _37466;
  wire _37468 = _37440 ^ _37467;
  wire _37469 = _37410 ^ _37468;
  wire _37470 = _9055 ^ _27621;
  wire _37471 = _9054 ^ _37470;
  wire _37472 = _1579 ^ _755;
  wire _37473 = _4623 ^ _9631;
  wire _37474 = _37472 ^ _37473;
  wire _37475 = _37471 ^ _37474;
  wire _37476 = _26789 ^ _13981;
  wire _37477 = uncoded_block[1553] ^ uncoded_block[1557];
  wire _37478 = _3912 ^ _37477;
  wire _37479 = _37478 ^ _7890;
  wire _37480 = _37476 ^ _37479;
  wire _37481 = _37475 ^ _37480;
  wire _37482 = _30869 ^ _30444;
  wire _37483 = _4651 ^ _10171;
  wire _37484 = _37483 ^ _9641;
  wire _37485 = _37482 ^ _37484;
  wire _37486 = _29994 ^ _14518;
  wire _37487 = _800 ^ _6040;
  wire _37488 = _3937 ^ _1633;
  wire _37489 = _37487 ^ _37488;
  wire _37490 = _37486 ^ _37489;
  wire _37491 = _37485 ^ _37490;
  wire _37492 = _37481 ^ _37491;
  wire _37493 = _12947 ^ _29147;
  wire _37494 = _20411 ^ _37493;
  wire _37495 = _12949 ^ _27651;
  wire _37496 = _6691 ^ _18030;
  wire _37497 = _37495 ^ _37496;
  wire _37498 = _37494 ^ _37497;
  wire _37499 = _14011 ^ _1653;
  wire _37500 = _25476 ^ _36269;
  wire _37501 = _37499 ^ _37500;
  wire _37502 = _833 ^ _4693;
  wire _37503 = _6705 ^ _3190;
  wire _37504 = _37502 ^ _37503;
  wire _37505 = _37501 ^ _37504;
  wire _37506 = _37498 ^ _37505;
  wire _37507 = _26832 ^ _15063;
  wire _37508 = _33020 ^ _37507;
  wire _37509 = _27671 ^ _1677;
  wire _37510 = _37509 ^ _21402;
  wire _37511 = _37508 ^ _37510;
  wire _37512 = _37506 ^ _37511;
  wire _37513 = _37492 ^ _37512;
  wire _37514 = _37469 ^ _37513;
  wire _37515 = _37353 ^ _37514;
  wire _37516 = _3209 ^ _866;
  wire _37517 = _6724 ^ _7956;
  wire _37518 = _37516 ^ _37517;
  wire _37519 = _8545 ^ _5426;
  wire _37520 = _35096 ^ _9143;
  wire _37521 = _37519 ^ _37520;
  wire _37522 = _37518 ^ _37521;
  wire _37523 = _15 ^ _14571;
  wire _37524 = _2468 ^ _888;
  wire _37525 = _37523 ^ _37524;
  wire _37526 = _10801 ^ _10806;
  wire _37527 = _9705 ^ _3241;
  wire _37528 = _37526 ^ _37527;
  wire _37529 = _37525 ^ _37528;
  wire _37530 = _37522 ^ _37529;
  wire _37531 = _7979 ^ _14586;
  wire _37532 = _37531 ^ _30933;
  wire _37533 = uncoded_block[99] ^ uncoded_block[105];
  wire _37534 = _46 ^ _37533;
  wire _37535 = _17580 ^ _37534;
  wire _37536 = _37532 ^ _37535;
  wire _37537 = uncoded_block[110] ^ uncoded_block[113];
  wire _37538 = _2491 ^ _37537;
  wire _37539 = _5455 ^ _12451;
  wire _37540 = _37538 ^ _37539;
  wire _37541 = _3257 ^ _11917;
  wire _37542 = _37540 ^ _37541;
  wire _37543 = _37536 ^ _37542;
  wire _37544 = _37530 ^ _37543;
  wire _37545 = _4760 ^ _5461;
  wire _37546 = _13573 ^ _70;
  wire _37547 = _37545 ^ _37546;
  wire _37548 = _3269 ^ _4048;
  wire _37549 = _37548 ^ _17601;
  wire _37550 = _37547 ^ _37549;
  wire _37551 = _30519 ^ _6788;
  wire _37552 = _37551 ^ _28035;
  wire _37553 = _10843 ^ _16114;
  wire _37554 = _4773 ^ _6800;
  wire _37555 = _37553 ^ _37554;
  wire _37556 = _37552 ^ _37555;
  wire _37557 = _37550 ^ _37556;
  wire _37558 = _95 ^ _1764;
  wire _37559 = _37558 ^ _27294;
  wire _37560 = _2540 ^ _9750;
  wire _37561 = _11409 ^ _2545;
  wire _37562 = _37560 ^ _37561;
  wire _37563 = _37559 ^ _37562;
  wire _37564 = _6168 ^ _1774;
  wire _37565 = _30087 ^ _7423;
  wire _37566 = _37564 ^ _37565;
  wire _37567 = _7425 ^ _4085;
  wire _37568 = _116 ^ _7434;
  wire _37569 = _37567 ^ _37568;
  wire _37570 = _37566 ^ _37569;
  wire _37571 = _37563 ^ _37570;
  wire _37572 = _37557 ^ _37571;
  wire _37573 = _37544 ^ _37572;
  wire _37574 = _4096 ^ _21007;
  wire _37575 = _22391 ^ _37574;
  wire _37576 = uncoded_block[282] ^ uncoded_block[287];
  wire _37577 = _5513 ^ _37576;
  wire _37578 = _21010 ^ _37577;
  wire _37579 = _37575 ^ _37578;
  wire _37580 = _992 ^ _16144;
  wire _37581 = uncoded_block[302] ^ uncoded_block[306];
  wire _37582 = _14133 ^ _37581;
  wire _37583 = _37580 ^ _37582;
  wire _37584 = _11439 ^ _4832;
  wire _37585 = _18613 ^ _37584;
  wire _37586 = _37583 ^ _37585;
  wire _37587 = _37579 ^ _37586;
  wire _37588 = uncoded_block[322] ^ uncoded_block[329];
  wire _37589 = _37588 ^ _15172;
  wire _37590 = _37589 ^ _12525;
  wire _37591 = uncoded_block[340] ^ uncoded_block[348];
  wire _37592 = _37591 ^ _5541;
  wire _37593 = _19092 ^ _33119;
  wire _37594 = _37592 ^ _37593;
  wire _37595 = _37590 ^ _37594;
  wire _37596 = _17163 ^ _3369;
  wire _37597 = _37596 ^ _21958;
  wire _37598 = _4854 ^ _4857;
  wire _37599 = _37598 ^ _9801;
  wire _37600 = _37597 ^ _37599;
  wire _37601 = _37595 ^ _37600;
  wire _37602 = _37587 ^ _37601;
  wire _37603 = _2615 ^ _3383;
  wire _37604 = _31870 ^ _1048;
  wire _37605 = _37603 ^ _37604;
  wire _37606 = _181 ^ _24243;
  wire _37607 = _37606 ^ _15198;
  wire _37608 = _37605 ^ _37607;
  wire _37609 = _21969 ^ _34374;
  wire _37610 = _10352 ^ _16187;
  wire _37611 = _37610 ^ _207;
  wire _37612 = _37609 ^ _37611;
  wire _37613 = _37608 ^ _37612;
  wire _37614 = _27756 ^ _2650;
  wire _37615 = _37614 ^ _8106;
  wire _37616 = _13665 ^ _221;
  wire _37617 = _15719 ^ _1086;
  wire _37618 = _37616 ^ _37617;
  wire _37619 = _37615 ^ _37618;
  wire _37620 = uncoded_block[490] ^ uncoded_block[493];
  wire _37621 = _7515 ^ _37620;
  wire _37622 = _30167 ^ _1097;
  wire _37623 = _37621 ^ _37622;
  wire _37624 = _2668 ^ _1892;
  wire _37625 = _37624 ^ _33579;
  wire _37626 = _37623 ^ _37625;
  wire _37627 = _37619 ^ _37626;
  wire _37628 = _37613 ^ _37627;
  wire _37629 = _37602 ^ _37628;
  wire _37630 = _37573 ^ _37629;
  wire _37631 = _8706 ^ _13152;
  wire _37632 = _37631 ^ _4923;
  wire _37633 = _9850 ^ _4217;
  wire _37634 = _9854 ^ _1909;
  wire _37635 = _37633 ^ _37634;
  wire _37636 = _37632 ^ _37635;
  wire _37637 = _2687 ^ _1123;
  wire _37638 = _3464 ^ _3467;
  wire _37639 = _37637 ^ _37638;
  wire _37640 = uncoded_block[568] ^ uncoded_block[574];
  wire _37641 = _37640 ^ _1931;
  wire _37642 = _37641 ^ _22013;
  wire _37643 = _37639 ^ _37642;
  wire _37644 = _37636 ^ _37643;
  wire _37645 = _9864 ^ _8148;
  wire _37646 = _37645 ^ _2708;
  wire _37647 = _3489 ^ _9870;
  wire _37648 = _12609 ^ _7564;
  wire _37649 = _37647 ^ _37648;
  wire _37650 = _37646 ^ _37649;
  wire _37651 = _3495 ^ _12618;
  wire _37652 = _13714 ^ _37651;
  wire _37653 = _1154 ^ _36847;
  wire _37654 = _1161 ^ _1956;
  wire _37655 = _37653 ^ _37654;
  wire _37656 = _37652 ^ _37655;
  wire _37657 = _37650 ^ _37656;
  wire _37658 = _37644 ^ _37657;
  wire _37659 = _6338 ^ _6341;
  wire _37660 = _37659 ^ _36021;
  wire _37661 = _16750 ^ _9357;
  wire _37662 = _37660 ^ _37661;
  wire _37663 = _6352 ^ _19191;
  wire _37664 = _322 ^ _13735;
  wire _37665 = _37663 ^ _37664;
  wire _37666 = _6985 ^ _19195;
  wire _37667 = _11562 ^ _6992;
  wire _37668 = _37666 ^ _37667;
  wire _37669 = _37665 ^ _37668;
  wire _37670 = _37662 ^ _37669;
  wire _37671 = uncoded_block[706] ^ uncoded_block[711];
  wire _37672 = _10447 ^ _37671;
  wire _37673 = _17266 ^ _6367;
  wire _37674 = _37672 ^ _37673;
  wire _37675 = _9369 ^ _3544;
  wire _37676 = _37675 ^ _12652;
  wire _37677 = _37674 ^ _37676;
  wire _37678 = uncoded_block[735] ^ uncoded_block[738];
  wire _37679 = _37678 ^ _5010;
  wire _37680 = _1209 ^ _37287;
  wire _37681 = _37679 ^ _37680;
  wire _37682 = _26579 ^ _13762;
  wire _37683 = _12113 ^ _34855;
  wire _37684 = _37682 ^ _37683;
  wire _37685 = _37681 ^ _37684;
  wire _37686 = _37677 ^ _37685;
  wire _37687 = _37670 ^ _37686;
  wire _37688 = _37658 ^ _37687;
  wire _37689 = _20165 ^ _19705;
  wire _37690 = _12673 ^ _4311;
  wire _37691 = _37689 ^ _37690;
  wire _37692 = uncoded_block[794] ^ uncoded_block[800];
  wire _37693 = _2019 ^ _37692;
  wire _37694 = _4317 ^ _16791;
  wire _37695 = _37693 ^ _37694;
  wire _37696 = _37691 ^ _37695;
  wire _37697 = _5042 ^ _2026;
  wire _37698 = uncoded_block[822] ^ uncoded_block[827];
  wire _37699 = _32388 ^ _37698;
  wire _37700 = _37697 ^ _37699;
  wire _37701 = uncoded_block[834] ^ uncoded_block[840];
  wire _37702 = _37701 ^ _2036;
  wire _37703 = _29793 ^ _37702;
  wire _37704 = _37700 ^ _37703;
  wire _37705 = _37696 ^ _37704;
  wire _37706 = _20188 ^ _2821;
  wire _37707 = _3600 ^ _2047;
  wire _37708 = _37706 ^ _37707;
  wire _37709 = uncoded_block[861] ^ uncoded_block[865];
  wire _37710 = _37709 ^ _5749;
  wire _37711 = _416 ^ _4347;
  wire _37712 = _37710 ^ _37711;
  wire _37713 = _37708 ^ _37712;
  wire _37714 = uncoded_block[896] ^ uncoded_block[901];
  wire _37715 = _5083 ^ _37714;
  wire _37716 = _19243 ^ _37715;
  wire _37717 = _1281 ^ _2070;
  wire _37718 = _19252 ^ _1287;
  wire _37719 = _37717 ^ _37718;
  wire _37720 = _37716 ^ _37719;
  wire _37721 = _37713 ^ _37720;
  wire _37722 = _37705 ^ _37721;
  wire _37723 = _3628 ^ _4368;
  wire _37724 = _37723 ^ _16829;
  wire _37725 = uncoded_block[936] ^ uncoded_block[942];
  wire _37726 = _449 ^ _37725;
  wire _37727 = uncoded_block[944] ^ uncoded_block[948];
  wire _37728 = _37727 ^ _4381;
  wire _37729 = _37726 ^ _37728;
  wire _37730 = _37724 ^ _37729;
  wire _37731 = _9438 ^ _14844;
  wire _37732 = _14330 ^ _37731;
  wire _37733 = _9981 ^ _22113;
  wire _37734 = _5114 ^ _11092;
  wire _37735 = _37733 ^ _37734;
  wire _37736 = _37732 ^ _37735;
  wire _37737 = _37730 ^ _37736;
  wire _37738 = _5790 ^ _1317;
  wire _37739 = _37738 ^ _34908;
  wire _37740 = _7691 ^ _6459;
  wire _37741 = _30293 ^ _37740;
  wire _37742 = _37739 ^ _37741;
  wire _37743 = uncoded_block[1011] ^ uncoded_block[1014];
  wire _37744 = _37743 ^ _5134;
  wire _37745 = _16853 ^ _12752;
  wire _37746 = _37744 ^ _37745;
  wire _37747 = _3675 ^ _34925;
  wire _37748 = _37747 ^ _8307;
  wire _37749 = _37746 ^ _37748;
  wire _37750 = _37742 ^ _37749;
  wire _37751 = _37737 ^ _37750;
  wire _37752 = _37722 ^ _37751;
  wire _37753 = _37688 ^ _37752;
  wire _37754 = _37630 ^ _37753;
  wire _37755 = uncoded_block[1050] ^ uncoded_block[1057];
  wire _37756 = _37755 ^ _521;
  wire _37757 = _35716 ^ _37756;
  wire _37758 = _8889 ^ _2143;
  wire _37759 = _23502 ^ _37758;
  wire _37760 = _37757 ^ _37759;
  wire _37761 = _20753 ^ _2149;
  wire _37762 = _12773 ^ _37761;
  wire _37763 = uncoded_block[1095] ^ uncoded_block[1102];
  wire _37764 = _31189 ^ _37763;
  wire _37765 = _37764 ^ _4449;
  wire _37766 = _37762 ^ _37765;
  wire _37767 = _37760 ^ _37766;
  wire _37768 = _550 ^ _1386;
  wire _37769 = _3713 ^ _14376;
  wire _37770 = _37768 ^ _37769;
  wire _37771 = _6500 ^ _8347;
  wire _37772 = _37770 ^ _37771;
  wire _37773 = _36139 ^ _5861;
  wire _37774 = _37773 ^ _18379;
  wire _37775 = _29439 ^ _8354;
  wire _37776 = _14389 ^ _2964;
  wire _37777 = _37775 ^ _37776;
  wire _37778 = _37774 ^ _37777;
  wire _37779 = _37772 ^ _37778;
  wire _37780 = _37767 ^ _37779;
  wire _37781 = _17390 ^ _9506;
  wire _37782 = _37781 ^ _32889;
  wire _37783 = _9508 ^ _2971;
  wire _37784 = _5879 ^ _37783;
  wire _37785 = _37782 ^ _37784;
  wire _37786 = _18389 ^ _23544;
  wire _37787 = _2204 ^ _37786;
  wire _37788 = uncoded_block[1216] ^ uncoded_block[1221];
  wire _37789 = _37788 ^ _2986;
  wire _37790 = _28298 ^ _37789;
  wire _37791 = _37787 ^ _37790;
  wire _37792 = _37785 ^ _37791;
  wire _37793 = _5894 ^ _14921;
  wire _37794 = _1443 ^ _10627;
  wire _37795 = _37793 ^ _37794;
  wire _37796 = uncoded_block[1243] ^ uncoded_block[1248];
  wire _37797 = _37796 ^ _11737;
  wire _37798 = _6546 ^ _7780;
  wire _37799 = _37797 ^ _37798;
  wire _37800 = _37795 ^ _37799;
  wire _37801 = _8970 ^ _22197;
  wire _37802 = _37801 ^ _30364;
  wire _37803 = _21281 ^ _24931;
  wire _37804 = _37802 ^ _37803;
  wire _37805 = _37800 ^ _37804;
  wire _37806 = _37792 ^ _37805;
  wire _37807 = _37780 ^ _37806;
  wire _37808 = _5243 ^ _24482;
  wire _37809 = _37808 ^ _25378;
  wire _37810 = _35380 ^ _3805;
  wire _37811 = _37810 ^ _10088;
  wire _37812 = _37809 ^ _37811;
  wire _37813 = uncoded_block[1321] ^ uncoded_block[1324];
  wire _37814 = _21293 ^ _37813;
  wire _37815 = _7201 ^ _23139;
  wire _37816 = _37814 ^ _37815;
  wire _37817 = _3820 ^ _3034;
  wire _37818 = _5261 ^ _13927;
  wire _37819 = _37817 ^ _37818;
  wire _37820 = _37816 ^ _37819;
  wire _37821 = _37812 ^ _37820;
  wire _37822 = _669 ^ _5272;
  wire _37823 = _673 ^ _22223;
  wire _37824 = _37822 ^ _37823;
  wire _37825 = _11224 ^ _11776;
  wire _37826 = _12305 ^ _29083;
  wire _37827 = _37825 ^ _37826;
  wire _37828 = _37824 ^ _37827;
  wire _37829 = _12311 ^ _691;
  wire _37830 = _694 ^ _5955;
  wire _37831 = _37829 ^ _37830;
  wire _37832 = _12315 ^ _4578;
  wire _37833 = _37832 ^ _5958;
  wire _37834 = _37831 ^ _37833;
  wire _37835 = _37828 ^ _37834;
  wire _37836 = _37821 ^ _37835;
  wire _37837 = uncoded_block[1421] ^ uncoded_block[1427];
  wire _37838 = _10120 ^ _37837;
  wire _37839 = _19399 ^ _37838;
  wire _37840 = _5968 ^ _10124;
  wire _37841 = _24521 ^ _27175;
  wire _37842 = _37840 ^ _37841;
  wire _37843 = _37839 ^ _37842;
  wire _37844 = uncoded_block[1448] ^ uncoded_block[1454];
  wire _37845 = _37844 ^ _3088;
  wire _37846 = _5313 ^ _18919;
  wire _37847 = _37845 ^ _37846;
  wire _37848 = _4603 ^ _1555;
  wire _37849 = _37848 ^ _14994;
  wire _37850 = _37847 ^ _37849;
  wire _37851 = _37843 ^ _37850;
  wire _37852 = _1563 ^ _13967;
  wire _37853 = _743 ^ _1571;
  wire _37854 = _37852 ^ _37853;
  wire _37855 = _18478 ^ _19892;
  wire _37856 = _7875 ^ _9621;
  wire _37857 = _37855 ^ _37856;
  wire _37858 = _37854 ^ _37857;
  wire _37859 = _9058 ^ _3900;
  wire _37860 = _5343 ^ _24994;
  wire _37861 = _37859 ^ _37860;
  wire _37862 = _15009 ^ _20387;
  wire _37863 = uncoded_block[1548] ^ uncoded_block[1556];
  wire _37864 = _2367 ^ _37863;
  wire _37865 = _37862 ^ _37864;
  wire _37866 = _37861 ^ _37865;
  wire _37867 = _37858 ^ _37866;
  wire _37868 = _37851 ^ _37867;
  wire _37869 = _37836 ^ _37868;
  wire _37870 = _37807 ^ _37869;
  wire _37871 = uncoded_block[1565] ^ uncoded_block[1567];
  wire _37872 = _773 ^ _37871;
  wire _37873 = _5363 ^ _21361;
  wire _37874 = _37872 ^ _37873;
  wire _37875 = _1615 ^ _25454;
  wire _37876 = _11839 ^ _37875;
  wire _37877 = _37874 ^ _37876;
  wire _37878 = _792 ^ _29550;
  wire _37879 = _12937 ^ _20406;
  wire _37880 = _37878 ^ _37879;
  wire _37881 = _9089 ^ _16031;
  wire _37882 = _37881 ^ _37081;
  wire _37883 = _37880 ^ _37882;
  wire _37884 = _37877 ^ _37883;
  wire _37885 = _6684 ^ _4665;
  wire _37886 = _37885 ^ _6687;
  wire _37887 = _2407 ^ _9661;
  wire _37888 = _20417 ^ _13508;
  wire _37889 = _37887 ^ _37888;
  wire _37890 = _37886 ^ _37889;
  wire _37891 = _4680 ^ _3175;
  wire _37892 = uncoded_block[1667] ^ uncoded_block[1672];
  wire _37893 = _7319 ^ _37892;
  wire _37894 = _37891 ^ _37893;
  wire _37895 = uncoded_block[1676] ^ uncoded_block[1681];
  wire _37896 = _8522 ^ _37895;
  wire _37897 = _37896 ^ _4695;
  wire _37898 = _37894 ^ _37897;
  wire _37899 = _37890 ^ _37898;
  wire _37900 = _37884 ^ _37899;
  wire _37901 = _28422 ^ _15064;
  wire _37902 = _33022 ^ _14030;
  wire _37903 = _37901 ^ _37902;
  wire _37904 = _37903 ^ uncoded_block[1722];
  wire _37905 = _37900 ^ _37904;
  wire _37906 = _37870 ^ _37905;
  wire _37907 = _37754 ^ _37906;
  wire _37908 = _4710 ^ _866;
  wire _37909 = _19959 ^ _19001;
  wire _37910 = _37908 ^ _37909;
  wire _37911 = _3998 ^ _872;
  wire _37912 = _9143 ^ _31363;
  wire _37913 = _37911 ^ _37912;
  wire _37914 = _37910 ^ _37913;
  wire _37915 = _21871 ^ _22;
  wire _37916 = _34281 ^ _37915;
  wire _37917 = _8554 ^ _13547;
  wire _37918 = _888 ^ _31790;
  wire _37919 = _37917 ^ _37918;
  wire _37920 = _37916 ^ _37919;
  wire _37921 = _37914 ^ _37920;
  wire _37922 = _34289 ^ _7367;
  wire _37923 = uncoded_block[72] ^ uncoded_block[79];
  wire _37924 = _37923 ^ _20472;
  wire _37925 = _37922 ^ _37924;
  wire _37926 = _15101 ^ _50;
  wire _37927 = _35114 ^ _37926;
  wire _37928 = _37925 ^ _37927;
  wire _37929 = _3253 ^ _33056;
  wire _37930 = _12451 ^ _33058;
  wire _37931 = _37929 ^ _37930;
  wire _37932 = _18095 ^ _15114;
  wire _37933 = _24172 ^ _37932;
  wire _37934 = _37931 ^ _37933;
  wire _37935 = _37928 ^ _37934;
  wire _37936 = _37921 ^ _37935;
  wire _37937 = _14082 ^ _10262;
  wire _37938 = _2514 ^ _8589;
  wire _37939 = _37937 ^ _37938;
  wire _37940 = _11390 ^ _4057;
  wire _37941 = _9195 ^ _4772;
  wire _37942 = _37940 ^ _37941;
  wire _37943 = _37939 ^ _37942;
  wire _37944 = _16116 ^ _8018;
  wire _37945 = _14096 ^ _37944;
  wire _37946 = _10278 ^ _14101;
  wire _37947 = _5489 ^ _2540;
  wire _37948 = _37946 ^ _37947;
  wire _37949 = _37945 ^ _37948;
  wire _37950 = _37943 ^ _37949;
  wire _37951 = _9750 ^ _8606;
  wire _37952 = _37951 ^ _19554;
  wire _37953 = _2550 ^ _6824;
  wire _37954 = _4082 ^ _37953;
  wire _37955 = _37952 ^ _37954;
  wire _37956 = _10860 ^ _35145;
  wire _37957 = _2556 ^ _13053;
  wire _37958 = _37956 ^ _37957;
  wire _37959 = uncoded_block[261] ^ uncoded_block[268];
  wire _37960 = _37959 ^ _16636;
  wire _37961 = _30098 ^ _37960;
  wire _37962 = _37958 ^ _37961;
  wire _37963 = _37955 ^ _37962;
  wire _37964 = _37950 ^ _37963;
  wire _37965 = _37936 ^ _37964;
  wire _37966 = _21479 ^ _4814;
  wire _37967 = _4105 ^ _15159;
  wire _37968 = _37966 ^ _37967;
  wire _37969 = _14652 ^ _3337;
  wire _37970 = _35160 ^ _37969;
  wire _37971 = _37968 ^ _37970;
  wire _37972 = _17642 ^ _4830;
  wire _37973 = _4832 ^ _15677;
  wire _37974 = _37972 ^ _37973;
  wire _37975 = _30117 ^ _2586;
  wire _37976 = _37975 ^ _10324;
  wire _37977 = _37974 ^ _37976;
  wire _37978 = _37971 ^ _37977;
  wire _37979 = _11450 ^ _6218;
  wire _37980 = _8652 ^ _13089;
  wire _37981 = _37979 ^ _37980;
  wire _37982 = _35170 ^ _1032;
  wire _37983 = uncoded_block[368] ^ uncoded_block[374];
  wire _37984 = _37983 ^ _10898;
  wire _37985 = _37982 ^ _37984;
  wire _37986 = _37981 ^ _37985;
  wire _37987 = _10899 ^ _6876;
  wire _37988 = uncoded_block[390] ^ uncoded_block[395];
  wire _37989 = _9255 ^ _37988;
  wire _37990 = _37987 ^ _37989;
  wire _37991 = uncoded_block[399] ^ uncoded_block[403];
  wire _37992 = _10910 ^ _37991;
  wire _37993 = _26045 ^ _3394;
  wire _37994 = _37992 ^ _37993;
  wire _37995 = _37990 ^ _37994;
  wire _37996 = _37986 ^ _37995;
  wire _37997 = _37978 ^ _37996;
  wire _37998 = _13112 ^ _14160;
  wire _37999 = _12551 ^ _14163;
  wire _38000 = _37998 ^ _37999;
  wire _38001 = _2638 ^ _201;
  wire _38002 = _5574 ^ _21052;
  wire _38003 = _38001 ^ _38002;
  wire _38004 = _38000 ^ _38003;
  wire _38005 = _1069 ^ _4883;
  wire _38006 = _38005 ^ _214;
  wire _38007 = _4890 ^ _21059;
  wire _38008 = _35973 ^ _38007;
  wire _38009 = _38006 ^ _38008;
  wire _38010 = _38004 ^ _38009;
  wire _38011 = _4188 ^ _24723;
  wire _38012 = _38011 ^ _9831;
  wire _38013 = _5600 ^ _27769;
  wire _38014 = _8698 ^ _25167;
  wire _38015 = _38013 ^ _38014;
  wire _38016 = _38012 ^ _38015;
  wire _38017 = _7531 ^ _9298;
  wire _38018 = _38017 ^ _29713;
  wire _38019 = _239 ^ _9309;
  wire _38020 = uncoded_block[540] ^ uncoded_block[547];
  wire _38021 = _6932 ^ _38020;
  wire _38022 = _38019 ^ _38021;
  wire _38023 = _38018 ^ _38022;
  wire _38024 = _38016 ^ _38023;
  wire _38025 = _38010 ^ _38024;
  wire _38026 = _37997 ^ _38025;
  wire _38027 = _37965 ^ _38026;
  wire _38028 = _23382 ^ _8724;
  wire _38029 = uncoded_block[562] ^ uncoded_block[566];
  wire _38030 = _4937 ^ _38029;
  wire _38031 = _38028 ^ _38030;
  wire _38032 = uncoded_block[567] ^ uncoded_block[573];
  wire _38033 = _38032 ^ _8731;
  wire _38034 = _38033 ^ _23834;
  wire _38035 = _38031 ^ _38034;
  wire _38036 = _35220 ^ _1141;
  wire _38037 = _38036 ^ _28516;
  wire _38038 = _4952 ^ _274;
  wire _38039 = _4240 ^ _17232;
  wire _38040 = _38038 ^ _38039;
  wire _38041 = _38037 ^ _38040;
  wire _38042 = _38035 ^ _38041;
  wire _38043 = _6960 ^ _4963;
  wire _38044 = _19663 ^ _38043;
  wire _38045 = _17238 ^ _30199;
  wire _38046 = uncoded_block[635] ^ uncoded_block[637];
  wire _38047 = _38046 ^ _6969;
  wire _38048 = _38045 ^ _38047;
  wire _38049 = _38044 ^ _38048;
  wire _38050 = _8751 ^ _6338;
  wire _38051 = _19177 ^ _6974;
  wire _38052 = _38050 ^ _38051;
  wire _38053 = _16249 ^ _3513;
  wire _38054 = _5670 ^ _15273;
  wire _38055 = _38053 ^ _38054;
  wire _38056 = _38052 ^ _38055;
  wire _38057 = _38049 ^ _38056;
  wire _38058 = _38042 ^ _38057;
  wire _38059 = _15775 ^ _319;
  wire _38060 = _5678 ^ _1974;
  wire _38061 = _38059 ^ _38060;
  wire _38062 = _18250 ^ _30214;
  wire _38063 = _20654 ^ _11565;
  wire _38064 = _38062 ^ _38063;
  wire _38065 = _38061 ^ _38064;
  wire _38066 = _12647 ^ _18259;
  wire _38067 = _2768 ^ _7002;
  wire _38068 = _38066 ^ _38067;
  wire _38069 = _1203 ^ _28930;
  wire _38070 = _35254 ^ _4298;
  wire _38071 = _38069 ^ _38070;
  wire _38072 = _38068 ^ _38071;
  wire _38073 = _38065 ^ _38072;
  wire _38074 = uncoded_block[768] ^ uncoded_block[778];
  wire _38075 = _364 ^ _38074;
  wire _38076 = _12673 ^ _371;
  wire _38077 = _38075 ^ _38076;
  wire _38078 = uncoded_block[787] ^ uncoded_block[791];
  wire _38079 = _38078 ^ _3574;
  wire _38080 = _14282 ^ _3576;
  wire _38081 = _38079 ^ _38080;
  wire _38082 = _38077 ^ _38081;
  wire _38083 = _32799 ^ _2026;
  wire _38084 = _35265 ^ _38083;
  wire _38085 = _7037 ^ _3587;
  wire _38086 = _33655 ^ _38085;
  wire _38087 = _38084 ^ _38086;
  wire _38088 = _38082 ^ _38087;
  wire _38089 = _38073 ^ _38088;
  wire _38090 = _38058 ^ _38089;
  wire _38091 = _12135 ^ _34467;
  wire _38092 = _9938 ^ _9405;
  wire _38093 = _38091 ^ _38092;
  wire _38094 = _6407 ^ _32809;
  wire _38095 = _38093 ^ _38094;
  wire _38096 = _2827 ^ _2830;
  wire _38097 = _26166 ^ _38096;
  wire _38098 = _36903 ^ _423;
  wire _38099 = _15338 ^ _38098;
  wire _38100 = _38097 ^ _38099;
  wire _38101 = _38095 ^ _38100;
  wire _38102 = _20701 ^ _29808;
  wire _38103 = _12156 ^ _38102;
  wire _38104 = _10508 ^ _2850;
  wire _38105 = _5762 ^ _18775;
  wire _38106 = _38104 ^ _38105;
  wire _38107 = _38103 ^ _38106;
  wire _38108 = _35296 ^ _2078;
  wire _38109 = _5101 ^ _7673;
  wire _38110 = _38108 ^ _38109;
  wire _38111 = _8271 ^ _23926;
  wire _38112 = _13266 ^ _8275;
  wire _38113 = _38111 ^ _38112;
  wire _38114 = _38110 ^ _38113;
  wire _38115 = _38107 ^ _38114;
  wire _38116 = _38101 ^ _38115;
  wire _38117 = _1307 ^ _25741;
  wire _38118 = _9981 ^ _8847;
  wire _38119 = _38117 ^ _38118;
  wire _38120 = _4397 ^ _8856;
  wire _38121 = _4396 ^ _38120;
  wire _38122 = _38119 ^ _38121;
  wire _38123 = uncoded_block[993] ^ uncoded_block[999];
  wire _38124 = _38123 ^ _24858;
  wire _38125 = _34913 ^ _4410;
  wire _38126 = _38124 ^ _38125;
  wire _38127 = _2894 ^ _5137;
  wire _38128 = _34107 ^ _38127;
  wire _38129 = _38126 ^ _38128;
  wire _38130 = _38122 ^ _38129;
  wire _38131 = _12752 ^ _498;
  wire _38132 = _12756 ^ _6474;
  wire _38133 = _38131 ^ _38132;
  wire _38134 = _19295 ^ _5147;
  wire _38135 = _23956 ^ _38134;
  wire _38136 = _38133 ^ _38135;
  wire _38137 = uncoded_block[1056] ^ uncoded_block[1059];
  wire _38138 = _4430 ^ _38137;
  wire _38139 = _3685 ^ _25773;
  wire _38140 = _38138 ^ _38139;
  wire _38141 = uncoded_block[1082] ^ uncoded_block[1087];
  wire _38142 = _2147 ^ _38141;
  wire _38143 = _27511 ^ _38142;
  wire _38144 = _38140 ^ _38143;
  wire _38145 = _38136 ^ _38144;
  wire _38146 = _38130 ^ _38145;
  wire _38147 = _38116 ^ _38146;
  wire _38148 = _38090 ^ _38147;
  wire _38149 = _38027 ^ _38148;
  wire _38150 = _1378 ^ _11139;
  wire _38151 = _36550 ^ _38150;
  wire _38152 = _12224 ^ _13318;
  wire _38153 = _38152 ^ _7134;
  wire _38154 = _38151 ^ _38153;
  wire _38155 = _5175 ^ _4455;
  wire _38156 = _8345 ^ _10593;
  wire _38157 = _38155 ^ _38156;
  wire _38158 = _16380 ^ _2953;
  wire _38159 = _38158 ^ _14892;
  wire _38160 = _38157 ^ _38159;
  wire _38161 = _38154 ^ _38160;
  wire _38162 = _2185 ^ _33736;
  wire _38163 = _38162 ^ _16892;
  wire _38164 = _5869 ^ _2967;
  wire _38165 = _38164 ^ _23991;
  wire _38166 = _38163 ^ _38165;
  wire _38167 = _33330 ^ _596;
  wire _38168 = _26688 ^ _38167;
  wire _38169 = uncoded_block[1197] ^ uncoded_block[1203];
  wire _38170 = uncoded_block[1204] ^ uncoded_block[1208];
  wire _38171 = _38169 ^ _38170;
  wire _38172 = _38171 ^ _35361;
  wire _38173 = _38168 ^ _38172;
  wire _38174 = _38166 ^ _38173;
  wire _38175 = _38161 ^ _38174;
  wire _38176 = _1436 ^ _31228;
  wire _38177 = _35363 ^ _38176;
  wire _38178 = _11732 ^ _10627;
  wire _38179 = _1449 ^ _1451;
  wire _38180 = _38178 ^ _38179;
  wire _38181 = _38177 ^ _38180;
  wire _38182 = _7178 ^ _627;
  wire _38183 = _7779 ^ _38182;
  wire _38184 = _7788 ^ _26718;
  wire _38185 = _30789 ^ _23123;
  wire _38186 = _38184 ^ _38185;
  wire _38187 = _38183 ^ _38186;
  wire _38188 = _38181 ^ _38187;
  wire _38189 = _25376 ^ _16423;
  wire _38190 = _14939 ^ _1479;
  wire _38191 = _29064 ^ _38190;
  wire _38192 = _38189 ^ _38191;
  wire _38193 = _14432 ^ _21293;
  wire _38194 = _35386 ^ _38193;
  wire _38195 = _8413 ^ _3822;
  wire _38196 = _17935 ^ _38195;
  wire _38197 = _38194 ^ _38196;
  wire _38198 = _38192 ^ _38197;
  wire _38199 = _38188 ^ _38198;
  wire _38200 = _38175 ^ _38199;
  wire _38201 = _10092 ^ _11218;
  wire _38202 = _5938 ^ _16942;
  wire _38203 = _38201 ^ _38202;
  wire _38204 = _5273 ^ _21306;
  wire _38205 = uncoded_block[1369] ^ uncoded_block[1375];
  wire _38206 = _38205 ^ _7217;
  wire _38207 = _38204 ^ _38206;
  wire _38208 = _38203 ^ _38207;
  wire _38209 = _16451 ^ _23154;
  wire _38210 = _692 ^ _694;
  wire _38211 = _38209 ^ _38210;
  wire _38212 = uncoded_block[1403] ^ uncoded_block[1409];
  wire _38213 = _5293 ^ _38212;
  wire _38214 = _38213 ^ _34601;
  wire _38215 = _38211 ^ _38214;
  wire _38216 = _38208 ^ _38215;
  wire _38217 = uncoded_block[1419] ^ uncoded_block[1423];
  wire _38218 = _38217 ^ _14466;
  wire _38219 = _38218 ^ _35415;
  wire _38220 = uncoded_block[1442] ^ uncoded_block[1448];
  wire _38221 = _38220 ^ _3865;
  wire _38222 = _21785 ^ _38221;
  wire _38223 = _38219 ^ _38222;
  wire _38224 = _22250 ^ _31285;
  wire _38225 = _726 ^ _5314;
  wire _38226 = _11255 ^ _1558;
  wire _38227 = _38225 ^ _38226;
  wire _38228 = _38224 ^ _38227;
  wire _38229 = _38223 ^ _38228;
  wire _38230 = _38216 ^ _38229;
  wire _38231 = uncoded_block[1484] ^ uncoded_block[1492];
  wire _38232 = _38231 ^ _12896;
  wire _38233 = _38232 ^ _9047;
  wire _38234 = _3111 ^ _23190;
  wire _38235 = _7875 ^ _5337;
  wire _38236 = _38234 ^ _38235;
  wire _38237 = _38233 ^ _38236;
  wire _38238 = _8473 ^ _13459;
  wire _38239 = _10717 ^ _38238;
  wire _38240 = uncoded_block[1534] ^ uncoded_block[1540];
  wire _38241 = _38240 ^ _7883;
  wire _38242 = _18488 ^ _38241;
  wire _38243 = _38239 ^ _38242;
  wire _38244 = _38237 ^ _38243;
  wire _38245 = _5355 ^ _13472;
  wire _38246 = _38245 ^ _31312;
  wire _38247 = uncoded_block[1558] ^ uncoded_block[1564];
  wire _38248 = uncoded_block[1565] ^ uncoded_block[1571];
  wire _38249 = _38247 ^ _38248;
  wire _38250 = _13478 ^ _6663;
  wire _38251 = _38249 ^ _38250;
  wire _38252 = _38246 ^ _38251;
  wire _38253 = _15537 ^ _1615;
  wire _38254 = _15030 ^ _38253;
  wire _38255 = _3145 ^ _12935;
  wire _38256 = _8499 ^ _6039;
  wire _38257 = _38255 ^ _38256;
  wire _38258 = _38254 ^ _38257;
  wire _38259 = _38252 ^ _38258;
  wire _38260 = _38244 ^ _38259;
  wire _38261 = _38230 ^ _38260;
  wire _38262 = _38200 ^ _38261;
  wire _38263 = _6677 ^ _12940;
  wire _38264 = _16032 ^ _805;
  wire _38265 = _38263 ^ _38264;
  wire _38266 = _13494 ^ _3161;
  wire _38267 = _3166 ^ _6049;
  wire _38268 = _38266 ^ _38267;
  wire _38269 = _38265 ^ _38268;
  wire _38270 = _3172 ^ _4678;
  wire _38271 = _33005 ^ _38270;
  wire _38272 = _1654 ^ _2422;
  wire _38273 = _9109 ^ _38272;
  wire _38274 = _38271 ^ _38273;
  wire _38275 = _38269 ^ _38274;
  wire _38276 = _3182 ^ _8522;
  wire _38277 = _7325 ^ _13517;
  wire _38278 = _38276 ^ _38277;
  wire _38279 = uncoded_block[1694] ^ uncoded_block[1700];
  wire _38280 = _3190 ^ _38279;
  wire _38281 = _34660 ^ _38280;
  wire _38282 = _38278 ^ _38281;
  wire _38283 = _30024 ^ _36700;
  wire _38284 = _38283 ^ uncoded_block[1718];
  wire _38285 = _38282 ^ _38284;
  wire _38286 = _38275 ^ _38285;
  wire _38287 = _38262 ^ _38286;
  wire _38288 = _38149 ^ _38287;
  wire _38289 = _4710 ^ _32201;
  wire _38290 = _6083 ^ _3998;
  wire _38291 = _38289 ^ _38290;
  wire _38292 = _4716 ^ _27998;
  wire _38293 = _13539 ^ _2462;
  wire _38294 = _38292 ^ _38293;
  wire _38295 = _38291 ^ _38294;
  wire _38296 = _21871 ^ _20457;
  wire _38297 = _32211 ^ _4726;
  wire _38298 = _38296 ^ _38297;
  wire _38299 = uncoded_block[54] ^ uncoded_block[57];
  wire _38300 = _38299 ^ _10806;
  wire _38301 = _38300 ^ _7368;
  wire _38302 = _38298 ^ _38301;
  wire _38303 = _38295 ^ _38302;
  wire _38304 = _12438 ^ _6749;
  wire _38305 = _35111 ^ _6755;
  wire _38306 = _38304 ^ _38305;
  wire _38307 = _17081 ^ _29608;
  wire _38308 = _38306 ^ _38307;
  wire _38309 = _15102 ^ _25519;
  wire _38310 = _7990 ^ _54;
  wire _38311 = _12451 ^ _9727;
  wire _38312 = _38310 ^ _38311;
  wire _38313 = _38309 ^ _38312;
  wire _38314 = _38308 ^ _38313;
  wire _38315 = _38303 ^ _38314;
  wire _38316 = _9729 ^ _2511;
  wire _38317 = _17594 ^ _38316;
  wire _38318 = uncoded_block[150] ^ uncoded_block[155];
  wire _38319 = _38318 ^ _12463;
  wire _38320 = uncoded_block[171] ^ uncoded_block[177];
  wire _38321 = _8589 ^ _38320;
  wire _38322 = _38319 ^ _38321;
  wire _38323 = _38317 ^ _38322;
  wire _38324 = _4770 ^ _13583;
  wire _38325 = _38324 ^ _35902;
  wire _38326 = uncoded_block[191] ^ uncoded_block[197];
  wire _38327 = _4773 ^ _38326;
  wire _38328 = _2537 ^ _4070;
  wire _38329 = _38327 ^ _38328;
  wire _38330 = _38325 ^ _38329;
  wire _38331 = _38323 ^ _38330;
  wire _38332 = uncoded_block[206] ^ uncoded_block[210];
  wire _38333 = _38332 ^ _19549;
  wire _38334 = _3296 ^ _102;
  wire _38335 = _38333 ^ _38334;
  wire _38336 = _104 ^ _3299;
  wire _38337 = _109 ^ _16125;
  wire _38338 = _38336 ^ _38337;
  wire _38339 = _38335 ^ _38338;
  wire _38340 = uncoded_block[237] ^ uncoded_block[241];
  wire _38341 = _38340 ^ _11952;
  wire _38342 = _38341 ^ _23304;
  wire _38343 = _11419 ^ _14639;
  wire _38344 = _38343 ^ _20521;
  wire _38345 = _38342 ^ _38344;
  wire _38346 = _38339 ^ _38345;
  wire _38347 = _38331 ^ _38346;
  wire _38348 = _38315 ^ _38347;
  wire _38349 = _20523 ^ _33099;
  wire _38350 = _38349 ^ _21010;
  wire _38351 = uncoded_block[281] ^ uncoded_block[289];
  wire _38352 = _38351 ^ _10876;
  wire _38353 = _6195 ^ _38352;
  wire _38354 = _38350 ^ _38353;
  wire _38355 = _2573 ^ _142;
  wire _38356 = _15668 ^ _3338;
  wire _38357 = _38355 ^ _38356;
  wire _38358 = _15168 ^ _2580;
  wire _38359 = _9780 ^ _2586;
  wire _38360 = _38358 ^ _38359;
  wire _38361 = _38357 ^ _38360;
  wire _38362 = _38354 ^ _38361;
  wire _38363 = uncoded_block[338] ^ uncoded_block[345];
  wire _38364 = _38363 ^ _1023;
  wire _38365 = _35556 ^ _38364;
  wire _38366 = uncoded_block[349] ^ uncoded_block[356];
  wire _38367 = _38366 ^ _6864;
  wire _38368 = _12530 ^ _21955;
  wire _38369 = _38367 ^ _38368;
  wire _38370 = _38365 ^ _38369;
  wire _38371 = _10896 ^ _4144;
  wire _38372 = _28091 ^ _10908;
  wire _38373 = _28845 ^ _26925;
  wire _38374 = _38372 ^ _38373;
  wire _38375 = _38371 ^ _38374;
  wire _38376 = _38370 ^ _38375;
  wire _38377 = _38362 ^ _38376;
  wire _38378 = _1051 ^ _5564;
  wire _38379 = _4161 ^ _14160;
  wire _38380 = _38378 ^ _38379;
  wire _38381 = _24248 ^ _6894;
  wire _38382 = _38381 ^ _10353;
  wire _38383 = _38380 ^ _38382;
  wire _38384 = _3404 ^ _5578;
  wire _38385 = _1864 ^ _19118;
  wire _38386 = _38384 ^ _38385;
  wire _38387 = _1079 ^ _12023;
  wire _38388 = _13128 ^ _38387;
  wire _38389 = _38386 ^ _38388;
  wire _38390 = _38383 ^ _38389;
  wire _38391 = _8110 ^ _21528;
  wire _38392 = _35588 ^ _38391;
  wire _38393 = _8117 ^ _1094;
  wire _38394 = _7517 ^ _38393;
  wire _38395 = _38392 ^ _38394;
  wire _38396 = _1097 ^ _6921;
  wire _38397 = uncoded_block[509] ^ uncoded_block[513];
  wire _38398 = _6922 ^ _38397;
  wire _38399 = _38396 ^ _38398;
  wire _38400 = uncoded_block[514] ^ uncoded_block[525];
  wire _38401 = _38400 ^ _4922;
  wire _38402 = _4925 ^ _10384;
  wire _38403 = _38401 ^ _38402;
  wire _38404 = _38399 ^ _38403;
  wire _38405 = _38395 ^ _38404;
  wire _38406 = _38390 ^ _38405;
  wire _38407 = _38377 ^ _38406;
  wire _38408 = _38348 ^ _38407;
  wire _38409 = _16215 ^ _3451;
  wire _38410 = _16715 ^ _6300;
  wire _38411 = _38409 ^ _38410;
  wire _38412 = _22004 ^ _15740;
  wire _38413 = _31907 ^ _9320;
  wire _38414 = _38412 ^ _38413;
  wire _38415 = _38411 ^ _38414;
  wire _38416 = _5635 ^ _6309;
  wire _38417 = _17221 ^ _4941;
  wire _38418 = _38416 ^ _38417;
  wire _38419 = _265 ^ _22012;
  wire _38420 = _38419 ^ _33602;
  wire _38421 = _38418 ^ _38420;
  wire _38422 = _38415 ^ _38421;
  wire _38423 = _18225 ^ _4953;
  wire _38424 = _3487 ^ _277;
  wire _38425 = _38423 ^ _38424;
  wire _38426 = _21098 ^ _3494;
  wire _38427 = _14222 ^ _38426;
  wire _38428 = _38425 ^ _38427;
  wire _38429 = uncoded_block[621] ^ uncoded_block[633];
  wire _38430 = _38429 ^ _4249;
  wire _38431 = _2727 ^ _6338;
  wire _38432 = _38430 ^ _38431;
  wire _38433 = _28908 ^ _8755;
  wire _38434 = _3514 ^ _308;
  wire _38435 = _38433 ^ _38434;
  wire _38436 = _38432 ^ _38435;
  wire _38437 = _38428 ^ _38436;
  wire _38438 = _38422 ^ _38437;
  wire _38439 = uncoded_block[667] ^ uncoded_block[672];
  wire _38440 = _1173 ^ _38439;
  wire _38441 = _17745 ^ _1181;
  wire _38442 = _38440 ^ _38441;
  wire _38443 = _6353 ^ _15281;
  wire _38444 = _38443 ^ _29755;
  wire _38445 = _38442 ^ _38444;
  wire _38446 = _6985 ^ _3529;
  wire _38447 = _4989 ^ _8189;
  wire _38448 = _38446 ^ _38447;
  wire _38449 = _4996 ^ _19201;
  wire _38450 = uncoded_block[717] ^ uncoded_block[720];
  wire _38451 = _38450 ^ _15292;
  wire _38452 = _38449 ^ _38451;
  wire _38453 = _38448 ^ _38452;
  wire _38454 = _38445 ^ _38453;
  wire _38455 = _4286 ^ _1991;
  wire _38456 = _38455 ^ _2771;
  wire _38457 = _1210 ^ _5016;
  wire _38458 = _20666 ^ _38457;
  wire _38459 = _38456 ^ _38458;
  wire _38460 = _1215 ^ _7016;
  wire _38461 = _38460 ^ _18744;
  wire _38462 = uncoded_block[772] ^ uncoded_block[777];
  wire _38463 = _11019 ^ _38462;
  wire _38464 = uncoded_block[778] ^ uncoded_block[782];
  wire _38465 = _38464 ^ _3570;
  wire _38466 = _38463 ^ _38465;
  wire _38467 = _38461 ^ _38466;
  wire _38468 = _38459 ^ _38467;
  wire _38469 = _38454 ^ _38468;
  wire _38470 = _38438 ^ _38469;
  wire _38471 = _1232 ^ _24804;
  wire _38472 = _1226 ^ _38471;
  wire _38473 = _4317 ^ _1238;
  wire _38474 = _38473 ^ _12681;
  wire _38475 = _38472 ^ _38474;
  wire _38476 = _4325 ^ _1242;
  wire _38477 = uncoded_block[827] ^ uncoded_block[833];
  wire _38478 = _397 ^ _38477;
  wire _38479 = _38476 ^ _38478;
  wire _38480 = _16293 ^ _4337;
  wire _38481 = uncoded_block[840] ^ uncoded_block[845];
  wire _38482 = _38481 ^ _19725;
  wire _38483 = _38480 ^ _38482;
  wire _38484 = _38479 ^ _38483;
  wire _38485 = _38475 ^ _38484;
  wire _38486 = _20692 ^ _9948;
  wire _38487 = _30257 ^ _38486;
  wire _38488 = _2828 ^ _416;
  wire _38489 = _14303 ^ _38488;
  wire _38490 = _38487 ^ _38489;
  wire _38491 = _2831 ^ _16815;
  wire _38492 = _16304 ^ _2054;
  wire _38493 = _38491 ^ _38492;
  wire _38494 = _11060 ^ _34081;
  wire _38495 = _38494 ^ _13803;
  wire _38496 = _38493 ^ _38495;
  wire _38497 = _38490 ^ _38496;
  wire _38498 = _38485 ^ _38497;
  wire _38499 = _7070 ^ _435;
  wire _38500 = uncoded_block[921] ^ uncoded_block[928];
  wire _38501 = _3631 ^ _38500;
  wire _38502 = _38499 ^ _38501;
  wire _38503 = _8835 ^ _2862;
  wire _38504 = uncoded_block[941] ^ uncoded_block[946];
  wire _38505 = _2083 ^ _38504;
  wire _38506 = _38503 ^ _38505;
  wire _38507 = _38502 ^ _38506;
  wire _38508 = _29387 ^ _5779;
  wire _38509 = _38508 ^ _34095;
  wire _38510 = _15363 ^ _468;
  wire _38511 = _16330 ^ _38510;
  wire _38512 = _38509 ^ _38511;
  wire _38513 = _38507 ^ _38512;
  wire _38514 = _17836 ^ _7689;
  wire _38515 = _1317 ^ _23938;
  wire _38516 = _38514 ^ _38515;
  wire _38517 = uncoded_block[998] ^ uncoded_block[1001];
  wire _38518 = _18333 ^ _38517;
  wire _38519 = _2112 ^ _2114;
  wire _38520 = _38518 ^ _38519;
  wire _38521 = _38516 ^ _38520;
  wire _38522 = _36532 ^ _35708;
  wire _38523 = _36106 ^ _38522;
  wire _38524 = uncoded_block[1022] ^ uncoded_block[1027];
  wire _38525 = _38524 ^ _26653;
  wire _38526 = _12199 ^ _12208;
  wire _38527 = _38525 ^ _38526;
  wire _38528 = _38523 ^ _38527;
  wire _38529 = _38521 ^ _38528;
  wire _38530 = _38513 ^ _38529;
  wire _38531 = _38498 ^ _38530;
  wire _38532 = _38470 ^ _38531;
  wire _38533 = _38408 ^ _38532;
  wire _38534 = _2134 ^ _2136;
  wire _38535 = uncoded_block[1058] ^ uncoded_block[1064];
  wire _38536 = _9465 ^ _38535;
  wire _38537 = _38534 ^ _38536;
  wire _38538 = uncoded_block[1066] ^ uncoded_block[1073];
  wire _38539 = _38538 ^ _6486;
  wire _38540 = _20251 ^ _2149;
  wire _38541 = _38539 ^ _38540;
  wire _38542 = _38537 ^ _38541;
  wire _38543 = _31189 ^ _10026;
  wire _38544 = _18365 ^ _546;
  wire _38545 = _38543 ^ _38544;
  wire _38546 = _3711 ^ _4451;
  wire _38547 = _23075 ^ _553;
  wire _38548 = _38546 ^ _38547;
  wire _38549 = _38545 ^ _38548;
  wire _38550 = _38542 ^ _38549;
  wire _38551 = _16376 ^ _15894;
  wire _38552 = _8343 ^ _13869;
  wire _38553 = _38551 ^ _38552;
  wire _38554 = _4465 ^ _27532;
  wire _38555 = _17381 ^ _38554;
  wire _38556 = _38553 ^ _38555;
  wire _38557 = uncoded_block[1152] ^ uncoded_block[1156];
  wire _38558 = _38557 ^ _24442;
  wire _38559 = _38558 ^ _3737;
  wire _38560 = _17392 ^ _4481;
  wire _38561 = uncoded_block[1182] ^ uncoded_block[1186];
  wire _38562 = _590 ^ _38561;
  wire _38563 = _38560 ^ _38562;
  wire _38564 = _38559 ^ _38563;
  wire _38565 = _38556 ^ _38564;
  wire _38566 = _38550 ^ _38565;
  wire _38567 = _2200 ^ _21257;
  wire _38568 = _1421 ^ _2974;
  wire _38569 = _38567 ^ _38568;
  wire _38570 = _1425 ^ _11171;
  wire _38571 = _1428 ^ _5889;
  wire _38572 = _38570 ^ _38571;
  wire _38573 = _38569 ^ _38572;
  wire _38574 = uncoded_block[1219] ^ uncoded_block[1224];
  wire _38575 = _38574 ^ _12819;
  wire _38576 = _38575 ^ _12266;
  wire _38577 = _30355 ^ _6546;
  wire _38578 = _35761 ^ _38577;
  wire _38579 = _38576 ^ _38578;
  wire _38580 = _38573 ^ _38579;
  wire _38581 = _3784 ^ _5235;
  wire _38582 = _13902 ^ _38581;
  wire _38583 = _7791 ^ _3793;
  wire _38584 = _19835 ^ _38583;
  wire _38585 = _38582 ^ _38584;
  wire _38586 = _23123 ^ _3797;
  wire _38587 = _5913 ^ _4529;
  wire _38588 = _38586 ^ _38587;
  wire _38589 = _645 ^ _8984;
  wire _38590 = uncoded_block[1306] ^ uncoded_block[1310];
  wire _38591 = _1472 ^ _38590;
  wire _38592 = _38589 ^ _38591;
  wire _38593 = _38588 ^ _38592;
  wire _38594 = _38585 ^ _38593;
  wire _38595 = _38580 ^ _38594;
  wire _38596 = _38566 ^ _38595;
  wire _38597 = _14430 ^ _9552;
  wire _38598 = _38597 ^ _24491;
  wire _38599 = uncoded_block[1329] ^ uncoded_block[1335];
  wire _38600 = _4545 ^ _38599;
  wire _38601 = _2276 ^ _1497;
  wire _38602 = _38600 ^ _38601;
  wire _38603 = _38598 ^ _38602;
  wire _38604 = _29929 ^ _18435;
  wire _38605 = _5272 ^ _23581;
  wire _38606 = uncoded_block[1368] ^ uncoded_block[1375];
  wire _38607 = _32106 ^ _38606;
  wire _38608 = _38605 ^ _38607;
  wire _38609 = _38604 ^ _38608;
  wire _38610 = _38603 ^ _38609;
  wire _38611 = _5284 ^ _9575;
  wire _38612 = _38611 ^ _20338;
  wire _38613 = uncoded_block[1392] ^ uncoded_block[1395];
  wire _38614 = _38613 ^ _30821;
  wire _38615 = _38614 ^ _5958;
  wire _38616 = _38612 ^ _38615;
  wire _38617 = _5961 ^ _20347;
  wire _38618 = _8438 ^ _17960;
  wire _38619 = _38617 ^ _38618;
  wire _38620 = _1526 ^ _3075;
  wire _38621 = _17468 ^ _2314;
  wire _38622 = _38620 ^ _38621;
  wire _38623 = _38619 ^ _38622;
  wire _38624 = _38616 ^ _38623;
  wire _38625 = _38610 ^ _38624;
  wire _38626 = uncoded_block[1443] ^ uncoded_block[1447];
  wire _38627 = _4590 ^ _38626;
  wire _38628 = _38627 ^ _26310;
  wire _38629 = _13437 ^ _21793;
  wire _38630 = _29519 ^ _4603;
  wire _38631 = _38629 ^ _38630;
  wire _38632 = _38628 ^ _38631;
  wire _38633 = _3881 ^ _1558;
  wire _38634 = _25426 ^ _13967;
  wire _38635 = _38633 ^ _38634;
  wire _38636 = uncoded_block[1499] ^ uncoded_block[1505];
  wire _38637 = _743 ^ _38636;
  wire _38638 = uncoded_block[1508] ^ uncoded_block[1511];
  wire _38639 = _3112 ^ _38638;
  wire _38640 = _38637 ^ _38639;
  wire _38641 = _38635 ^ _38640;
  wire _38642 = _38632 ^ _38641;
  wire _38643 = _9053 ^ _751;
  wire _38644 = _9058 ^ _17499;
  wire _38645 = _38643 ^ _38644;
  wire _38646 = _5344 ^ _12915;
  wire _38647 = uncoded_block[1538] ^ uncoded_block[1543];
  wire _38648 = _38647 ^ _4634;
  wire _38649 = _38646 ^ _38648;
  wire _38650 = _38645 ^ _38649;
  wire _38651 = _12920 ^ _22731;
  wire _38652 = _1597 ^ _774;
  wire _38653 = _38651 ^ _38652;
  wire _38654 = _20392 ^ _1606;
  wire _38655 = _18949 ^ _3924;
  wire _38656 = _38654 ^ _38655;
  wire _38657 = _38653 ^ _38656;
  wire _38658 = _38650 ^ _38657;
  wire _38659 = _38642 ^ _38658;
  wire _38660 = _38625 ^ _38659;
  wire _38661 = _38596 ^ _38660;
  wire _38662 = _30875 ^ _6674;
  wire _38663 = _38662 ^ _12374;
  wire _38664 = _1627 ^ _7908;
  wire _38665 = _25905 ^ _9095;
  wire _38666 = _38664 ^ _38665;
  wire _38667 = _38663 ^ _38666;
  wire _38668 = uncoded_block[1622] ^ uncoded_block[1627];
  wire _38669 = _38668 ^ _1636;
  wire _38670 = _5388 ^ _4668;
  wire _38671 = _38669 ^ _38670;
  wire _38672 = _4672 ^ _7313;
  wire _38673 = _38671 ^ _38672;
  wire _38674 = _38667 ^ _38673;
  wire _38675 = _4677 ^ _1653;
  wire _38676 = _38675 ^ _14535;
  wire _38677 = _9666 ^ _7928;
  wire _38678 = _11319 ^ _7325;
  wire _38679 = _38677 ^ _38678;
  wire _38680 = _38676 ^ _38679;
  wire _38681 = _10766 ^ _17040;
  wire _38682 = _11324 ^ _9675;
  wire _38683 = _38681 ^ _38682;
  wire _38684 = _9677 ^ _6068;
  wire _38685 = _38684 ^ _20921;
  wire _38686 = _38683 ^ _38685;
  wire _38687 = _38680 ^ _38686;
  wire _38688 = _38674 ^ _38687;
  wire _38689 = _1677 ^ _2444;
  wire _38690 = _38689 ^ uncoded_block[1722];
  wire _38691 = _38688 ^ _38690;
  wire _38692 = _38661 ^ _38691;
  wire _38693 = _38533 ^ _38692;
  wire _38694 = _22785 ^ _28746;
  wire _38695 = _15076 ^ _9694;
  wire _38696 = _11890 ^ _3227;
  wire _38697 = _38695 ^ _38696;
  wire _38698 = _38694 ^ _38697;
  wire _38699 = _21871 ^ _12425;
  wire _38700 = _8554 ^ _6101;
  wire _38701 = _38699 ^ _38700;
  wire _38702 = _5436 ^ _13552;
  wire _38703 = _7365 ^ _9705;
  wire _38704 = _38702 ^ _38703;
  wire _38705 = _38701 ^ _38704;
  wire _38706 = _38698 ^ _38705;
  wire _38707 = _35 ^ _897;
  wire _38708 = _38707 ^ _9709;
  wire _38709 = _13004 ^ _6755;
  wire _38710 = _15603 ^ _6115;
  wire _38711 = _38709 ^ _38710;
  wire _38712 = _38708 ^ _38711;
  wire _38713 = uncoded_block[100] ^ uncoded_block[103];
  wire _38714 = _38713 ^ _6120;
  wire _38715 = _48 ^ _38714;
  wire _38716 = _6122 ^ _20957;
  wire _38717 = _38716 ^ _18565;
  wire _38718 = _38715 ^ _38717;
  wire _38719 = _38712 ^ _38718;
  wire _38720 = _38706 ^ _38719;
  wire _38721 = uncoded_block[123] ^ uncoded_block[128];
  wire _38722 = _2501 ^ _38721;
  wire _38723 = uncoded_block[131] ^ uncoded_block[134];
  wire _38724 = _923 ^ _38723;
  wire _38725 = _38722 ^ _38724;
  wire _38726 = _8581 ^ _927;
  wire _38727 = _10830 ^ _14082;
  wire _38728 = _38726 ^ _38727;
  wire _38729 = _38725 ^ _38728;
  wire _38730 = _6782 ^ _19999;
  wire _38731 = _8589 ^ _2521;
  wire _38732 = _2522 ^ _940;
  wire _38733 = _38731 ^ _38732;
  wire _38734 = _38730 ^ _38733;
  wire _38735 = _38729 ^ _38734;
  wire _38736 = _1759 ^ _4773;
  wire _38737 = _5480 ^ _38736;
  wire _38738 = _9744 ^ _952;
  wire _38739 = _14101 ^ _3292;
  wire _38740 = _38738 ^ _38739;
  wire _38741 = _38737 ^ _38740;
  wire _38742 = uncoded_block[214] ^ uncoded_block[222];
  wire _38743 = _38742 ^ _8608;
  wire _38744 = _4081 ^ _2550;
  wire _38745 = _38743 ^ _38744;
  wire _38746 = _9756 ^ _10860;
  wire _38747 = _30090 ^ _38746;
  wire _38748 = _38745 ^ _38747;
  wire _38749 = _38741 ^ _38748;
  wire _38750 = _38735 ^ _38749;
  wire _38751 = _38720 ^ _38750;
  wire _38752 = _5505 ^ _14116;
  wire _38753 = _11419 ^ _1786;
  wire _38754 = _38752 ^ _38753;
  wire _38755 = uncoded_block[262] ^ uncoded_block[265];
  wire _38756 = _38755 ^ _7440;
  wire _38757 = _14642 ^ _6192;
  wire _38758 = _38756 ^ _38757;
  wire _38759 = _38754 ^ _38758;
  wire _38760 = _988 ^ _134;
  wire _38761 = _6195 ^ _38760;
  wire _38762 = uncoded_block[289] ^ uncoded_block[292];
  wire _38763 = _38762 ^ _24216;
  wire _38764 = _1810 ^ _12515;
  wire _38765 = _38763 ^ _38764;
  wire _38766 = _38761 ^ _38765;
  wire _38767 = _38759 ^ _38766;
  wire _38768 = _15668 ^ _8056;
  wire _38769 = _38768 ^ _11440;
  wire _38770 = _12520 ^ _35555;
  wire _38771 = _38769 ^ _38770;
  wire _38772 = _4838 ^ _11984;
  wire _38773 = _3355 ^ _2599;
  wire _38774 = _38772 ^ _38773;
  wire _38775 = _19092 ^ _2602;
  wire _38776 = _38775 ^ _21031;
  wire _38777 = _38774 ^ _38776;
  wire _38778 = _38771 ^ _38777;
  wire _38779 = _38767 ^ _38778;
  wire _38780 = _18161 ^ _19596;
  wire _38781 = _1841 ^ _31005;
  wire _38782 = _38781 ^ _22421;
  wire _38783 = _38780 ^ _38782;
  wire _38784 = _3388 ^ _5559;
  wire _38785 = uncoded_block[412] ^ uncoded_block[417];
  wire _38786 = _184 ^ _38785;
  wire _38787 = _38784 ^ _38786;
  wire _38788 = uncoded_block[425] ^ uncoded_block[431];
  wire _38789 = _8671 ^ _38788;
  wire _38790 = _25598 ^ _38789;
  wire _38791 = _38787 ^ _38790;
  wire _38792 = _38783 ^ _38791;
  wire _38793 = _4169 ^ _1863;
  wire _38794 = _13122 ^ _6259;
  wire _38795 = _38793 ^ _38794;
  wire _38796 = _4883 ^ _2650;
  wire _38797 = _7504 ^ _4181;
  wire _38798 = _38796 ^ _38797;
  wire _38799 = _38795 ^ _38798;
  wire _38800 = _13666 ^ _8109;
  wire _38801 = _1085 ^ _12028;
  wire _38802 = _38801 ^ _17197;
  wire _38803 = _38800 ^ _38802;
  wire _38804 = _38799 ^ _38803;
  wire _38805 = _38792 ^ _38804;
  wire _38806 = _38779 ^ _38805;
  wire _38807 = _38751 ^ _38806;
  wire _38808 = _3424 ^ _2665;
  wire _38809 = _2667 ^ _3434;
  wire _38810 = _38808 ^ _38809;
  wire _38811 = uncoded_block[509] ^ uncoded_block[518];
  wire _38812 = _5611 ^ _38811;
  wire _38813 = _18201 ^ _38812;
  wire _38814 = _38810 ^ _38813;
  wire _38815 = uncoded_block[524] ^ uncoded_block[529];
  wire _38816 = _8708 ^ _38815;
  wire _38817 = _38816 ^ _35603;
  wire _38818 = _25173 ^ _16715;
  wire _38819 = _38818 ^ _6302;
  wire _38820 = _38817 ^ _38819;
  wire _38821 = _38814 ^ _38820;
  wire _38822 = _1122 ^ _4937;
  wire _38823 = _5633 ^ _18682;
  wire _38824 = _38822 ^ _38823;
  wire _38825 = _8731 ^ _16727;
  wire _38826 = uncoded_block[587] ^ uncoded_block[592];
  wire _38827 = _31915 ^ _38826;
  wire _38828 = _38825 ^ _38827;
  wire _38829 = _38824 ^ _38828;
  wire _38830 = _6316 ^ _8149;
  wire _38831 = _9868 ^ _277;
  wire _38832 = _38830 ^ _38831;
  wire _38833 = _6323 ^ _17232;
  wire _38834 = _8744 ^ _4243;
  wire _38835 = _38833 ^ _38834;
  wire _38836 = _38832 ^ _38835;
  wire _38837 = _38829 ^ _38836;
  wire _38838 = _38821 ^ _38837;
  wire _38839 = _7568 ^ _8159;
  wire _38840 = _289 ^ _7577;
  wire _38841 = _38839 ^ _38840;
  wire _38842 = _294 ^ _15766;
  wire _38843 = _301 ^ _304;
  wire _38844 = _38842 ^ _38843;
  wire _38845 = _38841 ^ _38844;
  wire _38846 = uncoded_block[660] ^ uncoded_block[665];
  wire _38847 = _2738 ^ _38846;
  wire _38848 = _38847 ^ _4266;
  wire _38849 = _8177 ^ _10440;
  wire _38850 = _18247 ^ _321;
  wire _38851 = _38849 ^ _38850;
  wire _38852 = _38848 ^ _38851;
  wire _38853 = _38845 ^ _38852;
  wire _38854 = _18249 ^ _2754;
  wire _38855 = _2755 ^ _6360;
  wire _38856 = _38854 ^ _38855;
  wire _38857 = _333 ^ _33204;
  wire _38858 = _31525 ^ _1195;
  wire _38859 = _38857 ^ _38858;
  wire _38860 = _38856 ^ _38859;
  wire _38861 = _11006 ^ _5006;
  wire _38862 = _1206 ^ _1996;
  wire _38863 = _38861 ^ _38862;
  wire _38864 = _7601 ^ _38863;
  wire _38865 = _38860 ^ _38864;
  wire _38866 = _38853 ^ _38865;
  wire _38867 = _38838 ^ _38866;
  wire _38868 = _352 ^ _3550;
  wire _38869 = _1999 ^ _6378;
  wire _38870 = _38868 ^ _38869;
  wire _38871 = _15796 ^ _4302;
  wire _38872 = _38870 ^ _38871;
  wire _38873 = _5027 ^ _14271;
  wire _38874 = _31545 ^ _5715;
  wire _38875 = _38873 ^ _38874;
  wire _38876 = _3574 ^ _7029;
  wire _38877 = _38876 ^ _34063;
  wire _38878 = _38875 ^ _38877;
  wire _38879 = _38872 ^ _38878;
  wire _38880 = _15318 ^ _22525;
  wire _38881 = _27843 ^ _2032;
  wire _38882 = _38880 ^ _38881;
  wire _38883 = _15324 ^ _401;
  wire _38884 = _3591 ^ _38883;
  wire _38885 = _38882 ^ _38884;
  wire _38886 = _4337 ^ _10495;
  wire _38887 = _10498 ^ _2046;
  wire _38888 = _38886 ^ _38887;
  wire _38889 = uncoded_block[859] ^ uncoded_block[865];
  wire _38890 = _14300 ^ _38889;
  wire _38891 = _38890 ^ _33670;
  wire _38892 = _38888 ^ _38891;
  wire _38893 = _38885 ^ _38892;
  wire _38894 = _38879 ^ _38893;
  wire _38895 = _6416 ^ _5078;
  wire _38896 = _16304 ^ _2058;
  wire _38897 = _38895 ^ _38896;
  wire _38898 = uncoded_block[887] ^ uncoded_block[892];
  wire _38899 = _38898 ^ _2062;
  wire _38900 = _38899 ^ _21176;
  wire _38901 = _38897 ^ _38900;
  wire _38902 = uncoded_block[908] ^ uncoded_block[920];
  wire _38903 = _2065 ^ _38902;
  wire _38904 = _445 ^ _2076;
  wire _38905 = _38903 ^ _38904;
  wire _38906 = _448 ^ _8262;
  wire _38907 = _15355 ^ _456;
  wire _38908 = _38906 ^ _38907;
  wire _38909 = _38905 ^ _38908;
  wire _38910 = _38901 ^ _38909;
  wire _38911 = _5777 ^ _461;
  wire _38912 = _1308 ^ _10529;
  wire _38913 = _38911 ^ _38912;
  wire _38914 = _14844 ^ _9981;
  wire _38915 = uncoded_block[971] ^ uncoded_block[975];
  wire _38916 = _7088 ^ _38915;
  wire _38917 = _38914 ^ _38916;
  wire _38918 = _38913 ^ _38917;
  wire _38919 = _5789 ^ _29832;
  wire _38920 = _7093 ^ _24853;
  wire _38921 = _38919 ^ _38920;
  wire _38922 = _16846 ^ _16342;
  wire _38923 = _38921 ^ _38922;
  wire _38924 = _38918 ^ _38923;
  wire _38925 = _38910 ^ _38924;
  wire _38926 = _38894 ^ _38925;
  wire _38927 = _38867 ^ _38926;
  wire _38928 = _38807 ^ _38927;
  wire _38929 = uncoded_block[1002] ^ uncoded_block[1005];
  wire _38930 = _38929 ^ _2886;
  wire _38931 = _15860 ^ _19763;
  wire _38932 = _38930 ^ _38931;
  wire _38933 = _8872 ^ _18801;
  wire _38934 = _33705 ^ _38933;
  wire _38935 = _38932 ^ _38934;
  wire _38936 = _5806 ^ _12198;
  wire _38937 = uncoded_block[1041] ^ uncoded_block[1043];
  wire _38938 = _1345 ^ _38937;
  wire _38939 = _38936 ^ _38938;
  wire _38940 = _514 ^ _2134;
  wire _38941 = _38940 ^ _23501;
  wire _38942 = _38939 ^ _38941;
  wire _38943 = _38935 ^ _38942;
  wire _38944 = uncoded_block[1057] ^ uncoded_block[1061];
  wire _38945 = _38944 ^ _526;
  wire _38946 = _18359 ^ _530;
  wire _38947 = _38945 ^ _38946;
  wire _38948 = _21687 ^ _3696;
  wire _38949 = _38948 ^ _23070;
  wire _38950 = _38947 ^ _38949;
  wire _38951 = _10026 ^ _4444;
  wire _38952 = _38951 ^ _3709;
  wire _38953 = uncoded_block[1108] ^ uncoded_block[1112];
  wire _38954 = _38953 ^ _7133;
  wire _38955 = _1388 ^ _5854;
  wire _38956 = _38954 ^ _38955;
  wire _38957 = _38952 ^ _38956;
  wire _38958 = _38950 ^ _38957;
  wire _38959 = _38943 ^ _38958;
  wire _38960 = _23523 ^ _560;
  wire _38961 = _8345 ^ _35343;
  wire _38962 = _38960 ^ _38961;
  wire _38963 = uncoded_block[1144] ^ uncoded_block[1149];
  wire _38964 = uncoded_block[1150] ^ uncoded_block[1159];
  wire _38965 = _38963 ^ _38964;
  wire _38966 = _38965 ^ _10601;
  wire _38967 = _38962 ^ _38966;
  wire _38968 = _24449 ^ _27540;
  wire _38969 = _27545 ^ _6522;
  wire _38970 = uncoded_block[1193] ^ uncoded_block[1196];
  wire _38971 = _38970 ^ _11721;
  wire _38972 = _38969 ^ _38971;
  wire _38973 = _38968 ^ _38972;
  wire _38974 = _38967 ^ _38973;
  wire _38975 = _2982 ^ _10620;
  wire _38976 = _27551 ^ _38975;
  wire _38977 = _5894 ^ _2225;
  wire _38978 = _24005 ^ _38977;
  wire _38979 = _38976 ^ _38978;
  wire _38980 = _22651 ^ _5234;
  wire _38981 = _38179 ^ _38980;
  wire _38982 = _30781 ^ _38981;
  wire _38983 = _38979 ^ _38982;
  wire _38984 = _38974 ^ _38983;
  wire _38985 = _38959 ^ _38984;
  wire _38986 = _34163 ^ _2239;
  wire _38987 = _38986 ^ _22656;
  wire _38988 = _638 ^ _24023;
  wire _38989 = _12835 ^ _38988;
  wire _38990 = _38987 ^ _38989;
  wire _38991 = uncoded_block[1291] ^ uncoded_block[1294];
  wire _38992 = _4529 ^ _38991;
  wire _38993 = uncoded_block[1295] ^ uncoded_block[1297];
  wire _38994 = uncoded_block[1298] ^ uncoded_block[1302];
  wire _38995 = _38993 ^ _38994;
  wire _38996 = _38992 ^ _38995;
  wire _38997 = _22665 ^ _3807;
  wire _38998 = _3808 ^ _21748;
  wire _38999 = _38997 ^ _38998;
  wire _39000 = _38996 ^ _38999;
  wire _39001 = _38990 ^ _39000;
  wire _39002 = _15951 ^ _32513;
  wire _39003 = uncoded_block[1332] ^ uncoded_block[1338];
  wire _39004 = _39003 ^ _1497;
  wire _39005 = _39002 ^ _39004;
  wire _39006 = _7815 ^ _1498;
  wire _39007 = _5268 ^ _18436;
  wire _39008 = _39006 ^ _39007;
  wire _39009 = _39005 ^ _39008;
  wire _39010 = _10097 ^ _5273;
  wire _39011 = _679 ^ _3052;
  wire _39012 = _39010 ^ _39011;
  wire _39013 = _24954 ^ _3055;
  wire _39014 = _7219 ^ _19861;
  wire _39015 = _39013 ^ _39014;
  wire _39016 = _39012 ^ _39015;
  wire _39017 = _39009 ^ _39016;
  wire _39018 = _39001 ^ _39017;
  wire _39019 = _5950 ^ _7828;
  wire _39020 = _39019 ^ _7226;
  wire _39021 = _9585 ^ _7229;
  wire _39022 = _14969 ^ _39021;
  wire _39023 = _39020 ^ _39022;
  wire _39024 = _10120 ^ _3074;
  wire _39025 = _706 ^ _39024;
  wire _39026 = _14978 ^ _2318;
  wire _39027 = _1532 ^ _39026;
  wire _39028 = _39025 ^ _39027;
  wire _39029 = _39023 ^ _39028;
  wire _39030 = _4590 ^ _6619;
  wire _39031 = _16970 ^ _12335;
  wire _39032 = _39030 ^ _39031;
  wire _39033 = _2336 ^ _9602;
  wire _39034 = uncoded_block[1474] ^ uncoded_block[1483];
  wire _39035 = _35423 ^ _39034;
  wire _39036 = _39033 ^ _39035;
  wire _39037 = _39032 ^ _39036;
  wire _39038 = _17980 ^ _17489;
  wire _39039 = _13967 ^ _743;
  wire _39040 = _39038 ^ _39039;
  wire _39041 = uncoded_block[1506] ^ uncoded_block[1511];
  wire _39042 = _7259 ^ _39041;
  wire _39043 = _36650 ^ _39042;
  wire _39044 = _39040 ^ _39043;
  wire _39045 = _39037 ^ _39044;
  wire _39046 = _39029 ^ _39045;
  wire _39047 = _39018 ^ _39046;
  wire _39048 = _38985 ^ _39047;
  wire _39049 = _9053 ^ _9055;
  wire _39050 = uncoded_block[1533] ^ uncoded_block[1536];
  wire _39051 = _5999 ^ _39050;
  wire _39052 = _39049 ^ _39051;
  wire _39053 = _2365 ^ _1589;
  wire _39054 = _39053 ^ _23202;
  wire _39055 = _39052 ^ _39054;
  wire _39056 = _1597 ^ _11283;
  wire _39057 = _39056 ^ _3142;
  wire _39058 = _782 ^ _10171;
  wire _39059 = _39058 ^ _25455;
  wire _39060 = _39057 ^ _39059;
  wire _39061 = _39055 ^ _39060;
  wire _39062 = uncoded_block[1594] ^ uncoded_block[1597];
  wire _39063 = _39062 ^ _11847;
  wire _39064 = _798 ^ _10742;
  wire _39065 = _39063 ^ _39064;
  wire _39066 = _29997 ^ _12376;
  wire _39067 = _27210 ^ _39066;
  wire _39068 = _39065 ^ _39067;
  wire _39069 = _8508 ^ _23657;
  wire _39070 = _9099 ^ _7308;
  wire _39071 = _17527 ^ _12387;
  wire _39072 = _39070 ^ _39071;
  wire _39073 = _39069 ^ _39072;
  wire _39074 = _39068 ^ _39073;
  wire _39075 = _39061 ^ _39074;
  wire _39076 = _14011 ^ _12390;
  wire _39077 = _6055 ^ _3179;
  wire _39078 = _39076 ^ _39077;
  wire _39079 = _5399 ^ _19939;
  wire _39080 = _33862 ^ _9113;
  wire _39081 = _39079 ^ _39080;
  wire _39082 = _39078 ^ _39081;
  wire _39083 = uncoded_block[1683] ^ uncoded_block[1690];
  wire _39084 = _39083 ^ _3968;
  wire _39085 = _9677 ^ _25037;
  wire _39086 = _39084 ^ _39085;
  wire _39087 = _4700 ^ _16551;
  wire _39088 = _39087 ^ _30905;
  wire _39089 = _39086 ^ _39088;
  wire _39090 = _39082 ^ _39089;
  wire _39091 = _2441 ^ _17553;
  wire _39092 = _39091 ^ uncoded_block[1721];
  wire _39093 = _39090 ^ _39092;
  wire _39094 = _39075 ^ _39093;
  wire _39095 = _39048 ^ _39094;
  wire _39096 = _38928 ^ _39095;
  wire _39097 = _29176 ^ _33453;
  wire _39098 = _3998 ^ _14563;
  wire _39099 = _9694 ^ _6093;
  wire _39100 = _39098 ^ _39099;
  wire _39101 = _39097 ^ _39100;
  wire _39102 = _11 ^ _22333;
  wire _39103 = _3230 ^ _26850;
  wire _39104 = _39102 ^ _39103;
  wire _39105 = _1699 ^ _7969;
  wire _39106 = _31 ^ _6744;
  wire _39107 = _39105 ^ _39106;
  wire _39108 = _39104 ^ _39107;
  wire _39109 = _39101 ^ _39108;
  wire _39110 = _7367 ^ _5443;
  wire _39111 = _25955 ^ _41;
  wire _39112 = _39110 ^ _39111;
  wire _39113 = _14586 ^ _6755;
  wire _39114 = _6757 ^ _14068;
  wire _39115 = _39113 ^ _39114;
  wire _39116 = _39112 ^ _39115;
  wire _39117 = _7986 ^ _4034;
  wire _39118 = _4746 ^ _39117;
  wire _39119 = _7990 ^ _4750;
  wire _39120 = _39119 ^ _38722;
  wire _39121 = _39118 ^ _39120;
  wire _39122 = _39116 ^ _39121;
  wire _39123 = _39109 ^ _39122;
  wire _39124 = _923 ^ _21898;
  wire _39125 = _22819 ^ _3265;
  wire _39126 = _39124 ^ _39125;
  wire _39127 = _6780 ^ _1744;
  wire _39128 = uncoded_block[161] ^ uncoded_block[164];
  wire _39129 = _71 ^ _39128;
  wire _39130 = _39127 ^ _39129;
  wire _39131 = _39126 ^ _39130;
  wire _39132 = _8589 ^ _5473;
  wire _39133 = _938 ^ _1756;
  wire _39134 = _39132 ^ _39133;
  wire _39135 = _940 ^ _5477;
  wire _39136 = _18111 ^ _6155;
  wire _39137 = _39135 ^ _39136;
  wire _39138 = _39134 ^ _39137;
  wire _39139 = _39131 ^ _39138;
  wire _39140 = _2532 ^ _10849;
  wire _39141 = _3289 ^ _4070;
  wire _39142 = _39140 ^ _39141;
  wire _39143 = _956 ^ _959;
  wire _39144 = _14102 ^ _39143;
  wire _39145 = _39142 ^ _39144;
  wire _39146 = _10854 ^ _3299;
  wire _39147 = _21461 ^ _39146;
  wire _39148 = _4082 ^ _28051;
  wire _39149 = _39147 ^ _39148;
  wire _39150 = _39145 ^ _39149;
  wire _39151 = _39139 ^ _39150;
  wire _39152 = _39123 ^ _39151;
  wire _39153 = _2552 ^ _4797;
  wire _39154 = uncoded_block[249] ^ uncoded_block[252];
  wire _39155 = _8616 ^ _39154;
  wire _39156 = _39153 ^ _39155;
  wire _39157 = _1786 ^ _1788;
  wire _39158 = _4096 ^ _20523;
  wire _39159 = _39157 ^ _39158;
  wire _39160 = _39156 ^ _39159;
  wire _39161 = _985 ^ _6192;
  wire _39162 = _4814 ^ _988;
  wire _39163 = _39161 ^ _39162;
  wire _39164 = _8632 ^ _13069;
  wire _39165 = _15665 ^ _2577;
  wire _39166 = _39164 ^ _39165;
  wire _39167 = _39163 ^ _39166;
  wire _39168 = _39160 ^ _39167;
  wire _39169 = _12515 ^ _3334;
  wire _39170 = uncoded_block[312] ^ uncoded_block[314];
  wire _39171 = _8056 ^ _39170;
  wire _39172 = _39169 ^ _39171;
  wire _39173 = _6209 ^ _11444;
  wire _39174 = _28461 ^ _39173;
  wire _39175 = _39172 ^ _39174;
  wire _39176 = _1017 ^ _1825;
  wire _39177 = uncoded_block[349] ^ uncoded_block[357];
  wire _39178 = _18621 ^ _39177;
  wire _39179 = _39176 ^ _39178;
  wire _39180 = _3365 ^ _21955;
  wire _39181 = _39180 ^ _28085;
  wire _39182 = _39179 ^ _39181;
  wire _39183 = _39175 ^ _39182;
  wire _39184 = _39168 ^ _39183;
  wire _39185 = _6233 ^ _6876;
  wire _39186 = _31005 ^ _6239;
  wire _39187 = _39185 ^ _39186;
  wire _39188 = _16671 ^ _1048;
  wire _39189 = uncoded_block[401] ^ uncoded_block[409];
  wire _39190 = _39189 ^ _191;
  wire _39191 = _39188 ^ _39190;
  wire _39192 = _39187 ^ _39191;
  wire _39193 = _1055 ^ _4161;
  wire _39194 = _4163 ^ _8671;
  wire _39195 = _39193 ^ _39194;
  wire _39196 = _32297 ^ _3405;
  wire _39197 = uncoded_block[453] ^ uncoded_block[456];
  wire _39198 = _27756 ^ _39197;
  wire _39199 = _39196 ^ _39198;
  wire _39200 = _39195 ^ _39199;
  wire _39201 = _39192 ^ _39200;
  wire _39202 = _213 ^ _8681;
  wire _39203 = _9827 ^ _3416;
  wire _39204 = _39202 ^ _39203;
  wire _39205 = _4186 ^ _221;
  wire _39206 = _39205 ^ _19129;
  wire _39207 = _39204 ^ _39206;
  wire _39208 = _5598 ^ _13135;
  wire _39209 = _9832 ^ _1093;
  wire _39210 = _39208 ^ _39209;
  wire _39211 = _2668 ^ _5607;
  wire _39212 = _18200 ^ _39211;
  wire _39213 = _39210 ^ _39212;
  wire _39214 = _39207 ^ _39213;
  wire _39215 = _39201 ^ _39214;
  wire _39216 = _39184 ^ _39215;
  wire _39217 = _39152 ^ _39216;
  wire _39218 = _18203 ^ _26511;
  wire _39219 = _18206 ^ _9301;
  wire _39220 = _6929 ^ _9309;
  wire _39221 = _39219 ^ _39220;
  wire _39222 = _39218 ^ _39221;
  wire _39223 = _10957 ^ _23375;
  wire _39224 = _3468 ^ _13698;
  wire _39225 = _22005 ^ _39224;
  wire _39226 = _39223 ^ _39225;
  wire _39227 = _39222 ^ _39226;
  wire _39228 = _8732 ^ _28513;
  wire _39229 = _22012 ^ _1938;
  wire _39230 = _39229 ^ _34809;
  wire _39231 = _39228 ^ _39230;
  wire _39232 = uncoded_block[601] ^ uncoded_block[606];
  wire _39233 = uncoded_block[607] ^ uncoded_block[612];
  wire _39234 = _39232 ^ _39233;
  wire _39235 = _1149 ^ _281;
  wire _39236 = _39234 ^ _39235;
  wire _39237 = _6966 ^ _12071;
  wire _39238 = _29737 ^ _39237;
  wire _39239 = _39236 ^ _39238;
  wire _39240 = _39231 ^ _39239;
  wire _39241 = _39227 ^ _39240;
  wire _39242 = _3501 ^ _10984;
  wire _39243 = uncoded_block[642] ^ uncoded_block[646];
  wire _39244 = _39243 ^ _16247;
  wire _39245 = _39242 ^ _39244;
  wire _39246 = _302 ^ _3513;
  wire _39247 = _39246 ^ _13730;
  wire _39248 = _39245 ^ _39247;
  wire _39249 = _6349 ^ _319;
  wire _39250 = uncoded_block[688] ^ uncoded_block[691];
  wire _39251 = _5678 ^ _39250;
  wire _39252 = _39249 ^ _39251;
  wire _39253 = _30642 ^ _35245;
  wire _39254 = _39252 ^ _39253;
  wire _39255 = _39248 ^ _39254;
  wire _39256 = _1194 ^ _21595;
  wire _39257 = _39256 ^ _10456;
  wire _39258 = _11006 ^ _3547;
  wire _39259 = _7605 ^ _13208;
  wire _39260 = _39258 ^ _39259;
  wire _39261 = _39257 ^ _39260;
  wire _39262 = _13752 ^ _2002;
  wire _39263 = uncoded_block[763] ^ uncoded_block[773];
  wire _39264 = _5019 ^ _39263;
  wire _39265 = _39262 ^ _39264;
  wire _39266 = _14793 ^ _8790;
  wire _39267 = _14279 ^ _39266;
  wire _39268 = _39265 ^ _39267;
  wire _39269 = _39261 ^ _39268;
  wire _39270 = _39255 ^ _39269;
  wire _39271 = _39241 ^ _39270;
  wire _39272 = _2019 ^ _2799;
  wire _39273 = _6391 ^ _7628;
  wire _39274 = _39272 ^ _39273;
  wire _39275 = _24345 ^ _1238;
  wire _39276 = _39275 ^ _12681;
  wire _39277 = _39274 ^ _39276;
  wire _39278 = _12685 ^ _17794;
  wire _39279 = _9402 ^ _7043;
  wire _39280 = _2036 ^ _8808;
  wire _39281 = _39279 ^ _39280;
  wire _39282 = _39278 ^ _39281;
  wire _39283 = _39277 ^ _39282;
  wire _39284 = _13238 ^ _2046;
  wire _39285 = uncoded_block[856] ^ uncoded_block[859];
  wire _39286 = _39285 ^ _2824;
  wire _39287 = _39284 ^ _39286;
  wire _39288 = _2827 ^ _13791;
  wire _39289 = _39288 ^ _27455;
  wire _39290 = _39287 ^ _39289;
  wire _39291 = _5079 ^ _9416;
  wire _39292 = _428 ^ _1280;
  wire _39293 = _39291 ^ _39292;
  wire _39294 = uncoded_block[905] ^ uncoded_block[910];
  wire _39295 = _39294 ^ _435;
  wire _39296 = _39295 ^ _23025;
  wire _39297 = _39293 ^ _39296;
  wire _39298 = _39290 ^ _39297;
  wire _39299 = _39283 ^ _39298;
  wire _39300 = _31995 ^ _2857;
  wire _39301 = _39300 ^ _27055;
  wire _39302 = _7673 ^ _19747;
  wire _39303 = _12725 ^ _8274;
  wire _39304 = _39302 ^ _39303;
  wire _39305 = _39301 ^ _39304;
  wire _39306 = uncoded_block[961] ^ uncoded_block[966];
  wire _39307 = _9437 ^ _39306;
  wire _39308 = _7088 ^ _2877;
  wire _39309 = _39307 ^ _39308;
  wire _39310 = uncoded_block[979] ^ uncoded_block[985];
  wire _39311 = _39310 ^ _16338;
  wire _39312 = _28598 ^ _39311;
  wire _39313 = _39309 ^ _39312;
  wire _39314 = _39305 ^ _39313;
  wire _39315 = _1323 ^ _479;
  wire _39316 = _6457 ^ _2112;
  wire _39317 = _39315 ^ _39316;
  wire _39318 = _2114 ^ _15860;
  wire _39319 = _5131 ^ _8871;
  wire _39320 = _39318 ^ _39319;
  wire _39321 = _39317 ^ _39320;
  wire _39322 = _8872 ^ _36938;
  wire _39323 = uncoded_block[1035] ^ uncoded_block[1042];
  wire _39324 = _499 ^ _39323;
  wire _39325 = _39322 ^ _39324;
  wire _39326 = _2133 ^ _515;
  wire _39327 = _2914 ^ _11120;
  wire _39328 = _39326 ^ _39327;
  wire _39329 = _39325 ^ _39328;
  wire _39330 = _39321 ^ _39329;
  wire _39331 = _39314 ^ _39330;
  wire _39332 = _39299 ^ _39331;
  wire _39333 = _39271 ^ _39332;
  wire _39334 = _39217 ^ _39333;
  wire _39335 = _10569 ^ _1366;
  wire _39336 = _2146 ^ _7724;
  wire _39337 = _39335 ^ _39336;
  wire _39338 = uncoded_block[1090] ^ uncoded_block[1095];
  wire _39339 = _1374 ^ _39338;
  wire _39340 = _22607 ^ _39339;
  wire _39341 = _39337 ^ _39340;
  wire _39342 = _5843 ^ _15405;
  wire _39343 = _4450 ^ _13322;
  wire _39344 = _39342 ^ _39343;
  wire _39345 = _10587 ^ _12789;
  wire _39346 = _558 ^ _1393;
  wire _39347 = _39345 ^ _39346;
  wire _39348 = _39344 ^ _39347;
  wire _39349 = _39341 ^ _39348;
  wire _39350 = _23084 ^ _25333;
  wire _39351 = _8933 ^ _3727;
  wire _39352 = uncoded_block[1157] ^ uncoded_block[1165];
  wire _39353 = _39352 ^ _15907;
  wire _39354 = _39351 ^ _39353;
  wire _39355 = _39350 ^ _39354;
  wire _39356 = _17890 ^ _29887;
  wire _39357 = _8363 ^ _39356;
  wire _39358 = _15428 ^ _24910;
  wire _39359 = _21259 ^ _2206;
  wire _39360 = _39358 ^ _39359;
  wire _39361 = _39357 ^ _39360;
  wire _39362 = _39355 ^ _39361;
  wire _39363 = _39349 ^ _39362;
  wire _39364 = _7763 ^ _2210;
  wire _39365 = _7166 ^ _12813;
  wire _39366 = _39364 ^ _39365;
  wire _39367 = uncoded_block[1218] ^ uncoded_block[1226];
  wire _39368 = _605 ^ _39367;
  wire _39369 = _1440 ^ _2230;
  wire _39370 = _39368 ^ _39369;
  wire _39371 = _39366 ^ _39370;
  wire _39372 = _1451 ^ _8385;
  wire _39373 = _36991 ^ _39372;
  wire _39374 = uncoded_block[1260] ^ uncoded_block[1265];
  wire _39375 = _39374 ^ _3008;
  wire _39376 = _31657 ^ _39375;
  wire _39377 = _39373 ^ _39376;
  wire _39378 = _39371 ^ _39377;
  wire _39379 = uncoded_block[1271] ^ uncoded_block[1276];
  wire _39380 = uncoded_block[1277] ^ uncoded_block[1283];
  wire _39381 = _39379 ^ _39380;
  wire _39382 = uncoded_block[1293] ^ uncoded_block[1297];
  wire _39383 = _28317 ^ _39382;
  wire _39384 = _39381 ^ _39383;
  wire _39385 = _4532 ^ _8984;
  wire _39386 = _1472 ^ _1479;
  wire _39387 = _39385 ^ _39386;
  wire _39388 = _39384 ^ _39387;
  wire _39389 = _21748 ^ _15951;
  wire _39390 = _18878 ^ _39389;
  wire _39391 = uncoded_block[1330] ^ uncoded_block[1335];
  wire _39392 = _8411 ^ _39391;
  wire _39393 = uncoded_block[1338] ^ uncoded_block[1342];
  wire _39394 = _5259 ^ _39393;
  wire _39395 = _39392 ^ _39394;
  wire _39396 = _39390 ^ _39395;
  wire _39397 = _39388 ^ _39396;
  wire _39398 = _39378 ^ _39397;
  wire _39399 = _39363 ^ _39398;
  wire _39400 = _4556 ^ _11771;
  wire _39401 = _39400 ^ _28331;
  wire _39402 = _6587 ^ _5275;
  wire _39403 = _2284 ^ _8423;
  wire _39404 = _39402 ^ _39403;
  wire _39405 = _39401 ^ _39404;
  wire _39406 = uncoded_block[1374] ^ uncoded_block[1381];
  wire _39407 = _39406 ^ _19861;
  wire _39408 = _39407 ^ _37830;
  wire _39409 = _3841 ^ _8436;
  wire _39410 = uncoded_block[1415] ^ uncoded_block[1419];
  wire _39411 = _4580 ^ _39410;
  wire _39412 = _39409 ^ _39411;
  wire _39413 = _39408 ^ _39412;
  wire _39414 = _39405 ^ _39413;
  wire _39415 = _1526 ^ _3074;
  wire _39416 = _2308 ^ _14977;
  wire _39417 = _39415 ^ _39416;
  wire _39418 = _1541 ^ _3084;
  wire _39419 = _30405 ^ _39418;
  wire _39420 = _39417 ^ _39419;
  wire _39421 = _26763 ^ _11247;
  wire _39422 = _3088 ^ _3871;
  wire _39423 = _39421 ^ _39422;
  wire _39424 = _7247 ^ _733;
  wire _39425 = _39424 ^ _20864;
  wire _39426 = _39423 ^ _39425;
  wire _39427 = _39420 ^ _39426;
  wire _39428 = _39414 ^ _39427;
  wire _39429 = _3101 ^ _740;
  wire _39430 = _1565 ^ _11260;
  wire _39431 = _39429 ^ _39430;
  wire _39432 = _9618 ^ _7874;
  wire _39433 = _5334 ^ _13975;
  wire _39434 = _39432 ^ _39433;
  wire _39435 = _39431 ^ _39434;
  wire _39436 = _2357 ^ _755;
  wire _39437 = _5343 ^ _6002;
  wire _39438 = _39436 ^ _39437;
  wire _39439 = _16995 ^ _13472;
  wire _39440 = _6652 ^ _39439;
  wire _39441 = _39438 ^ _39440;
  wire _39442 = _39435 ^ _39441;
  wire _39443 = _6657 ^ _1596;
  wire _39444 = _774 ^ _16510;
  wire _39445 = _39443 ^ _39444;
  wire _39446 = _30870 ^ _24103;
  wire _39447 = _1609 ^ _2386;
  wire _39448 = _39446 ^ _39447;
  wire _39449 = _39445 ^ _39448;
  wire _39450 = uncoded_block[1592] ^ uncoded_block[1595];
  wire _39451 = _5368 ^ _39450;
  wire _39452 = _13486 ^ _3936;
  wire _39453 = _39451 ^ _39452;
  wire _39454 = _3153 ^ _800;
  wire _39455 = _3154 ^ _25905;
  wire _39456 = _39454 ^ _39455;
  wire _39457 = _39453 ^ _39456;
  wire _39458 = _39449 ^ _39457;
  wire _39459 = _39442 ^ _39458;
  wire _39460 = _39428 ^ _39459;
  wire _39461 = _39399 ^ _39460;
  wire _39462 = _808 ^ _5388;
  wire _39463 = _21833 ^ _39462;
  wire _39464 = _9659 ^ _3948;
  wire _39465 = uncoded_block[1648] ^ uncoded_block[1653];
  wire _39466 = _27651 ^ _39465;
  wire _39467 = _39464 ^ _39466;
  wire _39468 = _39463 ^ _39467;
  wire _39469 = _19471 ^ _3962;
  wire _39470 = _9110 ^ _39469;
  wire _39471 = _25029 ^ _39470;
  wire _39472 = _39468 ^ _39471;
  wire _39473 = _10202 ^ _3187;
  wire _39474 = _39473 ^ _21391;
  wire _39475 = _9675 ^ _1669;
  wire _39476 = _3973 ^ _3975;
  wire _39477 = _39475 ^ _39476;
  wire _39478 = _39474 ^ _39477;
  wire _39479 = _3976 ^ _852;
  wire _39480 = _33025 ^ _12976;
  wire _39481 = _39479 ^ _39480;
  wire _39482 = _39481 ^ uncoded_block[1722];
  wire _39483 = _39478 ^ _39482;
  wire _39484 = _39472 ^ _39483;
  wire _39485 = _39461 ^ _39484;
  wire _39486 = _39334 ^ _39485;
  wire _39487 = _1683 ^ _3;
  wire _39488 = _39487 ^ _7349;
  wire _39489 = _15075 ^ _5423;
  wire _39490 = _4716 ^ _19963;
  wire _39491 = _39489 ^ _39490;
  wire _39492 = _39488 ^ _39491;
  wire _39493 = _4001 ^ _17562;
  wire _39494 = _39493 ^ _22794;
  wire _39495 = _4008 ^ _7966;
  wire _39496 = _3233 ^ _4014;
  wire _39497 = _39495 ^ _39496;
  wire _39498 = _39494 ^ _39497;
  wire _39499 = _39492 ^ _39498;
  wire _39500 = _7969 ^ _7974;
  wire _39501 = _39500 ^ _3242;
  wire _39502 = _4020 ^ _14586;
  wire _39503 = _2484 ^ _8566;
  wire _39504 = _39502 ^ _39503;
  wire _39505 = _39501 ^ _39504;
  wire _39506 = _6115 ^ _14068;
  wire _39507 = _39506 ^ _17083;
  wire _39508 = _19520 ^ _16589;
  wire _39509 = _13571 ^ _20961;
  wire _39510 = _39508 ^ _39509;
  wire _39511 = _39507 ^ _39510;
  wire _39512 = _39505 ^ _39511;
  wire _39513 = _39499 ^ _39512;
  wire _39514 = _28448 ^ _33065;
  wire _39515 = _11918 ^ _2511;
  wire _39516 = _4046 ^ _1744;
  wire _39517 = _39515 ^ _39516;
  wire _39518 = _39514 ^ _39517;
  wire _39519 = _15623 ^ _7397;
  wire _39520 = _39519 ^ _15119;
  wire _39521 = _29208 ^ _5473;
  wire _39522 = _2521 ^ _6794;
  wire _39523 = _39521 ^ _39522;
  wire _39524 = _39520 ^ _39523;
  wire _39525 = _39518 ^ _39524;
  wire _39526 = _4062 ^ _2529;
  wire _39527 = _39526 ^ _4069;
  wire _39528 = _3289 ^ _8600;
  wire _39529 = uncoded_block[211] ^ uncoded_block[215];
  wire _39530 = _39529 ^ _1772;
  wire _39531 = _39528 ^ _39530;
  wire _39532 = _39527 ^ _39531;
  wire _39533 = _25990 ^ _16125;
  wire _39534 = _968 ^ _2552;
  wire _39535 = _39533 ^ _39534;
  wire _39536 = _8032 ^ _7432;
  wire _39537 = uncoded_block[251] ^ uncoded_block[256];
  wire _39538 = _39537 ^ _976;
  wire _39539 = _39536 ^ _39538;
  wire _39540 = _39535 ^ _39539;
  wire _39541 = _39532 ^ _39540;
  wire _39542 = _39525 ^ _39541;
  wire _39543 = _39513 ^ _39542;
  wire _39544 = _128 ^ _4814;
  wire _39545 = _25115 ^ _39544;
  wire _39546 = _11967 ^ _24212;
  wire _39547 = _5522 ^ _38762;
  wire _39548 = _39546 ^ _39547;
  wire _39549 = _39545 ^ _39548;
  wire _39550 = _995 ^ _137;
  wire _39551 = _39550 ^ _6203;
  wire _39552 = _143 ^ _21017;
  wire _39553 = _1003 ^ _3340;
  wire _39554 = _39552 ^ _39553;
  wire _39555 = _39551 ^ _39554;
  wire _39556 = _39549 ^ _39555;
  wire _39557 = _11439 ^ _29663;
  wire _39558 = _3347 ^ _1014;
  wire _39559 = _39557 ^ _39558;
  wire _39560 = uncoded_block[332] ^ uncoded_block[337];
  wire _39561 = _5534 ^ _39560;
  wire _39562 = _4840 ^ _2596;
  wire _39563 = _39561 ^ _39562;
  wire _39564 = _39559 ^ _39563;
  wire _39565 = _14662 ^ _1028;
  wire _39566 = _39565 ^ _3363;
  wire _39567 = uncoded_block[362] ^ uncoded_block[369];
  wire _39568 = _3365 ^ _39567;
  wire _39569 = _39568 ^ _35947;
  wire _39570 = _39566 ^ _39569;
  wire _39571 = _39564 ^ _39570;
  wire _39572 = _39556 ^ _39571;
  wire _39573 = _20056 ^ _1841;
  wire _39574 = _14677 ^ _19604;
  wire _39575 = _39573 ^ _39574;
  wire _39576 = _180 ^ _5559;
  wire _39577 = _12545 ^ _3391;
  wire _39578 = _39576 ^ _39577;
  wire _39579 = _39575 ^ _39578;
  wire _39580 = _28848 ^ _6888;
  wire _39581 = _17177 ^ _15704;
  wire _39582 = _9271 ^ _201;
  wire _39583 = _39581 ^ _39582;
  wire _39584 = _39580 ^ _39583;
  wire _39585 = _39579 ^ _39584;
  wire _39586 = uncoded_block[444] ^ uncoded_block[449];
  wire _39587 = _39586 ^ _209;
  wire _39588 = _5579 ^ _39587;
  wire _39589 = _1872 ^ _35196;
  wire _39590 = _39588 ^ _39589;
  wire _39591 = uncoded_block[468] ^ uncoded_block[477];
  wire _39592 = _39591 ^ _5592;
  wire _39593 = _4895 ^ _4897;
  wire _39594 = _39592 ^ _39593;
  wire _39595 = _13139 ^ _1097;
  wire _39596 = _29705 ^ _39595;
  wire _39597 = _39594 ^ _39596;
  wire _39598 = _39590 ^ _39597;
  wire _39599 = _39585 ^ _39598;
  wire _39600 = _39572 ^ _39599;
  wire _39601 = _39543 ^ _39600;
  wire _39602 = _7529 ^ _17694;
  wire _39603 = _3440 ^ _9841;
  wire _39604 = _39602 ^ _39603;
  wire _39605 = _1108 ^ _20099;
  wire _39606 = _39605 ^ _33588;
  wire _39607 = _39604 ^ _39606;
  wire _39608 = _14198 ^ _9854;
  wire _39609 = _39608 ^ _15235;
  wire _39610 = _247 ^ _3459;
  wire _39611 = uncoded_block[556] ^ uncoded_block[559];
  wire _39612 = _1122 ^ _39611;
  wire _39613 = _39610 ^ _39612;
  wire _39614 = _39609 ^ _39613;
  wire _39615 = _39607 ^ _39614;
  wire _39616 = _21555 ^ _7550;
  wire _39617 = uncoded_block[569] ^ uncoded_block[572];
  wire _39618 = _39617 ^ _262;
  wire _39619 = _39616 ^ _39618;
  wire _39620 = _6312 ^ _4947;
  wire _39621 = uncoded_block[591] ^ uncoded_block[596];
  wire _39622 = _1141 ^ _39621;
  wire _39623 = _39620 ^ _39622;
  wire _39624 = _39619 ^ _39623;
  wire _39625 = _7559 ^ _14219;
  wire _39626 = _4959 ^ _13713;
  wire _39627 = _4960 ^ _3499;
  wire _39628 = _39626 ^ _39627;
  wire _39629 = _39625 ^ _39628;
  wire _39630 = _39624 ^ _39629;
  wire _39631 = _39615 ^ _39630;
  wire _39632 = _4966 ^ _27803;
  wire _39633 = _10425 ^ _6341;
  wire _39634 = _28528 ^ _39633;
  wire _39635 = _39632 ^ _39634;
  wire _39636 = _16249 ^ _13726;
  wire _39637 = _9886 ^ _15775;
  wire _39638 = _39636 ^ _39637;
  wire _39639 = _21586 ^ _3526;
  wire _39640 = _18716 ^ _39250;
  wire _39641 = _39639 ^ _39640;
  wire _39642 = _39638 ^ _39641;
  wire _39643 = _39635 ^ _39642;
  wire _39644 = _3529 ^ _333;
  wire _39645 = _31519 ^ _39644;
  wire _39646 = uncoded_block[702] ^ uncoded_block[710];
  wire _39647 = _39646 ^ _4998;
  wire _39648 = _4999 ^ _5002;
  wire _39649 = _39647 ^ _39648;
  wire _39650 = _39645 ^ _39649;
  wire _39651 = uncoded_block[723] ^ uncoded_block[727];
  wire _39652 = _39651 ^ _30651;
  wire _39653 = _31087 ^ _39652;
  wire _39654 = _3549 ^ _13752;
  wire _39655 = _39654 ^ _2782;
  wire _39656 = _39653 ^ _39655;
  wire _39657 = _39650 ^ _39656;
  wire _39658 = _39643 ^ _39657;
  wire _39659 = _39631 ^ _39658;
  wire _39660 = _22514 ^ _38873;
  wire _39661 = uncoded_block[776] ^ uncoded_block[782];
  wire _39662 = _39661 ^ _4309;
  wire _39663 = _39662 ^ _27021;
  wire _39664 = _39660 ^ _39663;
  wire _39665 = _12126 ^ _8793;
  wire _39666 = _36474 ^ _39665;
  wire _39667 = _392 ^ _9397;
  wire _39668 = _12131 ^ _3588;
  wire _39669 = _39667 ^ _39668;
  wire _39670 = _39666 ^ _39669;
  wire _39671 = _39664 ^ _39670;
  wire _39672 = uncoded_block[828] ^ uncoded_block[835];
  wire _39673 = _39672 ^ _11043;
  wire _39674 = _39673 ^ _32395;
  wire _39675 = _4340 ^ _8809;
  wire _39676 = uncoded_block[858] ^ uncoded_block[862];
  wire _39677 = _7049 ^ _39676;
  wire _39678 = _39675 ^ _39677;
  wire _39679 = _39674 ^ _39678;
  wire _39680 = uncoded_block[865] ^ uncoded_block[870];
  wire _39681 = _9949 ^ _39680;
  wire _39682 = _1269 ^ _16815;
  wire _39683 = _39681 ^ _39682;
  wire _39684 = _2058 ^ _5083;
  wire _39685 = _5758 ^ _29809;
  wire _39686 = _39684 ^ _39685;
  wire _39687 = _39683 ^ _39686;
  wire _39688 = _39679 ^ _39687;
  wire _39689 = _39671 ^ _39688;
  wire _39690 = _3625 ^ _3628;
  wire _39691 = _16310 ^ _39690;
  wire _39692 = uncoded_block[920] ^ uncoded_block[922];
  wire _39693 = _3629 ^ _39692;
  wire _39694 = _39693 ^ _30698;
  wire _39695 = _39691 ^ _39694;
  wire _39696 = _2862 ^ _9971;
  wire _39697 = _456 ^ _14326;
  wire _39698 = _39696 ^ _39697;
  wire _39699 = _5779 ^ _461;
  wire _39700 = _39699 ^ _33267;
  wire _39701 = _39698 ^ _39700;
  wire _39702 = _39695 ^ _39701;
  wire _39703 = _1314 ^ _4390;
  wire _39704 = _38914 ^ _39703;
  wire _39705 = _8287 ^ _23938;
  wire _39706 = _38919 ^ _39705;
  wire _39707 = _39704 ^ _39706;
  wire _39708 = _28238 ^ _18335;
  wire _39709 = _8866 ^ _27077;
  wire _39710 = uncoded_block[1020] ^ uncoded_block[1025];
  wire _39711 = _8871 ^ _39710;
  wire _39712 = _39709 ^ _39711;
  wire _39713 = _39708 ^ _39712;
  wire _39714 = _39707 ^ _39713;
  wire _39715 = _39702 ^ _39714;
  wire _39716 = _39689 ^ _39715;
  wire _39717 = _39659 ^ _39716;
  wire _39718 = _39601 ^ _39717;
  wire _39719 = uncoded_block[1029] ^ uncoded_block[1034];
  wire _39720 = _39719 ^ _1342;
  wire _39721 = _5810 ^ _12208;
  wire _39722 = _39720 ^ _39721;
  wire _39723 = _515 ^ _14867;
  wire _39724 = _39723 ^ _5152;
  wire _39725 = _39722 ^ _39724;
  wire _39726 = _10566 ^ _14357;
  wire _39727 = _39726 ^ _26222;
  wire _39728 = _3692 ^ _3695;
  wire _39729 = _27515 ^ _5840;
  wire _39730 = _39728 ^ _39729;
  wire _39731 = _39727 ^ _39730;
  wire _39732 = _39725 ^ _39731;
  wire _39733 = _7129 ^ _543;
  wire _39734 = uncoded_block[1105] ^ uncoded_block[1109];
  wire _39735 = _7731 ^ _39734;
  wire _39736 = _39733 ^ _39735;
  wire _39737 = _7133 ^ _5175;
  wire _39738 = _12789 ^ _12791;
  wire _39739 = _39737 ^ _39738;
  wire _39740 = _39736 ^ _39739;
  wire _39741 = _9494 ^ _6501;
  wire _39742 = _39741 ^ _10594;
  wire _39743 = _25332 ^ _10597;
  wire _39744 = _39743 ^ _24900;
  wire _39745 = _39742 ^ _39744;
  wire _39746 = _39740 ^ _39745;
  wire _39747 = _39732 ^ _39746;
  wire _39748 = _11157 ^ _1404;
  wire _39749 = _39748 ^ _30339;
  wire _39750 = _2192 ^ _589;
  wire _39751 = _17888 ^ _39750;
  wire _39752 = _39749 ^ _39751;
  wire _39753 = uncoded_block[1185] ^ uncoded_block[1193];
  wire _39754 = _2195 ^ _39753;
  wire _39755 = _39754 ^ _28294;
  wire _39756 = _14912 ^ _10620;
  wire _39757 = _23541 ^ _39756;
  wire _39758 = _39755 ^ _39757;
  wire _39759 = _39752 ^ _39758;
  wire _39760 = _3766 ^ _5891;
  wire _39761 = _39760 ^ _8961;
  wire _39762 = _6536 ^ _18860;
  wire _39763 = _1449 ^ _8385;
  wire _39764 = _39762 ^ _39763;
  wire _39765 = _39761 ^ _39764;
  wire _39766 = uncoded_block[1255] ^ uncoded_block[1261];
  wire _39767 = _2235 ^ _39766;
  wire _39768 = _39767 ^ _24473;
  wire _39769 = uncoded_block[1267] ^ uncoded_block[1273];
  wire _39770 = _39769 ^ _9539;
  wire _39771 = _39770 ^ _3795;
  wire _39772 = _39768 ^ _39771;
  wire _39773 = _39765 ^ _39772;
  wire _39774 = _39759 ^ _39773;
  wire _39775 = _39747 ^ _39774;
  wire _39776 = _6557 ^ _24023;
  wire _39777 = _13380 ^ _38991;
  wire _39778 = _39776 ^ _39777;
  wire _39779 = _10647 ^ _646;
  wire _39780 = _3805 ^ _8991;
  wire _39781 = _39779 ^ _39780;
  wire _39782 = _39778 ^ _39781;
  wire _39783 = _8992 ^ _4539;
  wire _39784 = _39783 ^ _14944;
  wire _39785 = uncoded_block[1323] ^ uncoded_block[1336];
  wire _39786 = _39785 ^ _9563;
  wire _39787 = _2277 ^ _1498;
  wire _39788 = _39786 ^ _39787;
  wire _39789 = _39784 ^ _39788;
  wire _39790 = _39782 ^ _39789;
  wire _39791 = _5268 ^ _18434;
  wire _39792 = _5272 ^ _25393;
  wire _39793 = _39791 ^ _39792;
  wire _39794 = _10665 ^ _31686;
  wire _39795 = _39794 ^ _19390;
  wire _39796 = _39793 ^ _39795;
  wire _39797 = _32935 ^ _688;
  wire _39798 = _39797 ^ _23596;
  wire _39799 = _8432 ^ _2301;
  wire _39800 = _39798 ^ _39799;
  wire _39801 = _39796 ^ _39800;
  wire _39802 = _39790 ^ _39801;
  wire _39803 = _10118 ^ _13428;
  wire _39804 = _24515 ^ _39803;
  wire _39805 = uncoded_block[1426] ^ uncoded_block[1433];
  wire _39806 = _39805 ^ _3857;
  wire _39807 = _39806 ^ _32952;
  wire _39808 = _39804 ^ _39807;
  wire _39809 = _8450 ^ _3865;
  wire _39810 = _39809 ^ _18466;
  wire _39811 = _3089 ^ _2336;
  wire _39812 = _39811 ^ _9603;
  wire _39813 = _39810 ^ _39812;
  wire _39814 = _39808 ^ _39813;
  wire _39815 = _2344 ^ _5320;
  wire _39816 = _39815 ^ _17982;
  wire _39817 = _12344 ^ _4614;
  wire _39818 = _7259 ^ _19892;
  wire _39819 = _39817 ^ _39818;
  wire _39820 = _39816 ^ _39819;
  wire _39821 = _6643 ^ _12352;
  wire _39822 = _12904 ^ _39821;
  wire _39823 = uncoded_block[1526] ^ uncoded_block[1533];
  wire _39824 = _3118 ^ _39823;
  wire _39825 = _39824 ^ _21351;
  wire _39826 = _39822 ^ _39825;
  wire _39827 = _39820 ^ _39826;
  wire _39828 = _39814 ^ _39827;
  wire _39829 = _39802 ^ _39828;
  wire _39830 = _39775 ^ _39829;
  wire _39831 = _13471 ^ _767;
  wire _39832 = _32559 ^ _39831;
  wire _39833 = _9070 ^ _11281;
  wire _39834 = uncoded_block[1561] ^ uncoded_block[1567];
  wire _39835 = _1597 ^ _39834;
  wire _39836 = _39833 ^ _39835;
  wire _39837 = _39832 ^ _39836;
  wire _39838 = uncoded_block[1571] ^ uncoded_block[1579];
  wire _39839 = _7891 ^ _39838;
  wire _39840 = _5368 ^ _4653;
  wire _39841 = _39839 ^ _39840;
  wire _39842 = _791 ^ _4659;
  wire _39843 = _7902 ^ _801;
  wire _39844 = _39842 ^ _39843;
  wire _39845 = _39841 ^ _39844;
  wire _39846 = _39837 ^ _39845;
  wire _39847 = _6042 ^ _7297;
  wire _39848 = _7911 ^ _11853;
  wire _39849 = _39847 ^ _39848;
  wire _39850 = _4665 ^ _31749;
  wire _39851 = _7914 ^ _18513;
  wire _39852 = _39850 ^ _39851;
  wire _39853 = _39849 ^ _39852;
  wire _39854 = uncoded_block[1647] ^ uncoded_block[1651];
  wire _39855 = _2411 ^ _39854;
  wire _39856 = _18030 ^ _6055;
  wire _39857 = _39855 ^ _39856;
  wire _39858 = _1654 ^ _5399;
  wire _39859 = _7928 ^ _2423;
  wire _39860 = _39858 ^ _39859;
  wire _39861 = _39857 ^ _39860;
  wire _39862 = _39853 ^ _39861;
  wire _39863 = _39846 ^ _39862;
  wire _39864 = _3962 ^ _20427;
  wire _39865 = _7933 ^ _20429;
  wire _39866 = _39864 ^ _39865;
  wire _39867 = _9115 ^ _9118;
  wire _39868 = _8533 ^ _22314;
  wire _39869 = _39867 ^ _39868;
  wire _39870 = _39866 ^ _39869;
  wire _39871 = uncoded_block[1708] ^ uncoded_block[1712];
  wire _39872 = _2435 ^ _39871;
  wire _39873 = _1677 ^ uncoded_block[1719];
  wire _39874 = _39872 ^ _39873;
  wire _39875 = _39870 ^ _39874;
  wire _39876 = _39863 ^ _39875;
  wire _39877 = _39830 ^ _39876;
  wire _39878 = _39718 ^ _39877;
  wire _39879 = _17559 ^ _6086;
  wire _39880 = _37516 ^ _39879;
  wire _39881 = _871 ^ _5426;
  wire _39882 = _2459 ^ _15;
  wire _39883 = _39881 ^ _39882;
  wire _39884 = _39880 ^ _39883;
  wire _39885 = _14571 ^ _6099;
  wire _39886 = _1699 ^ _1703;
  wire _39887 = _39885 ^ _39886;
  wire _39888 = _9705 ^ _897;
  wire _39889 = _37526 ^ _39888;
  wire _39890 = _39887 ^ _39889;
  wire _39891 = _39884 ^ _39890;
  wire _39892 = _7979 ^ _17578;
  wire _39893 = _9713 ^ _19515;
  wire _39894 = _39892 ^ _39893;
  wire _39895 = _908 ^ _9718;
  wire _39896 = _38713 ^ _50;
  wire _39897 = _39895 ^ _39896;
  wire _39898 = _39894 ^ _39897;
  wire _39899 = uncoded_block[111] ^ uncoded_block[114];
  wire _39900 = _6123 ^ _39899;
  wire _39901 = _2495 ^ _2498;
  wire _39902 = _39900 ^ _39901;
  wire _39903 = uncoded_block[127] ^ uncoded_block[131];
  wire _39904 = _56 ^ _39903;
  wire _39905 = _924 ^ _926;
  wire _39906 = _39904 ^ _39905;
  wire _39907 = _39902 ^ _39906;
  wire _39908 = _39898 ^ _39907;
  wire _39909 = _39891 ^ _39908;
  wire _39910 = uncoded_block[138] ^ uncoded_block[141];
  wire _39911 = _1736 ^ _39910;
  wire _39912 = _15114 ^ _7392;
  wire _39913 = _39911 ^ _39912;
  wire _39914 = _14082 ^ _70;
  wire _39915 = _39914 ^ _37548;
  wire _39916 = _39913 ^ _39915;
  wire _39917 = _19042 ^ _6788;
  wire _39918 = _19535 ^ _39917;
  wire _39919 = uncoded_block[171] ^ uncoded_block[180];
  wire _39920 = _39919 ^ _28037;
  wire _39921 = uncoded_block[190] ^ uncoded_block[194];
  wire _39922 = _13588 ^ _39921;
  wire _39923 = _39920 ^ _39922;
  wire _39924 = _39918 ^ _39923;
  wire _39925 = _39916 ^ _39924;
  wire _39926 = _30961 ^ _26878;
  wire _39927 = _97 ^ _9750;
  wire _39928 = uncoded_block[218] ^ uncoded_block[224];
  wire _39929 = _39928 ^ _6168;
  wire _39930 = _39927 ^ _39929;
  wire _39931 = _39926 ^ _39930;
  wire _39932 = _1774 ^ _30087;
  wire _39933 = _5500 ^ _6172;
  wire _39934 = _39932 ^ _39933;
  wire _39935 = _35145 ^ _7432;
  wire _39936 = _39935 ^ _18597;
  wire _39937 = _39934 ^ _39936;
  wire _39938 = _39931 ^ _39937;
  wire _39939 = _39925 ^ _39938;
  wire _39940 = _39909 ^ _39939;
  wire _39941 = _6188 ^ _2566;
  wire _39942 = _13056 ^ _39941;
  wire _39943 = _18607 ^ _20529;
  wire _39944 = _39942 ^ _39943;
  wire _39945 = _31843 ^ _14133;
  wire _39946 = _31426 ^ _39945;
  wire _39947 = _14652 ^ _1002;
  wire _39948 = _3338 ^ _146;
  wire _39949 = _39947 ^ _39948;
  wire _39950 = _39946 ^ _39949;
  wire _39951 = _39944 ^ _39950;
  wire _39952 = _3347 ^ _30117;
  wire _39953 = _17150 ^ _39952;
  wire _39954 = _9235 ^ _4126;
  wire _39955 = _8065 ^ _9790;
  wire _39956 = _39954 ^ _39955;
  wire _39957 = _39953 ^ _39956;
  wire _39958 = _162 ^ _165;
  wire _39959 = _39958 ^ _28471;
  wire _39960 = _3369 ^ _16664;
  wire _39961 = uncoded_block[380] ^ uncoded_block[385];
  wire _39962 = _6233 ^ _39961;
  wire _39963 = _39960 ^ _39962;
  wire _39964 = _39959 ^ _39963;
  wire _39965 = _39957 ^ _39964;
  wire _39966 = _39951 ^ _39965;
  wire _39967 = _2613 ^ _2615;
  wire _39968 = _4152 ^ _2622;
  wire _39969 = _39967 ^ _39968;
  wire _39970 = _2623 ^ _34766;
  wire _39971 = _39970 ^ _9268;
  wire _39972 = _39969 ^ _39971;
  wire _39973 = _11477 ^ _8671;
  wire _39974 = _1062 ^ _13115;
  wire _39975 = _39973 ^ _39974;
  wire _39976 = uncoded_block[436] ^ uncoded_block[440];
  wire _39977 = _10352 ^ _39976;
  wire _39978 = _39977 ^ _207;
  wire _39979 = _39975 ^ _39978;
  wire _39980 = _39972 ^ _39979;
  wire _39981 = _10356 ^ _33565;
  wire _39982 = _1076 ^ _10926;
  wire _39983 = _39981 ^ _39982;
  wire _39984 = uncoded_block[467] ^ uncoded_block[473];
  wire _39985 = _11491 ^ _39984;
  wire _39986 = _11494 ^ _7513;
  wire _39987 = _39985 ^ _39986;
  wire _39988 = _39983 ^ _39987;
  wire _39989 = uncoded_block[482] ^ uncoded_block[486];
  wire _39990 = _39989 ^ _4194;
  wire _39991 = _3424 ^ _3432;
  wire _39992 = _39990 ^ _39991;
  wire _39993 = _34785 ^ _19135;
  wire _39994 = _1892 ^ _10376;
  wire _39995 = _39993 ^ _39994;
  wire _39996 = _39992 ^ _39995;
  wire _39997 = _39988 ^ _39996;
  wire _39998 = _39980 ^ _39997;
  wire _39999 = _39966 ^ _39998;
  wire _40000 = _39940 ^ _39999;
  wire _40001 = _10945 ^ _21992;
  wire _40002 = _1108 ^ _13684;
  wire _40003 = _40001 ^ _40002;
  wire _40004 = _1900 ^ _9850;
  wire _40005 = _40004 ^ _34800;
  wire _40006 = _40003 ^ _40005;
  wire _40007 = _244 ^ _6300;
  wire _40008 = uncoded_block[556] ^ uncoded_block[562];
  wire _40009 = _40008 ^ _32736;
  wire _40010 = _40007 ^ _40009;
  wire _40011 = uncoded_block[569] ^ uncoded_block[574];
  wire _40012 = _7550 ^ _40011;
  wire _40013 = _10967 ^ _24289;
  wire _40014 = _40012 ^ _40013;
  wire _40015 = _40010 ^ _40014;
  wire _40016 = _40006 ^ _40015;
  wire _40017 = _2706 ^ _5646;
  wire _40018 = _37645 ^ _40017;
  wire _40019 = _34017 ^ _37648;
  wire _40020 = _40018 ^ _40019;
  wire _40021 = _14744 ^ _30196;
  wire _40022 = _29318 ^ _5661;
  wire _40023 = uncoded_block[642] ^ uncoded_block[645];
  wire _40024 = _4255 ^ _40023;
  wire _40025 = _40022 ^ _40024;
  wire _40026 = _40021 ^ _40025;
  wire _40027 = _40020 ^ _40026;
  wire _40028 = _40016 ^ _40027;
  wire _40029 = _2730 ^ _6341;
  wire _40030 = uncoded_block[655] ^ uncoded_block[658];
  wire _40031 = _4975 ^ _40030;
  wire _40032 = _40029 ^ _40031;
  wire _40033 = _4261 ^ _15270;
  wire _40034 = _309 ^ _15775;
  wire _40035 = _40033 ^ _40034;
  wire _40036 = _40032 ^ _40035;
  wire _40037 = _10434 ^ _3521;
  wire _40038 = _40037 ^ _24773;
  wire _40039 = _1186 ^ _328;
  wire _40040 = _15777 ^ _40039;
  wire _40041 = _40038 ^ _40040;
  wire _40042 = _40036 ^ _40041;
  wire _40043 = _19195 ^ _19197;
  wire _40044 = uncoded_block[711] ^ uncoded_block[715];
  wire _40045 = _15783 ^ _40044;
  wire _40046 = _40043 ^ _40045;
  wire _40047 = _13745 ^ _24324;
  wire _40048 = _40046 ^ _40047;
  wire _40049 = _2768 ^ _37283;
  wire _40050 = _11572 ^ _40049;
  wire _40051 = _34048 ^ _3550;
  wire _40052 = _40051 ^ _20158;
  wire _40053 = _40050 ^ _40052;
  wire _40054 = _40048 ^ _40053;
  wire _40055 = _40042 ^ _40054;
  wire _40056 = _40028 ^ _40055;
  wire _40057 = _4301 ^ _33217;
  wire _40058 = _10467 ^ _40057;
  wire _40059 = _13766 ^ _17284;
  wire _40060 = _2015 ^ _8215;
  wire _40061 = _40059 ^ _40060;
  wire _40062 = _40058 ^ _40061;
  wire _40063 = _5033 ^ _8791;
  wire _40064 = _19223 ^ _4317;
  wire _40065 = _40063 ^ _40064;
  wire _40066 = _9394 ^ _15814;
  wire _40067 = _11596 ^ _10485;
  wire _40068 = _40066 ^ _40067;
  wire _40069 = _40065 ^ _40068;
  wire _40070 = _40062 ^ _40069;
  wire _40071 = uncoded_block[823] ^ uncoded_block[827];
  wire _40072 = _32388 ^ _40071;
  wire _40073 = _40072 ^ _11041;
  wire _40074 = _35668 ^ _2036;
  wire _40075 = _20188 ^ _6406;
  wire _40076 = _40074 ^ _40075;
  wire _40077 = _40073 ^ _40076;
  wire _40078 = _8237 ^ _3600;
  wire _40079 = _14300 ^ _3603;
  wire _40080 = _40078 ^ _40079;
  wire _40081 = _5749 ^ _1269;
  wire _40082 = _11620 ^ _31131;
  wire _40083 = _40081 ^ _40082;
  wire _40084 = _40080 ^ _40083;
  wire _40085 = _40077 ^ _40084;
  wire _40086 = _40070 ^ _40085;
  wire _40087 = uncoded_block[888] ^ uncoded_block[893];
  wire _40088 = _14821 ^ _40087;
  wire _40089 = _5758 ^ _8827;
  wire _40090 = _40088 ^ _40089;
  wire _40091 = _6428 ^ _1287;
  wire _40092 = _40091 ^ _37723;
  wire _40093 = _40090 ^ _40092;
  wire _40094 = _15841 ^ _1296;
  wire _40095 = _40094 ^ _19258;
  wire _40096 = _7080 ^ _2863;
  wire _40097 = uncoded_block[944] ^ uncoded_block[951];
  wire _40098 = _40097 ^ _14329;
  wire _40099 = _40096 ^ _40098;
  wire _40100 = _40095 ^ _40099;
  wire _40101 = _40093 ^ _40100;
  wire _40102 = uncoded_block[967] ^ uncoded_block[975];
  wire _40103 = _40102 ^ _5114;
  wire _40104 = _32006 ^ _40103;
  wire _40105 = _36518 ^ _8855;
  wire _40106 = _1317 ^ _8859;
  wire _40107 = _40105 ^ _40106;
  wire _40108 = _40104 ^ _40107;
  wire _40109 = uncoded_block[1001] ^ uncoded_block[1005];
  wire _40110 = _28241 ^ _40109;
  wire _40111 = _28238 ^ _40110;
  wire _40112 = _4410 ^ _2891;
  wire _40113 = uncoded_block[1024] ^ uncoded_block[1029];
  wire _40114 = _1333 ^ _40113;
  wire _40115 = _40112 ^ _40114;
  wire _40116 = _40111 ^ _40115;
  wire _40117 = _40108 ^ _40116;
  wire _40118 = _40101 ^ _40117;
  wire _40119 = _40086 ^ _40118;
  wire _40120 = _40056 ^ _40119;
  wire _40121 = _40000 ^ _40120;
  wire _40122 = _5806 ^ _22595;
  wire _40123 = _40122 ^ _1347;
  wire _40124 = uncoded_block[1044] ^ uncoded_block[1049];
  wire _40125 = _512 ^ _40124;
  wire _40126 = _9464 ^ _1360;
  wire _40127 = _40125 ^ _40126;
  wire _40128 = _40123 ^ _40127;
  wire _40129 = _6483 ^ _5825;
  wire _40130 = _3685 ^ _526;
  wire _40131 = _40129 ^ _40130;
  wire _40132 = _32035 ^ _5834;
  wire _40133 = _40132 ^ _34126;
  wire _40134 = _40131 ^ _40133;
  wire _40135 = _40128 ^ _40134;
  wire _40136 = _20253 ^ _11689;
  wire _40137 = _40136 ^ _24428;
  wire _40138 = _13318 ^ _2164;
  wire _40139 = _12782 ^ _5175;
  wire _40140 = _40138 ^ _40139;
  wire _40141 = _40137 ^ _40140;
  wire _40142 = _2944 ^ _19322;
  wire _40143 = _25328 ^ _40142;
  wire _40144 = _5859 ^ _5861;
  wire _40145 = _15419 ^ _40144;
  wire _40146 = _40143 ^ _40145;
  wire _40147 = _40141 ^ _40146;
  wire _40148 = _40135 ^ _40147;
  wire _40149 = _2185 ^ _3727;
  wire _40150 = _14892 ^ _40149;
  wire _40151 = _3728 ^ _2188;
  wire _40152 = _7151 ^ _9506;
  wire _40153 = _40151 ^ _40152;
  wire _40154 = _40150 ^ _40153;
  wire _40155 = _14901 ^ _3740;
  wire _40156 = _13882 ^ _35749;
  wire _40157 = _40155 ^ _40156;
  wire _40158 = _24910 ^ _7758;
  wire _40159 = _2209 ^ _10617;
  wire _40160 = _40158 ^ _40159;
  wire _40161 = _40157 ^ _40160;
  wire _40162 = _40154 ^ _40161;
  wire _40163 = _12813 ^ _14914;
  wire _40164 = _29045 ^ _12819;
  wire _40165 = _40163 ^ _40164;
  wire _40166 = uncoded_block[1230] ^ uncoded_block[1233];
  wire _40167 = _40166 ^ _3771;
  wire _40168 = _19827 ^ _10627;
  wire _40169 = _40167 ^ _40168;
  wire _40170 = _40165 ^ _40169;
  wire _40171 = _19829 ^ _4511;
  wire _40172 = _5231 ^ _6546;
  wire _40173 = _40171 ^ _40172;
  wire _40174 = _13902 ^ _8392;
  wire _40175 = _40173 ^ _40174;
  wire _40176 = _40170 ^ _40175;
  wire _40177 = _40162 ^ _40176;
  wire _40178 = _40148 ^ _40177;
  wire _40179 = _2246 ^ _7793;
  wire _40180 = _24931 ^ _37808;
  wire _40181 = _40179 ^ _40180;
  wire _40182 = _641 ^ _10646;
  wire _40183 = _4531 ^ _8984;
  wire _40184 = _40182 ^ _40183;
  wire _40185 = _3805 ^ _1479;
  wire _40186 = _6572 ^ _21293;
  wire _40187 = _40185 ^ _40186;
  wire _40188 = _40184 ^ _40187;
  wire _40189 = _40181 ^ _40188;
  wire _40190 = uncoded_block[1321] ^ uncoded_block[1325];
  wire _40191 = _40190 ^ _8997;
  wire _40192 = _40191 ^ _37817;
  wire _40193 = _669 ^ _32518;
  wire _40194 = _37818 ^ _40193;
  wire _40195 = _40192 ^ _40194;
  wire _40196 = _12857 ^ _5940;
  wire _40197 = _6588 ^ _1504;
  wire _40198 = _40196 ^ _40197;
  wire _40199 = _11224 ^ _10668;
  wire _40200 = _2289 ^ _5285;
  wire _40201 = _40199 ^ _40200;
  wire _40202 = _40198 ^ _40201;
  wire _40203 = _40195 ^ _40202;
  wire _40204 = _40189 ^ _40203;
  wire _40205 = _691 ^ _694;
  wire _40206 = _32112 ^ _40205;
  wire _40207 = _13938 ^ _3066;
  wire _40208 = _40207 ^ _29501;
  wire _40209 = _40206 ^ _40208;
  wire _40210 = _5958 ^ _706;
  wire _40211 = _10120 ^ _3853;
  wire _40212 = _2311 ^ _5968;
  wire _40213 = _40211 ^ _40212;
  wire _40214 = _40210 ^ _40213;
  wire _40215 = _40209 ^ _40214;
  wire _40216 = _1533 ^ _2314;
  wire _40217 = _40216 ^ _33384;
  wire _40218 = _9597 ^ _1544;
  wire _40219 = _40218 ^ _25869;
  wire _40220 = _40217 ^ _40219;
  wire _40221 = _24528 ^ _5983;
  wire _40222 = _40221 ^ _37848;
  wire _40223 = uncoded_block[1483] ^ uncoded_block[1489];
  wire _40224 = _2344 ^ _40223;
  wire _40225 = _40224 ^ _17490;
  wire _40226 = _40222 ^ _40225;
  wire _40227 = _40220 ^ _40226;
  wire _40228 = _40215 ^ _40227;
  wire _40229 = _40204 ^ _40228;
  wire _40230 = _40178 ^ _40229;
  wire _40231 = _7257 ^ _30421;
  wire _40232 = _5334 ^ _19897;
  wire _40233 = _40232 ^ _10720;
  wire _40234 = _40231 ^ _40233;
  wire _40235 = _15010 ^ _23201;
  wire _40236 = _4638 ^ _774;
  wire _40237 = _37864 ^ _40236;
  wire _40238 = _40235 ^ _40237;
  wire _40239 = _40234 ^ _40238;
  wire _40240 = _2376 ^ _16510;
  wire _40241 = _21361 ^ _18952;
  wire _40242 = _40240 ^ _40241;
  wire _40243 = uncoded_block[1583] ^ uncoded_block[1587];
  wire _40244 = _40243 ^ _14512;
  wire _40245 = _792 ^ _3934;
  wire _40246 = _40244 ^ _40245;
  wire _40247 = _40242 ^ _40246;
  wire _40248 = _6039 ^ _3153;
  wire _40249 = _4662 ^ _6679;
  wire _40250 = _40248 ^ _40249;
  wire _40251 = _24115 ^ _6684;
  wire _40252 = _40251 ^ _35461;
  wire _40253 = _40250 ^ _40252;
  wire _40254 = _40247 ^ _40253;
  wire _40255 = _40239 ^ _40254;
  wire _40256 = _812 ^ _2405;
  wire _40257 = uncoded_block[1637] ^ uncoded_block[1648];
  wire _40258 = _40257 ^ _24578;
  wire _40259 = _40256 ^ _40258;
  wire _40260 = _14011 ^ _13508;
  wire _40261 = _4680 ^ _823;
  wire _40262 = _40260 ^ _40261;
  wire _40263 = _40259 ^ _40262;
  wire _40264 = _22761 ^ _5399;
  wire _40265 = _3183 ^ _13517;
  wire _40266 = _40264 ^ _40265;
  wire _40267 = _3187 ^ _13519;
  wire _40268 = _8527 ^ _6068;
  wire _40269 = _40267 ^ _40268;
  wire _40270 = _40266 ^ _40269;
  wire _40271 = _40263 ^ _40270;
  wire _40272 = _15063 ^ _7335;
  wire _40273 = _40272 ^ _29581;
  wire _40274 = _14552 ^ _17553;
  wire _40275 = _40274 ^ uncoded_block[1721];
  wire _40276 = _40273 ^ _40275;
  wire _40277 = _40271 ^ _40276;
  wire _40278 = _40255 ^ _40277;
  wire _40279 = _40230 ^ _40278;
  wire _40280 = _40121 ^ _40279;
  wire _40281 = _3209 ^ _1683;
  wire _40282 = _1684 ^ _4713;
  wire _40283 = _40281 ^ _40282;
  wire _40284 = _868 ^ _6087;
  wire _40285 = _40284 ^ _32205;
  wire _40286 = _40283 ^ _40285;
  wire _40287 = uncoded_block[37] ^ uncoded_block[44];
  wire _40288 = _13543 ^ _40287;
  wire _40289 = _39099 ^ _40288;
  wire _40290 = _885 ^ _3233;
  wire _40291 = _14575 ^ _888;
  wire _40292 = _40290 ^ _40291;
  wire _40293 = _40289 ^ _40292;
  wire _40294 = _40286 ^ _40293;
  wire _40295 = _10806 ^ _2475;
  wire _40296 = _25506 ^ _40295;
  wire _40297 = uncoded_block[73] ^ uncoded_block[80];
  wire _40298 = _6745 ^ _40297;
  wire _40299 = _35111 ^ _4738;
  wire _40300 = _40298 ^ _40299;
  wire _40301 = _40296 ^ _40300;
  wire _40302 = _19515 ^ _4026;
  wire _40303 = _11909 ^ _4028;
  wire _40304 = _40302 ^ _40303;
  wire _40305 = uncoded_block[103] ^ uncoded_block[107];
  wire _40306 = _40305 ^ _2491;
  wire _40307 = _5453 ^ _25521;
  wire _40308 = _40306 ^ _40307;
  wire _40309 = _40304 ^ _40308;
  wire _40310 = _40301 ^ _40309;
  wire _40311 = _40294 ^ _40310;
  wire _40312 = uncoded_block[119] ^ uncoded_block[124];
  wire _40313 = _40312 ^ _1730;
  wire _40314 = _40313 ^ _6134;
  wire _40315 = _924 ^ _39910;
  wire _40316 = _15114 ^ _6780;
  wire _40317 = _40315 ^ _40316;
  wire _40318 = _40314 ^ _40317;
  wire _40319 = _1745 ^ _932;
  wire _40320 = _40319 ^ _13577;
  wire _40321 = _78 ^ _12467;
  wire _40322 = _4057 ^ _941;
  wire _40323 = _40321 ^ _40322;
  wire _40324 = _40320 ^ _40323;
  wire _40325 = _40318 ^ _40324;
  wire _40326 = _1761 ^ _17113;
  wire _40327 = _19549 ^ _6811;
  wire _40328 = uncoded_block[221] ^ uncoded_block[228];
  wire _40329 = _40328 ^ _1774;
  wire _40330 = _40327 ^ _40329;
  wire _40331 = _40326 ^ _40330;
  wire _40332 = uncoded_block[239] ^ uncoded_block[246];
  wire _40333 = _970 ^ _40332;
  wire _40334 = _11948 ^ _40333;
  wire _40335 = _20021 ^ _9761;
  wire _40336 = _40335 ^ _26892;
  wire _40337 = _40334 ^ _40336;
  wire _40338 = _40331 ^ _40337;
  wire _40339 = _40325 ^ _40338;
  wire _40340 = _40311 ^ _40339;
  wire _40341 = uncoded_block[263] ^ uncoded_block[267];
  wire _40342 = _40341 ^ _4811;
  wire _40343 = _9222 ^ _12506;
  wire _40344 = _40342 ^ _40343;
  wire _40345 = _4106 ^ _26011;
  wire _40346 = _40344 ^ _40345;
  wire _40347 = _4820 ^ _8636;
  wire _40348 = _40347 ^ _28068;
  wire _40349 = _5530 ^ _4123;
  wire _40350 = _1007 ^ _40349;
  wire _40351 = _40348 ^ _40350;
  wire _40352 = _40346 ^ _40351;
  wire _40353 = _1014 ^ _9235;
  wire _40354 = _9240 ^ _10323;
  wire _40355 = _40353 ^ _40354;
  wire _40356 = _4841 ^ _159;
  wire _40357 = _1023 ^ _36782;
  wire _40358 = _40356 ^ _40357;
  wire _40359 = _40355 ^ _40358;
  wire _40360 = uncoded_block[363] ^ uncoded_block[367];
  wire _40361 = _3365 ^ _40360;
  wire _40362 = _3363 ^ _40361;
  wire _40363 = _1036 ^ _6233;
  wire _40364 = _22415 ^ _40363;
  wire _40365 = _40362 ^ _40364;
  wire _40366 = _40359 ^ _40365;
  wire _40367 = _40352 ^ _40366;
  wire _40368 = _17661 ^ _2613;
  wire _40369 = _36788 ^ _40368;
  wire _40370 = _2615 ^ _19604;
  wire _40371 = _31870 ^ _181;
  wire _40372 = _40370 ^ _40371;
  wire _40373 = _40369 ^ _40372;
  wire _40374 = uncoded_block[410] ^ uncoded_block[415];
  wire _40375 = _24703 ^ _40374;
  wire _40376 = _40375 ^ _9268;
  wire _40377 = uncoded_block[429] ^ uncoded_block[435];
  wire _40378 = _40377 ^ _16187;
  wire _40379 = _6252 ^ _40378;
  wire _40380 = _40376 ^ _40379;
  wire _40381 = _40373 ^ _40380;
  wire _40382 = _5584 ^ _27354;
  wire _40383 = _17183 ^ _40382;
  wire _40384 = _4186 ^ _16692;
  wire _40385 = _12567 ^ _40384;
  wire _40386 = _40383 ^ _40385;
  wire _40387 = _21526 ^ _21528;
  wire _40388 = _12577 ^ _21987;
  wire _40389 = _40387 ^ _40388;
  wire _40390 = _5604 ^ _2668;
  wire _40391 = _40390 ^ _4206;
  wire _40392 = _40389 ^ _40391;
  wire _40393 = _40386 ^ _40392;
  wire _40394 = _40381 ^ _40393;
  wire _40395 = _40367 ^ _40394;
  wire _40396 = _40340 ^ _40395;
  wire _40397 = _23370 ^ _4918;
  wire _40398 = _1108 ^ _4922;
  wire _40399 = _40397 ^ _40398;
  wire _40400 = uncoded_block[534] ^ uncoded_block[540];
  wire _40401 = _9309 ^ _40400;
  wire _40402 = _40401 ^ _13691;
  wire _40403 = _40399 ^ _40402;
  wire _40404 = _3465 ^ _6309;
  wire _40405 = _31046 ^ _40404;
  wire _40406 = _21561 ^ _15748;
  wire _40407 = _40405 ^ _40406;
  wire _40408 = _40403 ^ _40407;
  wire _40409 = _18222 ^ _3480;
  wire _40410 = _25190 ^ _40409;
  wire _40411 = _12066 ^ _2707;
  wire _40412 = _11535 ^ _6325;
  wire _40413 = _40411 ^ _40412;
  wire _40414 = _40410 ^ _40413;
  wire _40415 = _22024 ^ _29318;
  wire _40416 = _12070 ^ _40415;
  wire _40417 = _8161 ^ _290;
  wire _40418 = uncoded_block[636] ^ uncoded_block[645];
  wire _40419 = _40418 ^ _10425;
  wire _40420 = _40417 ^ _40419;
  wire _40421 = _40416 ^ _40420;
  wire _40422 = _40414 ^ _40421;
  wire _40423 = _40408 ^ _40422;
  wire _40424 = _14234 ^ _302;
  wire _40425 = _40424 ^ _32757;
  wire _40426 = _4262 ^ _309;
  wire _40427 = uncoded_block[671] ^ uncoded_block[674];
  wire _40428 = _40427 ^ _12634;
  wire _40429 = _40426 ^ _40428;
  wire _40430 = _40425 ^ _40429;
  wire _40431 = _2751 ^ _13735;
  wire _40432 = _18248 ^ _40431;
  wire _40433 = _6990 ^ _10445;
  wire _40434 = uncoded_block[708] ^ uncoded_block[713];
  wire _40435 = _14255 ^ _40434;
  wire _40436 = _40433 ^ _40435;
  wire _40437 = _40432 ^ _40436;
  wire _40438 = _40430 ^ _40437;
  wire _40439 = _4999 ^ _17762;
  wire _40440 = _341 ^ _344;
  wire _40441 = _40439 ^ _40440;
  wire _40442 = _20153 ^ _352;
  wire _40443 = _29338 ^ _40442;
  wire _40444 = _40441 ^ _40443;
  wire _40445 = _5702 ^ _36873;
  wire _40446 = _5016 ^ _4298;
  wire _40447 = _40445 ^ _40446;
  wire _40448 = _31101 ^ _18744;
  wire _40449 = _40447 ^ _40448;
  wire _40450 = _40444 ^ _40449;
  wire _40451 = _40438 ^ _40450;
  wire _40452 = _40423 ^ _40451;
  wire _40453 = _11019 ^ _35257;
  wire _40454 = _13219 ^ _31106;
  wire _40455 = _40453 ^ _40454;
  wire _40456 = _1224 ^ _3574;
  wire _40457 = _14282 ^ _4316;
  wire _40458 = _40456 ^ _40457;
  wire _40459 = _40455 ^ _40458;
  wire _40460 = _34062 ^ _392;
  wire _40461 = _5729 ^ _29788;
  wire _40462 = _40460 ^ _40461;
  wire _40463 = _3587 ^ _7039;
  wire _40464 = _2033 ^ _16801;
  wire _40465 = _40463 ^ _40464;
  wire _40466 = _40462 ^ _40465;
  wire _40467 = _40459 ^ _40466;
  wire _40468 = _9938 ^ _2036;
  wire _40469 = _7047 ^ _4340;
  wire _40470 = _40468 ^ _40469;
  wire _40471 = _6406 ^ _2046;
  wire _40472 = _14300 ^ _6410;
  wire _40473 = _40471 ^ _40472;
  wire _40474 = _40470 ^ _40473;
  wire _40475 = _27452 ^ _35281;
  wire _40476 = _40475 ^ _12699;
  wire _40477 = _28212 ^ _13803;
  wire _40478 = _40476 ^ _40477;
  wire _40479 = _40474 ^ _40478;
  wire _40480 = _40467 ^ _40479;
  wire _40481 = _19251 ^ _435;
  wire _40482 = _12712 ^ _3631;
  wire _40483 = _40481 ^ _40482;
  wire _40484 = uncoded_block[921] ^ uncoded_block[924];
  wire _40485 = _40484 ^ _4370;
  wire _40486 = _40485 ^ _14837;
  wire _40487 = _40483 ^ _40486;
  wire _40488 = _1299 ^ _1302;
  wire _40489 = _460 ^ _2089;
  wire _40490 = _40488 ^ _40489;
  wire _40491 = _463 ^ _24388;
  wire _40492 = _11648 ^ _471;
  wire _40493 = _40491 ^ _40492;
  wire _40494 = _40490 ^ _40493;
  wire _40495 = _40487 ^ _40494;
  wire _40496 = _7093 ^ _1317;
  wire _40497 = uncoded_block[995] ^ uncoded_block[998];
  wire _40498 = _23939 ^ _40497;
  wire _40499 = _40496 ^ _40498;
  wire _40500 = _7691 ^ _2112;
  wire _40501 = _11661 ^ _4410;
  wire _40502 = _40500 ^ _40501;
  wire _40503 = _40499 ^ _40502;
  wire _40504 = _2117 ^ _9996;
  wire _40505 = _40504 ^ _32435;
  wire _40506 = _5138 ^ _12756;
  wire _40507 = _40506 ^ _503;
  wire _40508 = _40505 ^ _40507;
  wire _40509 = _40503 ^ _40508;
  wire _40510 = _40495 ^ _40509;
  wire _40511 = _40480 ^ _40510;
  wire _40512 = _40452 ^ _40511;
  wire _40513 = _40396 ^ _40512;
  wire _40514 = _24408 ^ _40124;
  wire _40515 = _40514 ^ _6480;
  wire _40516 = _12764 ^ _35719;
  wire _40517 = _15395 ^ _1366;
  wire _40518 = _40516 ^ _40517;
  wire _40519 = _40515 ^ _40518;
  wire _40520 = _12219 ^ _17363;
  wire _40521 = _18817 ^ _40520;
  wire _40522 = _19306 ^ _537;
  wire _40523 = _3704 ^ _545;
  wire _40524 = _40522 ^ _40523;
  wire _40525 = _40521 ^ _40524;
  wire _40526 = _40519 ^ _40525;
  wire _40527 = _30322 ^ _9488;
  wire _40528 = uncoded_block[1124] ^ uncoded_block[1126];
  wire _40529 = _40528 ^ _2945;
  wire _40530 = _25328 ^ _40529;
  wire _40531 = _40527 ^ _40530;
  wire _40532 = _14887 ^ _10593;
  wire _40533 = _16380 ^ _7141;
  wire _40534 = _40532 ^ _40533;
  wire _40535 = _24900 ^ _10044;
  wire _40536 = _40534 ^ _40535;
  wire _40537 = _40531 ^ _40536;
  wire _40538 = _40526 ^ _40537;
  wire _40539 = uncoded_block[1166] ^ uncoded_block[1169];
  wire _40540 = _40539 ^ _7154;
  wire _40541 = _14901 ^ _592;
  wire _40542 = _40540 ^ _40541;
  wire _40543 = _10053 ^ _4488;
  wire _40544 = _40543 ^ _14909;
  wire _40545 = _40542 ^ _40544;
  wire _40546 = _2974 ^ _24001;
  wire _40547 = _14914 ^ _4502;
  wire _40548 = _40546 ^ _40547;
  wire _40549 = _2226 ^ _19827;
  wire _40550 = _9523 ^ _40549;
  wire _40551 = _40548 ^ _40550;
  wire _40552 = _40545 ^ _40551;
  wire _40553 = _27129 ^ _33758;
  wire _40554 = _22651 ^ _624;
  wire _40555 = _40553 ^ _40554;
  wire _40556 = _3003 ^ _3786;
  wire _40557 = _40556 ^ _2246;
  wire _40558 = _40555 ^ _40557;
  wire _40559 = _2247 ^ _3011;
  wire _40560 = _6560 ^ _13380;
  wire _40561 = _40559 ^ _40560;
  wire _40562 = _18419 ^ _22662;
  wire _40563 = _40562 ^ _12284;
  wire _40564 = _40561 ^ _40563;
  wire _40565 = _40558 ^ _40564;
  wire _40566 = _40552 ^ _40565;
  wire _40567 = _40538 ^ _40566;
  wire _40568 = _14430 ^ _2262;
  wire _40569 = _34177 ^ _40568;
  wire _40570 = _3029 ^ _3032;
  wire _40571 = _657 ^ _5931;
  wire _40572 = _40570 ^ _40571;
  wire _40573 = _40569 ^ _40572;
  wire _40574 = _5262 ^ _3039;
  wire _40575 = _35781 ^ _40574;
  wire _40576 = _669 ^ _15473;
  wire _40577 = _15477 ^ _27157;
  wire _40578 = _40576 ^ _40577;
  wire _40579 = _40575 ^ _40578;
  wire _40580 = _40573 ^ _40579;
  wire _40581 = uncoded_block[1364] ^ uncoded_block[1367];
  wire _40582 = _40581 ^ _22224;
  wire _40583 = _40582 ^ _24506;
  wire _40584 = _3061 ^ _21771;
  wire _40585 = _7827 ^ _40584;
  wire _40586 = _40583 ^ _40585;
  wire _40587 = _5952 ^ _20835;
  wire _40588 = uncoded_block[1401] ^ uncoded_block[1407];
  wire _40589 = _40588 ^ _5957;
  wire _40590 = _40587 ^ _40589;
  wire _40591 = _4580 ^ _705;
  wire _40592 = _7842 ^ _32948;
  wire _40593 = _40591 ^ _40592;
  wire _40594 = _40590 ^ _40593;
  wire _40595 = _40586 ^ _40594;
  wire _40596 = _40580 ^ _40595;
  wire _40597 = _14467 ^ _3861;
  wire _40598 = _40597 ^ _35025;
  wire _40599 = _14983 ^ _3088;
  wire _40600 = _7241 ^ _9602;
  wire _40601 = _40599 ^ _40600;
  wire _40602 = _40598 ^ _40601;
  wire _40603 = uncoded_block[1468] ^ uncoded_block[1474];
  wire _40604 = _40603 ^ _3881;
  wire _40605 = _3100 ^ _5320;
  wire _40606 = _40604 ^ _40605;
  wire _40607 = uncoded_block[1491] ^ uncoded_block[1496];
  wire _40608 = _40607 ^ _3891;
  wire _40609 = _31716 ^ _40608;
  wire _40610 = _40606 ^ _40609;
  wire _40611 = _40602 ^ _40610;
  wire _40612 = uncoded_block[1504] ^ uncoded_block[1510];
  wire _40613 = _40612 ^ _7875;
  wire _40614 = _40613 ^ _7877;
  wire _40615 = _5341 ^ _8473;
  wire _40616 = _40615 ^ _39437;
  wire _40617 = _40614 ^ _40616;
  wire _40618 = _36235 ^ _19904;
  wire _40619 = _14496 ^ _6657;
  wire _40620 = _15527 ^ _40619;
  wire _40621 = _40618 ^ _40620;
  wire _40622 = _40617 ^ _40621;
  wire _40623 = _40611 ^ _40622;
  wire _40624 = _40596 ^ _40623;
  wire _40625 = _40567 ^ _40624;
  wire _40626 = _32985 ^ _2376;
  wire _40627 = _777 ^ _15026;
  wire _40628 = _40626 ^ _40627;
  wire _40629 = _17510 ^ _25009;
  wire _40630 = _40628 ^ _40629;
  wire _40631 = _29550 ^ _11847;
  wire _40632 = _34245 ^ _40631;
  wire _40633 = uncoded_block[1602] ^ uncoded_block[1607];
  wire _40634 = _40633 ^ _6040;
  wire _40635 = _801 ^ _10181;
  wire _40636 = _40634 ^ _40635;
  wire _40637 = _40632 ^ _40636;
  wire _40638 = _40630 ^ _40637;
  wire _40639 = _3160 ^ _5386;
  wire _40640 = _1636 ^ _6048;
  wire _40641 = _40639 ^ _40640;
  wire _40642 = _1641 ^ _12949;
  wire _40643 = _7309 ^ _12387;
  wire _40644 = _40642 ^ _40643;
  wire _40645 = _40641 ^ _40644;
  wire _40646 = _4680 ^ _2419;
  wire _40647 = _40260 ^ _40646;
  wire _40648 = _3182 ^ _36269;
  wire _40649 = _24585 ^ _40648;
  wire _40650 = _40647 ^ _40649;
  wire _40651 = _40645 ^ _40650;
  wire _40652 = _40638 ^ _40651;
  wire _40653 = _3186 ^ _4691;
  wire _40654 = _40653 ^ _19476;
  wire _40655 = _2435 ^ _3980;
  wire _40656 = _26833 ^ _40655;
  wire _40657 = _40654 ^ _40656;
  wire _40658 = _40657 ^ _23240;
  wire _40659 = _40652 ^ _40658;
  wire _40660 = _40625 ^ _40659;
  wire _40661 = _40513 ^ _40660;
  wire _40662 = _15582 ^ _18057;
  wire _40663 = _40662 ^ _18059;
  wire _40664 = _7351 ^ _10791;
  wire _40665 = _5427 ^ _11890;
  wire _40666 = _40664 ^ _40665;
  wire _40667 = _40663 ^ _40666;
  wire _40668 = _18548 ^ _8549;
  wire _40669 = _21416 ^ _5435;
  wire _40670 = _40668 ^ _40669;
  wire _40671 = _10238 ^ _31;
  wire _40672 = _10806 ^ _4728;
  wire _40673 = _40671 ^ _40672;
  wire _40674 = _40670 ^ _40673;
  wire _40675 = _40667 ^ _40674;
  wire _40676 = _26393 ^ _5443;
  wire _40677 = _40676 ^ _21885;
  wire _40678 = _14586 ^ _15603;
  wire _40679 = _1718 ^ _12443;
  wire _40680 = _40678 ^ _40679;
  wire _40681 = _40677 ^ _40680;
  wire _40682 = _49 ^ _2490;
  wire _40683 = _2491 ^ _7990;
  wire _40684 = _40682 ^ _40683;
  wire _40685 = uncoded_block[121] ^ uncoded_block[126];
  wire _40686 = _40685 ^ _8579;
  wire _40687 = _3263 ^ _9730;
  wire _40688 = _40686 ^ _40687;
  wire _40689 = _40684 ^ _40688;
  wire _40690 = _40681 ^ _40689;
  wire _40691 = _40675 ^ _40690;
  wire _40692 = _30945 ^ _6780;
  wire _40693 = _7397 ^ _4049;
  wire _40694 = _40692 ^ _40693;
  wire _40695 = _29208 ^ _15123;
  wire _40696 = _82 ^ _3281;
  wire _40697 = _40695 ^ _40696;
  wire _40698 = _40694 ^ _40697;
  wire _40699 = _20004 ^ _13588;
  wire _40700 = _40699 ^ _30079;
  wire _40701 = _28043 ^ _7415;
  wire _40702 = _14100 ^ _40701;
  wire _40703 = _40700 ^ _40702;
  wire _40704 = _40698 ^ _40703;
  wire _40705 = _6161 ^ _8606;
  wire _40706 = uncoded_block[225] ^ uncoded_block[233];
  wire _40707 = _40706 ^ _10289;
  wire _40708 = _40705 ^ _40707;
  wire _40709 = _4085 ^ _8617;
  wire _40710 = _10293 ^ _40709;
  wire _40711 = _40708 ^ _40710;
  wire _40712 = uncoded_block[252] ^ uncoded_block[256];
  wire _40713 = _40712 ^ _4095;
  wire _40714 = _15154 ^ _6192;
  wire _40715 = _40713 ^ _40714;
  wire _40716 = uncoded_block[282] ^ uncoded_block[286];
  wire _40717 = _10303 ^ _40716;
  wire _40718 = _38762 ^ _13615;
  wire _40719 = _40717 ^ _40718;
  wire _40720 = _40715 ^ _40719;
  wire _40721 = _40711 ^ _40720;
  wire _40722 = _40704 ^ _40721;
  wire _40723 = _40691 ^ _40722;
  wire _40724 = uncoded_block[306] ^ uncoded_block[313];
  wire _40725 = _142 ^ _40724;
  wire _40726 = uncoded_block[315] ^ uncoded_block[320];
  wire _40727 = _40726 ^ _8642;
  wire _40728 = _40725 ^ _40727;
  wire _40729 = _30117 ^ _4125;
  wire _40730 = _13629 ^ _6217;
  wire _40731 = _40729 ^ _40730;
  wire _40732 = _40728 ^ _40731;
  wire _40733 = uncoded_block[344] ^ uncoded_block[350];
  wire _40734 = _40733 ^ _15179;
  wire _40735 = uncoded_block[356] ^ uncoded_block[366];
  wire _40736 = _40735 ^ _1835;
  wire _40737 = _40734 ^ _40736;
  wire _40738 = uncoded_block[375] ^ uncoded_block[379];
  wire _40739 = _169 ^ _40738;
  wire _40740 = _40739 ^ _10337;
  wire _40741 = _40737 ^ _40740;
  wire _40742 = _40732 ^ _40741;
  wire _40743 = _2613 ^ _6239;
  wire _40744 = _40743 ^ _23782;
  wire _40745 = _24243 ^ _21508;
  wire _40746 = _24704 ^ _40745;
  wire _40747 = _40744 ^ _40746;
  wire _40748 = uncoded_block[417] ^ uncoded_block[422];
  wire _40749 = _40748 ^ _16184;
  wire _40750 = _9820 ^ _21049;
  wire _40751 = _40749 ^ _40750;
  wire _40752 = _9275 ^ _1075;
  wire _40753 = _3415 ^ _4890;
  wire _40754 = _40752 ^ _40753;
  wire _40755 = _40751 ^ _40754;
  wire _40756 = _40747 ^ _40755;
  wire _40757 = _40742 ^ _40756;
  wire _40758 = _1079 ^ _26944;
  wire _40759 = _3421 ^ _16693;
  wire _40760 = _40758 ^ _40759;
  wire _40761 = uncoded_block[488] ^ uncoded_block[494];
  wire _40762 = _8694 ^ _40761;
  wire _40763 = _5603 ^ _2667;
  wire _40764 = _40762 ^ _40763;
  wire _40765 = _40760 ^ _40764;
  wire _40766 = _3437 ^ _3439;
  wire _40767 = _8121 ^ _40766;
  wire _40768 = uncoded_block[515] ^ uncoded_block[528];
  wire _40769 = _40768 ^ _20603;
  wire _40770 = _4215 ^ _4217;
  wire _40771 = _40769 ^ _40770;
  wire _40772 = _40767 ^ _40771;
  wire _40773 = _40765 ^ _40772;
  wire _40774 = _7541 ^ _6300;
  wire _40775 = _40774 ^ _29301;
  wire _40776 = _1916 ^ _258;
  wire _40777 = _1126 ^ _39617;
  wire _40778 = _40776 ^ _40777;
  wire _40779 = _40775 ^ _40778;
  wire _40780 = _26528 ^ _4234;
  wire _40781 = _16723 ^ _40780;
  wire _40782 = _1142 ^ _278;
  wire _40783 = _12062 ^ _40782;
  wire _40784 = _40781 ^ _40783;
  wire _40785 = _40779 ^ _40784;
  wire _40786 = _40773 ^ _40785;
  wire _40787 = _40757 ^ _40786;
  wire _40788 = _40723 ^ _40787;
  wire _40789 = _7563 ^ _4243;
  wire _40790 = _40789 ^ _30196;
  wire _40791 = _1154 ^ _1156;
  wire _40792 = _30199 ^ _293;
  wire _40793 = _40791 ^ _40792;
  wire _40794 = _40790 ^ _40793;
  wire _40795 = _28528 ^ _12626;
  wire _40796 = _302 ^ _304;
  wire _40797 = _16747 ^ _14238;
  wire _40798 = _40796 ^ _40797;
  wire _40799 = _40795 ^ _40798;
  wire _40800 = _40794 ^ _40799;
  wire _40801 = _9355 ^ _311;
  wire _40802 = _1178 ^ _1180;
  wire _40803 = _40801 ^ _40802;
  wire _40804 = _3526 ^ _18249;
  wire _40805 = _12641 ^ _4995;
  wire _40806 = _40804 ^ _40805;
  wire _40807 = _40803 ^ _40806;
  wire _40808 = _3535 ^ _17266;
  wire _40809 = _9902 ^ _5693;
  wire _40810 = _40808 ^ _40809;
  wire _40811 = _11573 ^ _23425;
  wire _40812 = _20156 ^ _5013;
  wire _40813 = _40811 ^ _40812;
  wire _40814 = _40810 ^ _40813;
  wire _40815 = _40807 ^ _40814;
  wire _40816 = _40800 ^ _40815;
  wire _40817 = uncoded_block[750] ^ uncoded_block[753];
  wire _40818 = uncoded_block[755] ^ uncoded_block[761];
  wire _40819 = _40817 ^ _40818;
  wire _40820 = uncoded_block[766] ^ uncoded_block[771];
  wire _40821 = _364 ^ _40820;
  wire _40822 = _40819 ^ _40821;
  wire _40823 = _13219 ^ _1224;
  wire _40824 = _40823 ^ _22519;
  wire _40825 = _40822 ^ _40824;
  wire _40826 = _383 ^ _385;
  wire _40827 = _22071 ^ _392;
  wire _40828 = _40826 ^ _40827;
  wire _40829 = _2809 ^ _2812;
  wire _40830 = _28949 ^ _40829;
  wire _40831 = _40828 ^ _40830;
  wire _40832 = _40825 ^ _40831;
  wire _40833 = _4336 ^ _4339;
  wire _40834 = _1257 ^ _12141;
  wire _40835 = _40833 ^ _40834;
  wire _40836 = _2821 ^ _5066;
  wire _40837 = _7054 ^ _35281;
  wire _40838 = _40836 ^ _40837;
  wire _40839 = _40835 ^ _40838;
  wire _40840 = _33671 ^ _20696;
  wire _40841 = uncoded_block[888] ^ uncoded_block[892];
  wire _40842 = _8820 ^ _40841;
  wire _40843 = _40840 ^ _40842;
  wire _40844 = _14829 ^ _14316;
  wire _40845 = _6428 ^ _5762;
  wire _40846 = _40844 ^ _40845;
  wire _40847 = _40843 ^ _40846;
  wire _40848 = _40839 ^ _40847;
  wire _40849 = _40832 ^ _40848;
  wire _40850 = _40816 ^ _40849;
  wire _40851 = _8835 ^ _8262;
  wire _40852 = _38904 ^ _40851;
  wire _40853 = _24383 ^ _460;
  wire _40854 = _5779 ^ _10525;
  wire _40855 = _40853 ^ _40854;
  wire _40856 = _40852 ^ _40855;
  wire _40857 = _9981 ^ _28233;
  wire _40858 = uncoded_block[992] ^ uncoded_block[996];
  wire _40859 = _18329 ^ _40858;
  wire _40860 = _40857 ^ _40859;
  wire _40861 = _11101 ^ _2111;
  wire _40862 = _40861 ^ _18343;
  wire _40863 = _40860 ^ _40862;
  wire _40864 = _40856 ^ _40863;
  wire _40865 = _8871 ^ _27494;
  wire _40866 = _35706 ^ _40865;
  wire _40867 = _498 ^ _11668;
  wire _40868 = _1342 ^ _8306;
  wire _40869 = _40867 ^ _40868;
  wire _40870 = _40866 ^ _40869;
  wire _40871 = uncoded_block[1046] ^ uncoded_block[1051];
  wire _40872 = _40871 ^ _12762;
  wire _40873 = _4430 ^ _10566;
  wire _40874 = _40872 ^ _40873;
  wire _40875 = _2917 ^ _6485;
  wire _40876 = uncoded_block[1071] ^ uncoded_block[1078];
  wire _40877 = uncoded_block[1079] ^ uncoded_block[1083];
  wire _40878 = _40876 ^ _40877;
  wire _40879 = _40875 ^ _40878;
  wire _40880 = _40874 ^ _40879;
  wire _40881 = _40870 ^ _40880;
  wire _40882 = _40864 ^ _40881;
  wire _40883 = _4438 ^ _23508;
  wire _40884 = uncoded_block[1096] ^ uncoded_block[1104];
  wire _40885 = _40884 ^ _3708;
  wire _40886 = _40883 ^ _40885;
  wire _40887 = _1385 ^ _8917;
  wire _40888 = _3713 ^ _7736;
  wire _40889 = _40887 ^ _40888;
  wire _40890 = _40886 ^ _40889;
  wire _40891 = _8342 ^ _23981;
  wire _40892 = _40891 ^ _38961;
  wire _40893 = _2953 ^ _10597;
  wire _40894 = uncoded_block[1148] ^ uncoded_block[1157];
  wire _40895 = _40894 ^ _22627;
  wire _40896 = _40893 ^ _40895;
  wire _40897 = _40892 ^ _40896;
  wire _40898 = _40890 ^ _40897;
  wire _40899 = uncoded_block[1174] ^ uncoded_block[1179];
  wire _40900 = _40899 ^ _4482;
  wire _40901 = _18844 ^ _40900;
  wire _40902 = _5200 ^ _4488;
  wire _40903 = uncoded_block[1195] ^ uncoded_block[1202];
  wire _40904 = uncoded_block[1203] ^ uncoded_block[1208];
  wire _40905 = _40903 ^ _40904;
  wire _40906 = _40902 ^ _40905;
  wire _40907 = _40901 ^ _40906;
  wire _40908 = uncoded_block[1210] ^ uncoded_block[1217];
  wire _40909 = _40908 ^ _10059;
  wire _40910 = _7168 ^ _4504;
  wire _40911 = _40909 ^ _40910;
  wire _40912 = _22188 ^ _3772;
  wire _40913 = uncoded_block[1240] ^ uncoded_block[1247];
  wire _40914 = uncoded_block[1248] ^ uncoded_block[1254];
  wire _40915 = _40913 ^ _40914;
  wire _40916 = _40912 ^ _40915;
  wire _40917 = _40911 ^ _40916;
  wire _40918 = _40907 ^ _40917;
  wire _40919 = _40898 ^ _40918;
  wire _40920 = _40882 ^ _40919;
  wire _40921 = _40850 ^ _40920;
  wire _40922 = _40788 ^ _40921;
  wire _40923 = _35373 ^ _38581;
  wire _40924 = _22197 ^ _5907;
  wire _40925 = uncoded_block[1287] ^ uncoded_block[1292];
  wire _40926 = _6556 ^ _40925;
  wire _40927 = _40924 ^ _40926;
  wire _40928 = _40923 ^ _40927;
  wire _40929 = _13388 ^ _6571;
  wire _40930 = _40929 ^ _24938;
  wire _40931 = _21748 ^ _3028;
  wire _40932 = uncoded_block[1322] ^ uncoded_block[1326];
  wire _40933 = uncoded_block[1327] ^ uncoded_block[1332];
  wire _40934 = _40932 ^ _40933;
  wire _40935 = _40931 ^ _40934;
  wire _40936 = _40930 ^ _40935;
  wire _40937 = _40928 ^ _40936;
  wire _40938 = _21298 ^ _1501;
  wire _40939 = _26731 ^ _40938;
  wire _40940 = _14442 ^ _33363;
  wire _40941 = uncoded_block[1355] ^ uncoded_block[1359];
  wire _40942 = _40941 ^ _10665;
  wire _40943 = _40940 ^ _40942;
  wire _40944 = _40939 ^ _40943;
  wire _40945 = uncoded_block[1370] ^ uncoded_block[1374];
  wire _40946 = _10668 ^ _40945;
  wire _40947 = _9573 ^ _4564;
  wire _40948 = _40946 ^ _40947;
  wire _40949 = uncoded_block[1386] ^ uncoded_block[1397];
  wire _40950 = _10108 ^ _40949;
  wire _40951 = _40950 ^ _23159;
  wire _40952 = _40948 ^ _40951;
  wire _40953 = _40944 ^ _40952;
  wire _40954 = _40937 ^ _40953;
  wire _40955 = _11236 ^ _4580;
  wire _40956 = uncoded_block[1415] ^ uncoded_block[1421];
  wire _40957 = _40956 ^ _2308;
  wire _40958 = _40955 ^ _40957;
  wire _40959 = _22242 ^ _23169;
  wire _40960 = _27172 ^ _40959;
  wire _40961 = _40958 ^ _40960;
  wire _40962 = _3084 ^ _717;
  wire _40963 = _2326 ^ _13440;
  wire _40964 = _40962 ^ _40963;
  wire _40965 = _7247 ^ _14989;
  wire _40966 = _4604 ^ _2344;
  wire _40967 = _40965 ^ _40966;
  wire _40968 = _40964 ^ _40967;
  wire _40969 = _40961 ^ _40968;
  wire _40970 = _5988 ^ _5329;
  wire _40971 = uncoded_block[1498] ^ uncoded_block[1505];
  wire _40972 = _6631 ^ _40971;
  wire _40973 = _40970 ^ _40972;
  wire _40974 = uncoded_block[1506] ^ uncoded_block[1512];
  wire _40975 = _40974 ^ _18480;
  wire _40976 = _40975 ^ _10150;
  wire _40977 = _40973 ^ _40976;
  wire _40978 = _13978 ^ _31309;
  wire _40979 = uncoded_block[1546] ^ uncoded_block[1556];
  wire _40980 = _6651 ^ _40979;
  wire _40981 = _40978 ^ _40980;
  wire _40982 = _1597 ^ _2376;
  wire _40983 = _4644 ^ _16020;
  wire _40984 = _40982 ^ _40983;
  wire _40985 = _40981 ^ _40984;
  wire _40986 = _40977 ^ _40985;
  wire _40987 = _40969 ^ _40986;
  wire _40988 = _40954 ^ _40987;
  wire _40989 = uncoded_block[1574] ^ uncoded_block[1581];
  wire _40990 = _40989 ^ _15537;
  wire _40991 = _4653 ^ _791;
  wire _40992 = _40990 ^ _40991;
  wire _40993 = _39062 ^ _1621;
  wire _40994 = _3153 ^ _6677;
  wire _40995 = _40993 ^ _40994;
  wire _40996 = _40992 ^ _40995;
  wire _40997 = _7906 ^ _17020;
  wire _40998 = uncoded_block[1621] ^ uncoded_block[1627];
  wire _40999 = _12376 ^ _40998;
  wire _41000 = _40997 ^ _40999;
  wire _41001 = uncoded_block[1646] ^ uncoded_block[1652];
  wire _41002 = _24576 ^ _41001;
  wire _41003 = _39462 ^ _41002;
  wire _41004 = _41000 ^ _41003;
  wire _41005 = _40996 ^ _41004;
  wire _41006 = _4678 ^ _29569;
  wire _41007 = _16537 ^ _4687;
  wire _41008 = _41006 ^ _41007;
  wire _41009 = uncoded_block[1671] ^ uncoded_block[1675];
  wire _41010 = uncoded_block[1677] ^ uncoded_block[1682];
  wire _41011 = _41009 ^ _41010;
  wire _41012 = _14543 ^ _10768;
  wire _41013 = _41011 ^ _41012;
  wire _41014 = _41008 ^ _41013;
  wire _41015 = _8533 ^ _20920;
  wire _41016 = _29576 ^ _41015;
  wire _41017 = _15063 ^ _19953;
  wire _41018 = _854 ^ _3988;
  wire _41019 = _41017 ^ _41018;
  wire _41020 = _41016 ^ _41019;
  wire _41021 = _41014 ^ _41020;
  wire _41022 = _41005 ^ _41021;
  wire _41023 = _41022 ^ uncoded_block[1722];
  wire _41024 = _40988 ^ _41023;
  wire _41025 = _40922 ^ _41024;
  wire _41026 = uncoded_block[1] ^ uncoded_block[7];
  wire _41027 = _41026 ^ _18057;
  wire _41028 = _41027 ^ _36289;
  wire _41029 = _10226 ^ _7353;
  wire _41030 = _9694 ^ _1693;
  wire _41031 = _41029 ^ _41030;
  wire _41032 = _41028 ^ _41031;
  wire _41033 = _15080 ^ _879;
  wire _41034 = _41033 ^ _20;
  wire _41035 = _7968 ^ _16572;
  wire _41036 = _12426 ^ _41035;
  wire _41037 = _41034 ^ _41036;
  wire _41038 = _41032 ^ _41037;
  wire _41039 = _13553 ^ _34688;
  wire _41040 = _41039 ^ _29190;
  wire _41041 = _2481 ^ _4735;
  wire _41042 = _41041 ^ _12441;
  wire _41043 = _41040 ^ _41042;
  wire _41044 = uncoded_block[89] ^ uncoded_block[94];
  wire _41045 = _41044 ^ _6758;
  wire _41046 = _41045 ^ _40303;
  wire _41047 = _1721 ^ _4034;
  wire _41048 = _41047 ^ _21435;
  wire _41049 = _41046 ^ _41048;
  wire _41050 = _41043 ^ _41049;
  wire _41051 = _41038 ^ _41050;
  wire _41052 = _20963 ^ _25075;
  wire _41053 = _15618 ^ _41052;
  wire _41054 = _3265 ^ _11924;
  wire _41055 = _14082 ^ _31393;
  wire _41056 = _41054 ^ _41055;
  wire _41057 = _41053 ^ _41056;
  wire _41058 = _4048 ^ _20975;
  wire _41059 = _4054 ^ _1751;
  wire _41060 = _41058 ^ _41059;
  wire _41061 = uncoded_block[173] ^ uncoded_block[176];
  wire _41062 = _6788 ^ _41061;
  wire _41063 = _41062 ^ _39135;
  wire _41064 = _41060 ^ _41063;
  wire _41065 = _41057 ^ _41064;
  wire _41066 = _86 ^ _4062;
  wire _41067 = _41066 ^ _13589;
  wire _41068 = uncoded_block[195] ^ uncoded_block[198];
  wire _41069 = _4776 ^ _41068;
  wire _41070 = _41069 ^ _22839;
  wire _41071 = _41067 ^ _41070;
  wire _41072 = _8600 ^ _19549;
  wire _41073 = _8606 ^ _7419;
  wire _41074 = _41072 ^ _41073;
  wire _41075 = _17118 ^ _6821;
  wire _41076 = _33088 ^ _7425;
  wire _41077 = _41075 ^ _41076;
  wire _41078 = _41074 ^ _41077;
  wire _41079 = _41071 ^ _41078;
  wire _41080 = _41065 ^ _41079;
  wire _41081 = _41051 ^ _41080;
  wire _41082 = _10860 ^ _1781;
  wire _41083 = _11954 ^ _20520;
  wire _41084 = _41082 ^ _41083;
  wire _41085 = _7441 ^ _19570;
  wire _41086 = _26443 ^ _41085;
  wire _41087 = _41084 ^ _41086;
  wire _41088 = _7446 ^ _8632;
  wire _41089 = _15159 ^ _995;
  wire _41090 = _41088 ^ _41089;
  wire _41091 = uncoded_block[303] ^ uncoded_block[307];
  wire _41092 = _21483 ^ _41091;
  wire _41093 = _21017 ^ _3338;
  wire _41094 = _41092 ^ _41093;
  wire _41095 = _41090 ^ _41094;
  wire _41096 = _41087 ^ _41095;
  wire _41097 = _1008 ^ _3346;
  wire _41098 = _3342 ^ _41097;
  wire _41099 = _2583 ^ _6213;
  wire _41100 = _41099 ^ _12525;
  wire _41101 = _41098 ^ _41100;
  wire _41102 = uncoded_block[344] ^ uncoded_block[349];
  wire _41103 = _11450 ^ _41102;
  wire _41104 = uncoded_block[358] ^ uncoded_block[365];
  wire _41105 = _13089 ^ _41104;
  wire _41106 = _41103 ^ _41105;
  wire _41107 = _15183 ^ _1035;
  wire _41108 = _41107 ^ _36376;
  wire _41109 = _41106 ^ _41108;
  wire _41110 = _41101 ^ _41109;
  wire _41111 = _41096 ^ _41110;
  wire _41112 = _2613 ^ _6879;
  wire _41113 = _1843 ^ _41112;
  wire _41114 = _3384 ^ _2623;
  wire _41115 = _5559 ^ _6244;
  wire _41116 = _41114 ^ _41115;
  wire _41117 = _41113 ^ _41116;
  wire _41118 = _4158 ^ _14159;
  wire _41119 = _4164 ^ _35576;
  wire _41120 = _41119 ^ _37610;
  wire _41121 = _41118 ^ _41120;
  wire _41122 = _41117 ^ _41121;
  wire _41123 = _17181 ^ _6259;
  wire _41124 = _12562 ^ _35583;
  wire _41125 = _41123 ^ _41124;
  wire _41126 = _4185 ^ _21059;
  wire _41127 = _1082 ^ _13132;
  wire _41128 = _41126 ^ _41127;
  wire _41129 = _41125 ^ _41128;
  wire _41130 = uncoded_block[484] ^ uncoded_block[488];
  wire _41131 = uncoded_block[489] ^ uncoded_block[497];
  wire _41132 = _41130 ^ _41131;
  wire _41133 = _1087 ^ _41132;
  wire _41134 = _4905 ^ _8700;
  wire _41135 = _6283 ^ _9298;
  wire _41136 = _41134 ^ _41135;
  wire _41137 = _41133 ^ _41136;
  wire _41138 = _41129 ^ _41137;
  wire _41139 = _41122 ^ _41138;
  wire _41140 = _41111 ^ _41139;
  wire _41141 = _41081 ^ _41140;
  wire _41142 = _19638 ^ _10947;
  wire _41143 = uncoded_block[529] ^ uncoded_block[536];
  wire _41144 = _41143 ^ _6293;
  wire _41145 = _41142 ^ _41144;
  wire _41146 = _1117 ^ _12592;
  wire _41147 = uncoded_block[550] ^ uncoded_block[554];
  wire _41148 = _41147 ^ _8724;
  wire _41149 = _41146 ^ _41148;
  wire _41150 = _41145 ^ _41149;
  wire _41151 = _6940 ^ _9319;
  wire _41152 = _41151 ^ _34804;
  wire _41153 = _4224 ^ _8731;
  wire _41154 = _11526 ^ _1138;
  wire _41155 = _41153 ^ _41154;
  wire _41156 = _41152 ^ _41155;
  wire _41157 = _41150 ^ _41156;
  wire _41158 = _3478 ^ _4234;
  wire _41159 = _4231 ^ _41158;
  wire _41160 = _8150 ^ _9869;
  wire _41161 = _41159 ^ _41160;
  wire _41162 = uncoded_block[605] ^ uncoded_block[610];
  wire _41163 = _41162 ^ _3492;
  wire _41164 = _41163 ^ _12613;
  wire _41165 = _1949 ^ _17734;
  wire _41166 = _41164 ^ _41165;
  wire _41167 = _41161 ^ _41166;
  wire _41168 = _41157 ^ _41167;
  wire _41169 = _3501 ^ _5661;
  wire _41170 = _26545 ^ _1163;
  wire _41171 = _41169 ^ _41170;
  wire _41172 = _296 ^ _2730;
  wire _41173 = _19181 ^ _9352;
  wire _41174 = _41172 ^ _41173;
  wire _41175 = _41171 ^ _41174;
  wire _41176 = _10990 ^ _311;
  wire _41177 = _41176 ^ _27810;
  wire _41178 = uncoded_block[686] ^ uncoded_block[693];
  wire _41179 = _26995 ^ _41178;
  wire _41180 = uncoded_block[694] ^ uncoded_block[698];
  wire _41181 = uncoded_block[700] ^ uncoded_block[704];
  wire _41182 = _41180 ^ _41181;
  wire _41183 = _41179 ^ _41182;
  wire _41184 = _41177 ^ _41183;
  wire _41185 = _41175 ^ _41184;
  wire _41186 = uncoded_block[707] ^ uncoded_block[713];
  wire _41187 = _3533 ^ _41186;
  wire _41188 = _41187 ^ _1196;
  wire _41189 = _1984 ^ _18259;
  wire _41190 = _5693 ^ _7002;
  wire _41191 = _41189 ^ _41190;
  wire _41192 = _41188 ^ _41191;
  wire _41193 = uncoded_block[734] ^ uncoded_block[736];
  wire _41194 = _41193 ^ _7005;
  wire _41195 = _23870 ^ _7006;
  wire _41196 = _41194 ^ _41195;
  wire _41197 = _1210 ^ _21605;
  wire _41198 = _20666 ^ _41197;
  wire _41199 = _41196 ^ _41198;
  wire _41200 = _41192 ^ _41199;
  wire _41201 = _41185 ^ _41200;
  wire _41202 = _41168 ^ _41201;
  wire _41203 = _7015 ^ _359;
  wire _41204 = _8781 ^ _364;
  wire _41205 = _41203 ^ _41204;
  wire _41206 = _5709 ^ _2791;
  wire _41207 = _5711 ^ _2014;
  wire _41208 = _41206 ^ _41207;
  wire _41209 = _41205 ^ _41208;
  wire _41210 = uncoded_block[781] ^ uncoded_block[786];
  wire _41211 = _368 ^ _41210;
  wire _41212 = _19709 ^ _6391;
  wire _41213 = _41211 ^ _41212;
  wire _41214 = _7029 ^ _7629;
  wire _41215 = _12127 ^ _1238;
  wire _41216 = _41214 ^ _41215;
  wire _41217 = _41213 ^ _41216;
  wire _41218 = _41209 ^ _41217;
  wire _41219 = _4324 ^ _3584;
  wire _41220 = _37697 ^ _41219;
  wire _41221 = _3587 ^ _12686;
  wire _41222 = _41221 ^ _35272;
  wire _41223 = _41220 ^ _41222;
  wire _41224 = _15330 ^ _37709;
  wire _41225 = _30254 ^ _41224;
  wire _41226 = _5071 ^ _5749;
  wire _41227 = _416 ^ _2835;
  wire _41228 = _41226 ^ _41227;
  wire _41229 = _41225 ^ _41228;
  wire _41230 = _41223 ^ _41229;
  wire _41231 = _41218 ^ _41230;
  wire _41232 = _11056 ^ _5082;
  wire _41233 = _35287 ^ _8250;
  wire _41234 = _41232 ^ _41233;
  wire _41235 = _5089 ^ _8254;
  wire _41236 = _41235 ^ _37326;
  wire _41237 = _41234 ^ _41236;
  wire _41238 = uncoded_block[918] ^ uncoded_block[923];
  wire _41239 = _7665 ^ _41238;
  wire _41240 = uncoded_block[925] ^ uncoded_block[931];
  wire _41241 = _41240 ^ _8262;
  wire _41242 = _41239 ^ _41241;
  wire _41243 = _9972 ^ _457;
  wire _41244 = _41242 ^ _41243;
  wire _41245 = _41237 ^ _41244;
  wire _41246 = _460 ^ _2869;
  wire _41247 = _8277 ^ _5783;
  wire _41248 = _41246 ^ _41247;
  wire _41249 = _12180 ^ _36515;
  wire _41250 = _32427 ^ _5792;
  wire _41251 = _41249 ^ _41250;
  wire _41252 = _41248 ^ _41251;
  wire _41253 = _18331 ^ _2884;
  wire _41254 = _23946 ^ _25757;
  wire _41255 = _41253 ^ _41254;
  wire _41256 = _41252 ^ _41255;
  wire _41257 = _41245 ^ _41256;
  wire _41258 = _41231 ^ _41257;
  wire _41259 = _41202 ^ _41258;
  wire _41260 = _41141 ^ _41259;
  wire _41261 = _487 ^ _8296;
  wire _41262 = _1331 ^ _2894;
  wire _41263 = _41261 ^ _41262;
  wire _41264 = _5137 ^ _495;
  wire _41265 = _12756 ^ _502;
  wire _41266 = _41264 ^ _41265;
  wire _41267 = _41263 ^ _41266;
  wire _41268 = _15387 ^ _22132;
  wire _41269 = _41268 ^ _31177;
  wire _41270 = _521 ^ _2142;
  wire _41271 = _17858 ^ _41270;
  wire _41272 = _41269 ^ _41271;
  wire _41273 = _41267 ^ _41272;
  wire _41274 = _7722 ^ _2924;
  wire _41275 = _17863 ^ _41274;
  wire _41276 = _20753 ^ _22149;
  wire _41277 = _18818 ^ _41276;
  wire _41278 = _41275 ^ _41277;
  wire _41279 = _1377 ^ _11139;
  wire _41280 = _8910 ^ _549;
  wire _41281 = _41279 ^ _41280;
  wire _41282 = _2938 ^ _10587;
  wire _41283 = _4452 ^ _41282;
  wire _41284 = _41281 ^ _41283;
  wire _41285 = _41278 ^ _41284;
  wire _41286 = _41273 ^ _41285;
  wire _41287 = _15894 ^ _4460;
  wire _41288 = uncoded_block[1137] ^ uncoded_block[1142];
  wire _41289 = _41288 ^ _2179;
  wire _41290 = _41287 ^ _41289;
  wire _41291 = _8932 ^ _8937;
  wire _41292 = uncoded_block[1159] ^ uncoded_block[1172];
  wire _41293 = _9500 ^ _41292;
  wire _41294 = _41291 ^ _41293;
  wire _41295 = _41290 ^ _41294;
  wire _41296 = uncoded_block[1173] ^ uncoded_block[1177];
  wire _41297 = _41296 ^ _27539;
  wire _41298 = _8944 ^ _9508;
  wire _41299 = _41297 ^ _41298;
  wire _41300 = _5203 ^ _24910;
  wire _41301 = _13886 ^ _13349;
  wire _41302 = _41300 ^ _41301;
  wire _41303 = _41299 ^ _41302;
  wire _41304 = _41295 ^ _41303;
  wire _41305 = _11171 ^ _1427;
  wire _41306 = _5213 ^ _606;
  wire _41307 = _41305 ^ _41306;
  wire _41308 = _4502 ^ _3769;
  wire _41309 = _3771 ^ _15441;
  wire _41310 = _41308 ^ _41309;
  wire _41311 = _41307 ^ _41310;
  wire _41312 = _10627 ^ _2995;
  wire _41313 = _6538 ^ _6543;
  wire _41314 = _41312 ^ _41313;
  wire _41315 = _6547 ^ _36994;
  wire _41316 = _41314 ^ _41315;
  wire _41317 = _41311 ^ _41316;
  wire _41318 = _41304 ^ _41317;
  wire _41319 = _41286 ^ _41318;
  wire _41320 = _7179 ^ _26718;
  wire _41321 = _3787 ^ _41320;
  wire _41322 = _6560 ^ _5913;
  wire _41323 = _27136 ^ _41322;
  wire _41324 = _41321 ^ _41323;
  wire _41325 = uncoded_block[1290] ^ uncoded_block[1294];
  wire _41326 = _41325 ^ _7799;
  wire _41327 = _648 ^ _6572;
  wire _41328 = _41326 ^ _41327;
  wire _41329 = _8407 ^ _1483;
  wire _41330 = _2262 ^ _3028;
  wire _41331 = _41329 ^ _41330;
  wire _41332 = _41328 ^ _41331;
  wire _41333 = _41324 ^ _41332;
  wire _41334 = _12289 ^ _40571;
  wire _41335 = _2277 ^ _7815;
  wire _41336 = _36183 ^ _41335;
  wire _41337 = _41334 ^ _41336;
  wire _41338 = _1498 ^ _664;
  wire _41339 = _5269 ^ _3042;
  wire _41340 = _41338 ^ _41339;
  wire _41341 = _33788 ^ _2284;
  wire _41342 = _39010 ^ _41341;
  wire _41343 = _41340 ^ _41342;
  wire _41344 = _41337 ^ _41343;
  wire _41345 = _41333 ^ _41344;
  wire _41346 = uncoded_block[1368] ^ uncoded_block[1376];
  wire _41347 = _41346 ^ _2290;
  wire _41348 = _16451 ^ _5950;
  wire _41349 = _41347 ^ _41348;
  wire _41350 = _5952 ^ _4572;
  wire _41351 = _41350 ^ _31694;
  wire _41352 = _41349 ^ _41351;
  wire _41353 = _13420 ^ _17461;
  wire _41354 = _38217 ^ _709;
  wire _41355 = _41353 ^ _41354;
  wire _41356 = _10684 ^ _1533;
  wire _41357 = _15982 ^ _2319;
  wire _41358 = _41356 ^ _41357;
  wire _41359 = _41355 ^ _41358;
  wire _41360 = _41352 ^ _41359;
  wire _41361 = _11246 ^ _2329;
  wire _41362 = _2335 ^ _9602;
  wire _41363 = _41361 ^ _41362;
  wire _41364 = uncoded_block[1471] ^ uncoded_block[1479];
  wire _41365 = _7247 ^ _41364;
  wire _41366 = _12342 ^ _7861;
  wire _41367 = _41365 ^ _41366;
  wire _41368 = _41363 ^ _41367;
  wire _41369 = uncoded_block[1492] ^ uncoded_block[1495];
  wire _41370 = _7251 ^ _41369;
  wire _41371 = uncoded_block[1498] ^ uncoded_block[1508];
  wire _41372 = _41371 ^ _750;
  wire _41373 = _41370 ^ _41372;
  wire _41374 = _19429 ^ _14488;
  wire _41375 = _754 ^ _3122;
  wire _41376 = _41374 ^ _41375;
  wire _41377 = _41373 ^ _41376;
  wire _41378 = _41368 ^ _41377;
  wire _41379 = _41360 ^ _41378;
  wire _41380 = _41345 ^ _41379;
  wire _41381 = _41319 ^ _41380;
  wire _41382 = _22266 ^ _6006;
  wire _41383 = _27626 ^ _16995;
  wire _41384 = _41382 ^ _41383;
  wire _41385 = _13472 ^ _6657;
  wire _41386 = _41385 ^ _16509;
  wire _41387 = _41384 ^ _41386;
  wire _41388 = _3139 ^ _777;
  wire _41389 = _4647 ^ _782;
  wire _41390 = _41388 ^ _41389;
  wire _41391 = uncoded_block[1578] ^ uncoded_block[1586];
  wire _41392 = _41391 ^ _21827;
  wire _41393 = _41392 ^ _15037;
  wire _41394 = _41390 ^ _41393;
  wire _41395 = _41387 ^ _41394;
  wire _41396 = _14000 ^ _5380;
  wire _41397 = _3157 ^ _10181;
  wire _41398 = _41396 ^ _41397;
  wire _41399 = _7298 ^ _3941;
  wire _41400 = _807 ^ _11307;
  wire _41401 = _41399 ^ _41400;
  wire _41402 = _41398 ^ _41401;
  wire _41403 = _12383 ^ _4673;
  wire _41404 = _16530 ^ _41403;
  wire _41405 = _2412 ^ _3953;
  wire _41406 = _820 ^ _822;
  wire _41407 = _41405 ^ _41406;
  wire _41408 = _41404 ^ _41407;
  wire _41409 = _41402 ^ _41408;
  wire _41410 = _41395 ^ _41409;
  wire _41411 = _6055 ^ _1654;
  wire _41412 = uncoded_block[1668] ^ uncoded_block[1672];
  wire _41413 = _7319 ^ _41412;
  wire _41414 = _41411 ^ _41413;
  wire _41415 = _5401 ^ _11321;
  wire _41416 = uncoded_block[1684] ^ uncoded_block[1689];
  wire _41417 = _17040 ^ _41416;
  wire _41418 = _41415 ^ _41417;
  wire _41419 = _41414 ^ _41418;
  wire _41420 = _7331 ^ _14024;
  wire _41421 = _1669 ^ _3973;
  wire _41422 = _41420 ^ _41421;
  wire _41423 = uncoded_block[1702] ^ uncoded_block[1711];
  wire _41424 = _41423 ^ _852;
  wire _41425 = _7944 ^ uncoded_block[1717];
  wire _41426 = _41424 ^ _41425;
  wire _41427 = _41422 ^ _41426;
  wire _41428 = _41419 ^ _41427;
  wire _41429 = _41410 ^ _41428;
  wire _41430 = _41381 ^ _41429;
  wire _41431 = _41260 ^ _41430;
  wire _41432 = _866 ^ _18057;
  wire _41433 = _41432 ^ _18059;
  wire _41434 = uncoded_block[21] ^ uncoded_block[26];
  wire _41435 = _10226 ^ _41434;
  wire _41436 = _19965 ^ _18;
  wire _41437 = _41435 ^ _41436;
  wire _41438 = _41433 ^ _41437;
  wire _41439 = _19 ^ _12425;
  wire _41440 = _6099 ^ _4726;
  wire _41441 = _41439 ^ _41440;
  wire _41442 = _2472 ^ _894;
  wire _41443 = _34 ^ _26393;
  wire _41444 = _41442 ^ _41443;
  wire _41445 = _41441 ^ _41444;
  wire _41446 = _41438 ^ _41445;
  wire _41447 = _14060 ^ _4735;
  wire _41448 = _2483 ^ _14065;
  wire _41449 = _41447 ^ _41448;
  wire _41450 = _8567 ^ _3249;
  wire _41451 = _7377 ^ _1721;
  wire _41452 = _41450 ^ _41451;
  wire _41453 = _41449 ^ _41452;
  wire _41454 = uncoded_block[107] ^ uncoded_block[111];
  wire _41455 = _41454 ^ _6763;
  wire _41456 = uncoded_block[114] ^ uncoded_block[118];
  wire _41457 = _41456 ^ _12451;
  wire _41458 = _41455 ^ _41457;
  wire _41459 = _11374 ^ _1735;
  wire _41460 = _41459 ^ _11917;
  wire _41461 = _41458 ^ _41460;
  wire _41462 = _41453 ^ _41461;
  wire _41463 = _41446 ^ _41462;
  wire _41464 = _4760 ^ _16600;
  wire _41465 = _4046 ^ _14082;
  wire _41466 = _41464 ^ _41465;
  wire _41467 = _33487 ^ _79;
  wire _41468 = _36324 ^ _41467;
  wire _41469 = _41466 ^ _41468;
  wire _41470 = _5473 ^ _940;
  wire _41471 = _2525 ^ _4062;
  wire _41472 = _41470 ^ _41471;
  wire _41473 = uncoded_block[189] ^ uncoded_block[192];
  wire _41474 = uncoded_block[193] ^ uncoded_block[202];
  wire _41475 = _41473 ^ _41474;
  wire _41476 = _4070 ^ _4780;
  wire _41477 = _41475 ^ _41476;
  wire _41478 = _41472 ^ _41477;
  wire _41479 = _41469 ^ _41478;
  wire _41480 = _4071 ^ _1767;
  wire _41481 = _41480 ^ _8607;
  wire _41482 = uncoded_block[227] ^ uncoded_block[234];
  wire _41483 = _35912 ^ _41482;
  wire _41484 = _18125 ^ _9756;
  wire _41485 = _41483 ^ _41484;
  wire _41486 = _41481 ^ _41485;
  wire _41487 = _11952 ^ _14116;
  wire _41488 = _41487 ^ _35149;
  wire _41489 = _8620 ^ _25108;
  wire _41490 = _41489 ^ _26443;
  wire _41491 = _41488 ^ _41490;
  wire _41492 = _41486 ^ _41491;
  wire _41493 = _41479 ^ _41492;
  wire _41494 = _41463 ^ _41493;
  wire _41495 = _4102 ^ _5513;
  wire _41496 = _41495 ^ _37967;
  wire _41497 = _2577 ^ _7453;
  wire _41498 = _18139 ^ _41497;
  wire _41499 = _41496 ^ _41498;
  wire _41500 = uncoded_block[311] ^ uncoded_block[316];
  wire _41501 = _21017 ^ _41500;
  wire _41502 = uncoded_block[322] ^ uncoded_block[325];
  wire _41503 = _6850 ^ _41502;
  wire _41504 = _41501 ^ _41503;
  wire _41505 = _1014 ^ _11983;
  wire _41506 = _1821 ^ _8646;
  wire _41507 = _41505 ^ _41506;
  wire _41508 = _41504 ^ _41507;
  wire _41509 = _41499 ^ _41508;
  wire _41510 = _4844 ^ _5541;
  wire _41511 = _17650 ^ _41510;
  wire _41512 = _36782 ^ _2602;
  wire _41513 = uncoded_block[365] ^ uncoded_block[369];
  wire _41514 = _6864 ^ _41513;
  wire _41515 = _41512 ^ _41514;
  wire _41516 = _41511 ^ _41515;
  wire _41517 = _29257 ^ _10899;
  wire _41518 = _41517 ^ _1843;
  wire _41519 = _3380 ^ _12541;
  wire _41520 = _1847 ^ _2622;
  wire _41521 = _41519 ^ _41520;
  wire _41522 = _41518 ^ _41521;
  wire _41523 = _41516 ^ _41522;
  wire _41524 = _41509 ^ _41523;
  wire _41525 = uncoded_block[403] ^ uncoded_block[406];
  wire _41526 = _41525 ^ _27341;
  wire _41527 = _41526 ^ _26487;
  wire _41528 = _35963 ^ _28104;
  wire _41529 = _41527 ^ _41528;
  wire _41530 = _10356 ^ _4176;
  wire _41531 = _28489 ^ _41530;
  wire _41532 = _1070 ^ _212;
  wire _41533 = _41532 ^ _39202;
  wire _41534 = _41531 ^ _41533;
  wire _41535 = _41529 ^ _41534;
  wire _41536 = _32711 ^ _1880;
  wire _41537 = uncoded_block[474] ^ uncoded_block[478];
  wire _41538 = _41537 ^ _1085;
  wire _41539 = _41538 ^ _39593;
  wire _41540 = _41536 ^ _41539;
  wire _41541 = _5600 ^ _10937;
  wire _41542 = _6919 ^ _21067;
  wire _41543 = _41541 ^ _41542;
  wire _41544 = _7521 ^ _12034;
  wire _41545 = _41544 ^ _35989;
  wire _41546 = _41543 ^ _41545;
  wire _41547 = _41540 ^ _41546;
  wire _41548 = _41535 ^ _41547;
  wire _41549 = _41524 ^ _41548;
  wire _41550 = _41494 ^ _41549;
  wire _41551 = _22447 ^ _40002;
  wire _41552 = _19146 ^ _24278;
  wire _41553 = _41551 ^ _41552;
  wire _41554 = uncoded_block[543] ^ uncoded_block[547];
  wire _41555 = _1115 ^ _41554;
  wire _41556 = _1912 ^ _25182;
  wire _41557 = _41555 ^ _41556;
  wire _41558 = _1126 ^ _7550;
  wire _41559 = _36418 ^ _41558;
  wire _41560 = _41557 ^ _41559;
  wire _41561 = _41553 ^ _41560;
  wire _41562 = _7551 ^ _10399;
  wire _41563 = _4229 ^ _1933;
  wire _41564 = _41562 ^ _41563;
  wire _41565 = _4233 ^ _1938;
  wire _41566 = _17721 ^ _8736;
  wire _41567 = _41565 ^ _41566;
  wire _41568 = _41564 ^ _41567;
  wire _41569 = _3489 ^ _277;
  wire _41570 = uncoded_block[608] ^ uncoded_block[612];
  wire _41571 = _41570 ^ _7567;
  wire _41572 = _41569 ^ _41571;
  wire _41573 = _1946 ^ _14224;
  wire _41574 = _41573 ^ _22026;
  wire _41575 = _41572 ^ _41574;
  wire _41576 = _41568 ^ _41575;
  wire _41577 = _41561 ^ _41576;
  wire _41578 = _6969 ^ _2730;
  wire _41579 = _40417 ^ _41578;
  wire _41580 = _6344 ^ _10990;
  wire _41581 = _32755 ^ _41580;
  wire _41582 = _41579 ^ _41581;
  wire _41583 = _1177 ^ _1181;
  wire _41584 = uncoded_block[687] ^ uncoded_block[691];
  wire _41585 = _12636 ^ _41584;
  wire _41586 = _41583 ^ _41585;
  wire _41587 = _4272 ^ _41180;
  wire _41588 = _11562 ^ _11564;
  wire _41589 = _41587 ^ _41588;
  wire _41590 = _41586 ^ _41589;
  wire _41591 = _41582 ^ _41590;
  wire _41592 = _14772 ^ _17763;
  wire _41593 = _5005 ^ _352;
  wire _41594 = _15301 ^ _1210;
  wire _41595 = _41593 ^ _41594;
  wire _41596 = _41592 ^ _41595;
  wire _41597 = _12663 ^ _13213;
  wire _41598 = _364 ^ _13215;
  wire _41599 = _41597 ^ _41598;
  wire _41600 = _9382 ^ _13219;
  wire _41601 = _12668 ^ _41600;
  wire _41602 = _41599 ^ _41601;
  wire _41603 = _41596 ^ _41602;
  wire _41604 = _41591 ^ _41603;
  wire _41605 = _41577 ^ _41604;
  wire _41606 = _13221 ^ _27021;
  wire _41607 = uncoded_block[790] ^ uncoded_block[795];
  wire _41608 = _41607 ^ _382;
  wire _41609 = _385 ^ _22071;
  wire _41610 = _41608 ^ _41609;
  wire _41611 = _41606 ^ _41610;
  wire _41612 = uncoded_block[806] ^ uncoded_block[812];
  wire _41613 = _41612 ^ _10485;
  wire _41614 = _1241 ^ _15320;
  wire _41615 = _41613 ^ _41614;
  wire _41616 = _1247 ^ _4331;
  wire _41617 = _2035 ^ _7640;
  wire _41618 = _41616 ^ _41617;
  wire _41619 = _41615 ^ _41618;
  wire _41620 = _41611 ^ _41619;
  wire _41621 = uncoded_block[845] ^ uncoded_block[849];
  wire _41622 = _41621 ^ _14814;
  wire _41623 = _41622 ^ _20693;
  wire _41624 = _9949 ^ _11618;
  wire _41625 = _6415 ^ _1269;
  wire _41626 = _41624 ^ _41625;
  wire _41627 = _41623 ^ _41626;
  wire _41628 = uncoded_block[876] ^ uncoded_block[880];
  wire _41629 = _41628 ^ _2061;
  wire _41630 = uncoded_block[897] ^ uncoded_block[905];
  wire _41631 = _1277 ^ _41630;
  wire _41632 = _41629 ^ _41631;
  wire _41633 = _9421 ^ _9424;
  wire _41634 = _41633 ^ _17819;
  wire _41635 = _41632 ^ _41634;
  wire _41636 = _41627 ^ _41635;
  wire _41637 = _41620 ^ _41636;
  wire _41638 = _439 ^ _31995;
  wire _41639 = _41638 ^ _31582;
  wire _41640 = _455 ^ _3643;
  wire _41641 = _40096 ^ _41640;
  wire _41642 = _41639 ^ _41641;
  wire _41643 = _4385 ^ _14844;
  wire _41644 = _34095 ^ _41643;
  wire _41645 = _9981 ^ _36515;
  wire _41646 = _5112 ^ _4391;
  wire _41647 = _41645 ^ _41646;
  wire _41648 = _41644 ^ _41647;
  wire _41649 = _41642 ^ _41648;
  wire _41650 = _6451 ^ _23938;
  wire _41651 = _9442 ^ _41650;
  wire _41652 = _2882 ^ _8293;
  wire _41653 = _5798 ^ _3666;
  wire _41654 = _41652 ^ _41653;
  wire _41655 = _41651 ^ _41654;
  wire _41656 = _2890 ^ _11663;
  wire _41657 = _41656 ^ _21208;
  wire _41658 = _495 ^ _9459;
  wire _41659 = _2908 ^ _6475;
  wire _41660 = _41658 ^ _41659;
  wire _41661 = _41657 ^ _41660;
  wire _41662 = _41655 ^ _41661;
  wire _41663 = _41649 ^ _41662;
  wire _41664 = _41637 ^ _41663;
  wire _41665 = _41605 ^ _41664;
  wire _41666 = _41550 ^ _41665;
  wire _41667 = _23498 ^ _515;
  wire _41668 = uncoded_block[1054] ^ uncoded_block[1060];
  wire _41669 = _13844 ^ _41668;
  wire _41670 = _41667 ^ _41669;
  wire _41671 = _20749 ^ _5829;
  wire _41672 = _41670 ^ _41671;
  wire _41673 = uncoded_block[1073] ^ uncoded_block[1079];
  wire _41674 = _41673 ^ _530;
  wire _41675 = _1373 ^ _4440;
  wire _41676 = _41674 ^ _41675;
  wire _41677 = _11137 ^ _16878;
  wire _41678 = _8910 ^ _2161;
  wire _41679 = _41677 ^ _41678;
  wire _41680 = _41676 ^ _41679;
  wire _41681 = _41672 ^ _41680;
  wire _41682 = _4450 ^ _7133;
  wire _41683 = _29427 ^ _13327;
  wire _41684 = _41682 ^ _41683;
  wire _41685 = _14380 ^ _8346;
  wire _41686 = _9495 ^ _41685;
  wire _41687 = _41684 ^ _41686;
  wire _41688 = _18377 ^ _8932;
  wire _41689 = _41688 ^ _20271;
  wire _41690 = uncoded_block[1156] ^ uncoded_block[1161];
  wire _41691 = _41690 ^ _2964;
  wire _41692 = _41691 ^ _4477;
  wire _41693 = _41689 ^ _41692;
  wire _41694 = _41687 ^ _41693;
  wire _41695 = _41681 ^ _41694;
  wire _41696 = uncoded_block[1169] ^ uncoded_block[1176];
  wire _41697 = uncoded_block[1177] ^ uncoded_block[1188];
  wire _41698 = _41696 ^ _41697;
  wire _41699 = _41698 ^ _10613;
  wire _41700 = _1421 ^ _1424;
  wire _41701 = _41700 ^ _28297;
  wire _41702 = _41699 ^ _41701;
  wire _41703 = _2217 ^ _27911;
  wire _41704 = _41703 ^ _32074;
  wire _41705 = _7774 ^ _2995;
  wire _41706 = _8959 ^ _41705;
  wire _41707 = _41704 ^ _41706;
  wire _41708 = _41702 ^ _41707;
  wire _41709 = _6543 ^ _32082;
  wire _41710 = _41709 ^ _6549;
  wire _41711 = _2239 ^ _1459;
  wire _41712 = _3010 ^ _15455;
  wire _41713 = _41711 ^ _41712;
  wire _41714 = _41710 ^ _41713;
  wire _41715 = _4529 ^ _39382;
  wire _41716 = _14939 ^ _22665;
  wire _41717 = _41715 ^ _41716;
  wire _41718 = _3807 ^ _1480;
  wire _41719 = uncoded_block[1318] ^ uncoded_block[1323];
  wire _41720 = _20314 ^ _41719;
  wire _41721 = _41718 ^ _41720;
  wire _41722 = _41717 ^ _41721;
  wire _41723 = _41714 ^ _41722;
  wire _41724 = _41708 ^ _41723;
  wire _41725 = _41695 ^ _41724;
  wire _41726 = _1489 ^ _8998;
  wire _41727 = _4551 ^ _13399;
  wire _41728 = _41726 ^ _41727;
  wire _41729 = _5262 ^ _14442;
  wire _41730 = _33363 ^ _12857;
  wire _41731 = _41729 ^ _41730;
  wire _41732 = _41728 ^ _41731;
  wire _41733 = _4559 ^ _1504;
  wire _41734 = _41733 ^ _3048;
  wire _41735 = _3052 ^ _9573;
  wire _41736 = _5285 ^ _15483;
  wire _41737 = _41735 ^ _41736;
  wire _41738 = _41734 ^ _41737;
  wire _41739 = _41732 ^ _41738;
  wire _41740 = _19864 ^ _13938;
  wire _41741 = _1517 ^ _2300;
  wire _41742 = _41740 ^ _41741;
  wire _41743 = _5957 ^ _10117;
  wire _41744 = _41743 ^ _36628;
  wire _41745 = _41742 ^ _41744;
  wire _41746 = uncoded_block[1422] ^ uncoded_block[1431];
  wire _41747 = uncoded_block[1432] ^ uncoded_block[1438];
  wire _41748 = _41746 ^ _41747;
  wire _41749 = _24065 ^ _11246;
  wire _41750 = _41748 ^ _41749;
  wire _41751 = _2328 ^ _22252;
  wire _41752 = _3870 ^ _20855;
  wire _41753 = _41751 ^ _41752;
  wire _41754 = _41750 ^ _41753;
  wire _41755 = _41745 ^ _41754;
  wire _41756 = _41739 ^ _41755;
  wire _41757 = uncoded_block[1474] ^ uncoded_block[1479];
  wire _41758 = _5983 ^ _41757;
  wire _41759 = _14479 ^ _16981;
  wire _41760 = _41758 ^ _41759;
  wire _41761 = _12896 ^ _3890;
  wire _41762 = uncoded_block[1501] ^ uncoded_block[1504];
  wire _41763 = _6634 ^ _41762;
  wire _41764 = _41761 ^ _41763;
  wire _41765 = _41760 ^ _41764;
  wire _41766 = _11264 ^ _750;
  wire _41767 = _41766 ^ _14489;
  wire _41768 = uncoded_block[1521] ^ uncoded_block[1528];
  wire _41769 = _754 ^ _41768;
  wire _41770 = _5344 ^ _6005;
  wire _41771 = _41769 ^ _41770;
  wire _41772 = _41767 ^ _41771;
  wire _41773 = _41765 ^ _41772;
  wire _41774 = _7883 ^ _3912;
  wire _41775 = _32973 ^ _41774;
  wire _41776 = _25001 ^ _1596;
  wire _41777 = _13991 ^ _29986;
  wire _41778 = _41776 ^ _41777;
  wire _41779 = _41775 ^ _41778;
  wire _41780 = _21361 ^ _13479;
  wire _41781 = _41780 ^ _7899;
  wire _41782 = _4653 ^ _11292;
  wire _41783 = _41782 ^ _32168;
  wire _41784 = _41781 ^ _41783;
  wire _41785 = _41779 ^ _41784;
  wire _41786 = _41773 ^ _41785;
  wire _41787 = _41756 ^ _41786;
  wire _41788 = _41725 ^ _41787;
  wire _41789 = _10742 ^ _31740;
  wire _41790 = _41789 ^ _31326;
  wire _41791 = _3160 ^ _14006;
  wire _41792 = _41791 ^ _17524;
  wire _41793 = _41790 ^ _41792;
  wire _41794 = _7914 ^ _10754;
  wire _41795 = _41794 ^ _9104;
  wire _41796 = _4673 ^ _9661;
  wire _41797 = _9662 ^ _10761;
  wire _41798 = _41796 ^ _41797;
  wire _41799 = _41795 ^ _41798;
  wire _41800 = _41793 ^ _41799;
  wire _41801 = uncoded_block[1661] ^ uncoded_block[1665];
  wire _41802 = _41801 ^ _10200;
  wire _41803 = _41009 ^ _20427;
  wire _41804 = _41802 ^ _41803;
  wire _41805 = _17040 ^ _10205;
  wire _41806 = _18041 ^ _5409;
  wire _41807 = _41805 ^ _41806;
  wire _41808 = _41804 ^ _41807;
  wire _41809 = _39476 ^ _7939;
  wire _41810 = _3980 ^ _3200;
  wire _41811 = _855 ^ _12976;
  wire _41812 = _41810 ^ _41811;
  wire _41813 = _41809 ^ _41812;
  wire _41814 = _41808 ^ _41813;
  wire _41815 = _41800 ^ _41814;
  wire _41816 = _41815 ^ uncoded_block[1722];
  wire _41817 = _41788 ^ _41816;
  wire _41818 = _41666 ^ _41817;
  wire _41819 = _21407 ^ _3993;
  wire _41820 = _41819 ^ _7349;
  wire _41821 = _4713 ^ _7351;
  wire _41822 = _41821 ^ _37113;
  wire _41823 = _41820 ^ _41822;
  wire _41824 = _11890 ^ _13543;
  wire _41825 = _18549 ^ _7965;
  wire _41826 = _41824 ^ _41825;
  wire _41827 = _3232 ^ _23255;
  wire _41828 = _33039 ^ _41827;
  wire _41829 = _41826 ^ _41828;
  wire _41830 = _41823 ^ _41829;
  wire _41831 = _7969 ^ _6742;
  wire _41832 = _41831 ^ _9706;
  wire _41833 = _33467 ^ _22805;
  wire _41834 = _14586 ^ _42;
  wire _41835 = _41833 ^ _41834;
  wire _41836 = _41832 ^ _41835;
  wire _41837 = _6115 ^ _12443;
  wire _41838 = _4028 ^ _1721;
  wire _41839 = _41837 ^ _41838;
  wire _41840 = _6122 ^ _53;
  wire _41841 = _54 ^ _10819;
  wire _41842 = _41840 ^ _41841;
  wire _41843 = _41839 ^ _41842;
  wire _41844 = _41836 ^ _41843;
  wire _41845 = _41830 ^ _41844;
  wire _41846 = uncoded_block[124] ^ uncoded_block[128];
  wire _41847 = _41846 ^ _923;
  wire _41848 = _41847 ^ _17594;
  wire _41849 = _1736 ^ _6776;
  wire _41850 = uncoded_block[152] ^ uncoded_block[159];
  wire _41851 = _70 ^ _41850;
  wire _41852 = _41849 ^ _41851;
  wire _41853 = _41848 ^ _41852;
  wire _41854 = _78 ^ _29624;
  wire _41855 = uncoded_block[176] ^ uncoded_block[180];
  wire _41856 = _8591 ^ _41855;
  wire _41857 = _41854 ^ _41856;
  wire _41858 = _7409 ^ _3283;
  wire _41859 = _41858 ^ _35529;
  wire _41860 = _41857 ^ _41859;
  wire _41861 = _41853 ^ _41860;
  wire _41862 = _97 ^ _3296;
  wire _41863 = _22839 ^ _41862;
  wire _41864 = _2545 ^ _41482;
  wire _41865 = _19055 ^ _41864;
  wire _41866 = _41863 ^ _41865;
  wire _41867 = _22852 ^ _7433;
  wire _41868 = _1786 ^ _4096;
  wire _41869 = _26000 ^ _33099;
  wire _41870 = _41868 ^ _41869;
  wire _41871 = _41867 ^ _41870;
  wire _41872 = _41866 ^ _41871;
  wire _41873 = _41861 ^ _41872;
  wire _41874 = _41845 ^ _41873;
  wire _41875 = _4102 ^ _2568;
  wire _41876 = uncoded_block[278] ^ uncoded_block[281];
  wire _41877 = _41876 ^ _4105;
  wire _41878 = _41875 ^ _41877;
  wire _41879 = _20038 ^ _10312;
  wire _41880 = _11969 ^ _41879;
  wire _41881 = _41878 ^ _41880;
  wire _41882 = _14133 ^ _1000;
  wire _41883 = _1813 ^ _4832;
  wire _41884 = _41882 ^ _41883;
  wire _41885 = uncoded_block[323] ^ uncoded_block[328];
  wire _41886 = _41885 ^ _2586;
  wire _41887 = uncoded_block[336] ^ uncoded_block[340];
  wire _41888 = _2587 ^ _41887;
  wire _41889 = _41886 ^ _41888;
  wire _41890 = _41884 ^ _41889;
  wire _41891 = _41881 ^ _41890;
  wire _41892 = _159 ^ _5541;
  wire _41893 = _41892 ^ _22878;
  wire _41894 = _41104 ^ _169;
  wire _41895 = _29257 ^ _7474;
  wire _41896 = _41894 ^ _41895;
  wire _41897 = _41893 ^ _41896;
  wire _41898 = _7476 ^ _1039;
  wire _41899 = _41898 ^ _8662;
  wire _41900 = _19606 ^ _3392;
  wire _41901 = _41899 ^ _41900;
  wire _41902 = _41897 ^ _41901;
  wire _41903 = _41891 ^ _41902;
  wire _41904 = _4163 ^ _6889;
  wire _41905 = _17673 ^ _41904;
  wire _41906 = _6255 ^ _13122;
  wire _41907 = _15199 ^ _41906;
  wire _41908 = _41905 ^ _41907;
  wire _41909 = uncoded_block[452] ^ uncoded_block[455];
  wire _41910 = _1866 ^ _41909;
  wire _41911 = _41910 ^ _18185;
  wire _41912 = _6906 ^ _2657;
  wire _41913 = _36805 ^ _41912;
  wire _41914 = _41911 ^ _41913;
  wire _41915 = _41908 ^ _41914;
  wire _41916 = _14180 ^ _7517;
  wire _41917 = uncoded_block[492] ^ uncoded_block[502];
  wire _41918 = _41917 ^ _12034;
  wire _41919 = _7531 ^ _20598;
  wire _41920 = _41918 ^ _41919;
  wire _41921 = _41916 ^ _41920;
  wire _41922 = _1901 ^ _16215;
  wire _41923 = _4211 ^ _41922;
  wire _41924 = _6932 ^ _24279;
  wire _41925 = _8132 ^ _41554;
  wire _41926 = _41924 ^ _41925;
  wire _41927 = _41923 ^ _41926;
  wire _41928 = _41921 ^ _41927;
  wire _41929 = _41915 ^ _41928;
  wire _41930 = _41903 ^ _41929;
  wire _41931 = _41874 ^ _41930;
  wire _41932 = uncoded_block[556] ^ uncoded_block[561];
  wire _41933 = _1912 ^ _41932;
  wire _41934 = _32327 ^ _7550;
  wire _41935 = _41933 ^ _41934;
  wire _41936 = _262 ^ _11526;
  wire _41937 = _26092 ^ _41936;
  wire _41938 = _41935 ^ _41937;
  wire _41939 = _6947 ^ _9325;
  wire _41940 = _41939 ^ _14734;
  wire _41941 = uncoded_block[597] ^ uncoded_block[601];
  wire _41942 = _20618 ^ _41941;
  wire _41943 = _2709 ^ _1146;
  wire _41944 = _41942 ^ _41943;
  wire _41945 = _41940 ^ _41944;
  wire _41946 = _41938 ^ _41945;
  wire _41947 = _20626 ^ _7564;
  wire _41948 = uncoded_block[616] ^ uncoded_block[622];
  wire _41949 = _41948 ^ _2720;
  wire _41950 = _41947 ^ _41949;
  wire _41951 = _1953 ^ _36435;
  wire _41952 = _6336 ^ _2729;
  wire _41953 = _41951 ^ _41952;
  wire _41954 = _41950 ^ _41953;
  wire _41955 = uncoded_block[646] ^ uncoded_block[652];
  wire _41956 = _41955 ^ _4975;
  wire _41957 = uncoded_block[659] ^ uncoded_block[663];
  wire _41958 = uncoded_block[668] ^ uncoded_block[676];
  wire _41959 = _41957 ^ _41958;
  wire _41960 = _41956 ^ _41959;
  wire _41961 = _1968 ^ _1971;
  wire _41962 = _41961 ^ _26555;
  wire _41963 = _41960 ^ _41962;
  wire _41964 = _41954 ^ _41963;
  wire _41965 = _41946 ^ _41964;
  wire _41966 = _4271 ^ _6357;
  wire _41967 = _2755 ^ _19195;
  wire _41968 = _41966 ^ _41967;
  wire _41969 = _11563 ^ _18256;
  wire _41970 = _41968 ^ _41969;
  wire _41971 = _8192 ^ _30645;
  wire _41972 = _41971 ^ _3545;
  wire _41973 = _1202 ^ _7605;
  wire _41974 = _20156 ^ _1998;
  wire _41975 = _41973 ^ _41974;
  wire _41976 = _41972 ^ _41975;
  wire _41977 = _41970 ^ _41976;
  wire _41978 = _8209 ^ _21605;
  wire _41979 = _41978 ^ _13214;
  wire _41980 = _8213 ^ _7021;
  wire _41981 = _25687 ^ _41980;
  wire _41982 = _41979 ^ _41981;
  wire _41983 = _2794 ^ _3570;
  wire _41984 = _41983 ^ _36881;
  wire _41985 = _8223 ^ _7029;
  wire _41986 = _41985 ^ _11595;
  wire _41987 = _41984 ^ _41986;
  wire _41988 = _41982 ^ _41987;
  wire _41989 = _41977 ^ _41988;
  wire _41990 = _41965 ^ _41989;
  wire _41991 = _10483 ^ _5046;
  wire _41992 = _27843 ^ _14291;
  wire _41993 = _41991 ^ _41992;
  wire _41994 = _3590 ^ _4331;
  wire _41995 = _41994 ^ _17296;
  wire _41996 = _41993 ^ _41995;
  wire _41997 = _5057 ^ _4339;
  wire _41998 = _41997 ^ _11611;
  wire _41999 = _12146 ^ _29368;
  wire _42000 = _5066 ^ _6412;
  wire _42001 = _41999 ^ _42000;
  wire _42002 = _41998 ^ _42001;
  wire _42003 = _41996 ^ _42002;
  wire _42004 = _1266 ^ _416;
  wire _42005 = _2831 ^ _8820;
  wire _42006 = _42004 ^ _42005;
  wire _42007 = _35678 ^ _19735;
  wire _42008 = _42007 ^ _1282;
  wire _42009 = _42006 ^ _42008;
  wire _42010 = _1284 ^ _19252;
  wire _42011 = _42010 ^ _13256;
  wire _42012 = _3632 ^ _35296;
  wire _42013 = _42012 ^ _2080;
  wire _42014 = _42011 ^ _42013;
  wire _42015 = _42009 ^ _42014;
  wire _42016 = _42003 ^ _42015;
  wire _42017 = _18321 ^ _2087;
  wire _42018 = _34496 ^ _2090;
  wire _42019 = _1308 ^ _7088;
  wire _42020 = _42018 ^ _42019;
  wire _42021 = _42017 ^ _42020;
  wire _42022 = uncoded_block[971] ^ uncoded_block[977];
  wire _42023 = _42022 ^ _11092;
  wire _42024 = _476 ^ _5118;
  wire _42025 = _42023 ^ _42024;
  wire _42026 = _16338 ^ _25289;
  wire _42027 = uncoded_block[996] ^ uncoded_block[1002];
  wire _42028 = _42027 ^ _6459;
  wire _42029 = _42026 ^ _42028;
  wire _42030 = _42025 ^ _42029;
  wire _42031 = _42021 ^ _42030;
  wire _42032 = _4409 ^ _2117;
  wire _42033 = _9996 ^ _8871;
  wire _42034 = _42032 ^ _42033;
  wire _42035 = _35320 ^ _5810;
  wire _42036 = _1346 ^ _2130;
  wire _42037 = _42035 ^ _42036;
  wire _42038 = _42034 ^ _42037;
  wire _42039 = uncoded_block[1047] ^ uncoded_block[1051];
  wire _42040 = _2133 ^ _42039;
  wire _42041 = _12762 ^ _4430;
  wire _42042 = _42040 ^ _42041;
  wire _42043 = _519 ^ _6483;
  wire _42044 = uncoded_block[1061] ^ uncoded_block[1066];
  wire _42045 = _42044 ^ _8892;
  wire _42046 = _42043 ^ _42045;
  wire _42047 = _42042 ^ _42046;
  wire _42048 = _42038 ^ _42047;
  wire _42049 = _42031 ^ _42048;
  wire _42050 = _42016 ^ _42049;
  wire _42051 = _41990 ^ _42050;
  wire _42052 = _41931 ^ _42051;
  wire _42053 = _12770 ^ _5162;
  wire _42054 = uncoded_block[1081] ^ uncoded_block[1085];
  wire _42055 = _42054 ^ _3696;
  wire _42056 = _42053 ^ _42055;
  wire _42057 = _5843 ^ _543;
  wire _42058 = _39339 ^ _42057;
  wire _42059 = _42056 ^ _42058;
  wire _42060 = _546 ^ _550;
  wire _42061 = _1386 ^ _30326;
  wire _42062 = _42060 ^ _42061;
  wire _42063 = _2942 ^ _33312;
  wire _42064 = _6499 ^ _8929;
  wire _42065 = _42063 ^ _42064;
  wire _42066 = _42062 ^ _42065;
  wire _42067 = _42059 ^ _42066;
  wire _42068 = _5862 ^ _8933;
  wire _42069 = _2954 ^ _42068;
  wire _42070 = _3727 ^ _5190;
  wire _42071 = _3733 ^ _3736;
  wire _42072 = _42070 ^ _42071;
  wire _42073 = _42069 ^ _42072;
  wire _42074 = _13338 ^ _14901;
  wire _42075 = _13882 ^ _3749;
  wire _42076 = _42074 ^ _42075;
  wire _42077 = _38970 ^ _2974;
  wire _42078 = _1425 ^ _5209;
  wire _42079 = _42077 ^ _42078;
  wire _42080 = _42076 ^ _42079;
  wire _42081 = _42073 ^ _42080;
  wire _42082 = _42067 ^ _42081;
  wire _42083 = _3762 ^ _1432;
  wire _42084 = uncoded_block[1222] ^ uncoded_block[1229];
  wire _42085 = _10059 ^ _42084;
  wire _42086 = _42083 ^ _42085;
  wire _42087 = _10067 ^ _1448;
  wire _42088 = _24465 ^ _42087;
  wire _42089 = _42086 ^ _42088;
  wire _42090 = _5231 ^ _20801;
  wire _42091 = _38179 ^ _42090;
  wire _42092 = _14418 ^ _627;
  wire _42093 = _2245 ^ _1463;
  wire _42094 = _42092 ^ _42093;
  wire _42095 = _42091 ^ _42094;
  wire _42096 = _42089 ^ _42095;
  wire _42097 = uncoded_block[1279] ^ uncoded_block[1283];
  wire _42098 = _5908 ^ _42097;
  wire _42099 = _28317 ^ _8980;
  wire _42100 = _42098 ^ _42099;
  wire _42101 = _3017 ^ _18870;
  wire _42102 = _2254 ^ _648;
  wire _42103 = _42101 ^ _42102;
  wire _42104 = _42100 ^ _42103;
  wire _42105 = _7802 ^ _7804;
  wire _42106 = _21293 ^ _4543;
  wire _42107 = _42105 ^ _42106;
  wire _42108 = _7201 ^ _5256;
  wire _42109 = _42108 ^ _22218;
  wire _42110 = _42107 ^ _42109;
  wire _42111 = _42104 ^ _42110;
  wire _42112 = _42096 ^ _42111;
  wire _42113 = _42082 ^ _42112;
  wire _42114 = _1501 ^ _5269;
  wire _42115 = uncoded_block[1351] ^ uncoded_block[1356];
  wire _42116 = _42115 ^ _5940;
  wire _42117 = _42114 ^ _42116;
  wire _42118 = _3045 ^ _2283;
  wire _42119 = _3052 ^ _3054;
  wire _42120 = _42118 ^ _42119;
  wire _42121 = _42117 ^ _42120;
  wire _42122 = _26743 ^ _3834;
  wire _42123 = _10108 ^ _12867;
  wire _42124 = _42122 ^ _42123;
  wire _42125 = _18901 ^ _12315;
  wire _42126 = _42125 ^ _28691;
  wire _42127 = _42124 ^ _42126;
  wire _42128 = _42121 ^ _42127;
  wire _42129 = _10117 ^ _2306;
  wire _42130 = _16463 ^ _32948;
  wire _42131 = _42129 ^ _42130;
  wire _42132 = _9591 ^ _22242;
  wire _42133 = _42132 ^ _14980;
  wire _42134 = _42131 ^ _42133;
  wire _42135 = _22700 ^ _25868;
  wire _42136 = _7243 ^ _7247;
  wire _42137 = _3090 ^ _42136;
  wire _42138 = _42135 ^ _42137;
  wire _42139 = _42134 ^ _42138;
  wire _42140 = _42128 ^ _42139;
  wire _42141 = _13446 ^ _15994;
  wire _42142 = _16978 ^ _42141;
  wire _42143 = _7861 ^ _16981;
  wire _42144 = _41369 ^ _10712;
  wire _42145 = _42143 ^ _42144;
  wire _42146 = _42142 ^ _42145;
  wire _42147 = _15002 ^ _3115;
  wire _42148 = _17493 ^ _42147;
  wire _42149 = uncoded_block[1528] ^ uncoded_block[1539];
  wire _42150 = _3900 ^ _42149;
  wire _42151 = _34223 ^ _42150;
  wire _42152 = _42148 ^ _42151;
  wire _42153 = _42146 ^ _42152;
  wire _42154 = _3128 ^ _17998;
  wire _42155 = _767 ^ _28378;
  wire _42156 = _42154 ^ _42155;
  wire _42157 = _36240 ^ _27202;
  wire _42158 = _2379 ^ _782;
  wire _42159 = _42157 ^ _42158;
  wire _42160 = _42156 ^ _42159;
  wire _42161 = _20397 ^ _5368;
  wire _42162 = uncoded_block[1591] ^ uncoded_block[1597];
  wire _42163 = _42162 ^ _11295;
  wire _42164 = _42161 ^ _42163;
  wire _42165 = _3151 ^ _3153;
  wire _42166 = uncoded_block[1607] ^ uncoded_block[1611];
  wire _42167 = _42166 ^ _7908;
  wire _42168 = _42165 ^ _42167;
  wire _42169 = _42164 ^ _42168;
  wire _42170 = _42160 ^ _42169;
  wire _42171 = _42153 ^ _42170;
  wire _42172 = _42140 ^ _42171;
  wire _42173 = _42113 ^ _42172;
  wire _42174 = _7298 ^ _13494;
  wire _42175 = _12947 ^ _1639;
  wire _42176 = _42174 ^ _42175;
  wire _42177 = uncoded_block[1632] ^ uncoded_block[1637];
  wire _42178 = _42177 ^ _7308;
  wire _42179 = _13500 ^ _5394;
  wire _42180 = _42178 ^ _42179;
  wire _42181 = _42176 ^ _42180;
  wire _42182 = _6691 ^ _3172;
  wire _42183 = _42182 ^ _37888;
  wire _42184 = _41411 ^ _7320;
  wire _42185 = _42183 ^ _42184;
  wire _42186 = _42181 ^ _42185;
  wire _42187 = uncoded_block[1670] ^ uncoded_block[1674];
  wire _42188 = _42187 ^ _33862;
  wire _42189 = _20427 ^ _3965;
  wire _42190 = _42188 ^ _42189;
  wire _42191 = uncoded_block[1689] ^ uncoded_block[1694];
  wire _42192 = _42191 ^ _11327;
  wire _42193 = _845 ^ _3976;
  wire _42194 = _42192 ^ _42193;
  wire _42195 = _42190 ^ _42194;
  wire _42196 = _30908 ^ _2443;
  wire _42197 = _3981 ^ _42196;
  wire _42198 = _42197 ^ _12977;
  wire _42199 = _42195 ^ _42198;
  wire _42200 = _42186 ^ _42199;
  wire _42201 = _42173 ^ _42200;
  wire _42202 = _42052 ^ _42201;
  wire _42203 = _2 ^ _19960;
  wire _42204 = uncoded_block[10] ^ uncoded_block[14];
  wire _42205 = _42204 ^ _9692;
  wire _42206 = _3217 ^ _13539;
  wire _42207 = _42205 ^ _42206;
  wire _42208 = _42203 ^ _42207;
  wire _42209 = _875 ^ _18548;
  wire _42210 = _42209 ^ _12991;
  wire _42211 = _6099 ^ _25;
  wire _42212 = _15084 ^ _42211;
  wire _42213 = _42210 ^ _42212;
  wire _42214 = _42208 ^ _42213;
  wire _42215 = uncoded_block[66] ^ uncoded_block[73];
  wire _42216 = _31 ^ _42215;
  wire _42217 = _39 ^ _2481;
  wire _42218 = _42216 ^ _42217;
  wire _42219 = _28438 ^ _9713;
  wire _42220 = uncoded_block[90] ^ uncoded_block[100];
  wire _42221 = _42220 ^ _2490;
  wire _42222 = _42219 ^ _42221;
  wire _42223 = _42218 ^ _42222;
  wire _42224 = _37135 ^ _2498;
  wire _42225 = _18562 ^ _42224;
  wire _42226 = _7386 ^ _32634;
  wire _42227 = _42226 ^ _14078;
  wire _42228 = _42225 ^ _42227;
  wire _42229 = _42223 ^ _42228;
  wire _42230 = _42214 ^ _42229;
  wire _42231 = uncoded_block[141] ^ uncoded_block[144];
  wire _42232 = _42231 ^ _14082;
  wire _42233 = _8003 ^ _14085;
  wire _42234 = _42232 ^ _42233;
  wire _42235 = _11392 ^ _2524;
  wire _42236 = _33073 ^ _42235;
  wire _42237 = _42234 ^ _42236;
  wire _42238 = _8009 ^ _13583;
  wire _42239 = _42238 ^ _22369;
  wire _42240 = uncoded_block[193] ^ uncoded_block[201];
  wire _42241 = _42240 ^ _3289;
  wire _42242 = _33082 ^ _17116;
  wire _42243 = _42241 ^ _42242;
  wire _42244 = _42239 ^ _42243;
  wire _42245 = _42237 ^ _42244;
  wire _42246 = _35912 ^ _6814;
  wire _42247 = _1774 ^ _8029;
  wire _42248 = _42246 ^ _42247;
  wire _42249 = _6824 ^ _6179;
  wire _42250 = _4087 ^ _11419;
  wire _42251 = _42249 ^ _42250;
  wire _42252 = _42248 ^ _42251;
  wire _42253 = _20023 ^ _20520;
  wire _42254 = _977 ^ _1792;
  wire _42255 = _42253 ^ _42254;
  wire _42256 = _3320 ^ _19570;
  wire _42257 = _7445 ^ _10304;
  wire _42258 = _42256 ^ _42257;
  wire _42259 = _42255 ^ _42258;
  wire _42260 = _42252 ^ _42259;
  wire _42261 = _42245 ^ _42260;
  wire _42262 = _42230 ^ _42261;
  wire _42263 = _13066 ^ _22861;
  wire _42264 = _4820 ^ _138;
  wire _42265 = _35933 ^ _8055;
  wire _42266 = _42264 ^ _42265;
  wire _42267 = _42263 ^ _42266;
  wire _42268 = _5528 ^ _39170;
  wire _42269 = _3341 ^ _1008;
  wire _42270 = _42268 ^ _42269;
  wire _42271 = _18147 ^ _2586;
  wire _42272 = _3348 ^ _42271;
  wire _42273 = _42270 ^ _42272;
  wire _42274 = _42267 ^ _42273;
  wire _42275 = _22873 ^ _26026;
  wire _42276 = _42275 ^ _37979;
  wire _42277 = uncoded_block[351] ^ uncoded_block[355];
  wire _42278 = _161 ^ _42277;
  wire _42279 = _21030 ^ _168;
  wire _42280 = _42278 ^ _42279;
  wire _42281 = _42276 ^ _42280;
  wire _42282 = uncoded_block[367] ^ uncoded_block[373];
  wire _42283 = _42282 ^ _4141;
  wire _42284 = _12538 ^ _1045;
  wire _42285 = _42283 ^ _42284;
  wire _42286 = uncoded_block[392] ^ uncoded_block[395];
  wire _42287 = _42286 ^ _1849;
  wire _42288 = uncoded_block[402] ^ uncoded_block[407];
  wire _42289 = _181 ^ _42288;
  wire _42290 = _42287 ^ _42289;
  wire _42291 = _42285 ^ _42290;
  wire _42292 = _42281 ^ _42291;
  wire _42293 = _42274 ^ _42292;
  wire _42294 = _35182 ^ _22897;
  wire _42295 = uncoded_block[423] ^ uncoded_block[427];
  wire _42296 = _42295 ^ _2638;
  wire _42297 = _6255 ^ _5574;
  wire _42298 = _42296 ^ _42297;
  wire _42299 = _42294 ^ _42298;
  wire _42300 = uncoded_block[440] ^ uncoded_block[446];
  wire _42301 = _42300 ^ _11486;
  wire _42302 = _42301 ^ _26058;
  wire _42303 = _5584 ^ _8681;
  wire _42304 = uncoded_block[469] ^ uncoded_block[474];
  wire _42305 = uncoded_block[475] ^ uncoded_block[480];
  wire _42306 = _42304 ^ _42305;
  wire _42307 = _42303 ^ _42306;
  wire _42308 = _42302 ^ _42307;
  wire _42309 = _42299 ^ _42308;
  wire _42310 = _18658 ^ _14701;
  wire _42311 = uncoded_block[499] ^ uncoded_block[505];
  wire _42312 = _42311 ^ _5611;
  wire _42313 = _3433 ^ _42312;
  wire _42314 = _42310 ^ _42313;
  wire _42315 = _20598 ^ _3444;
  wire _42316 = _8123 ^ _42315;
  wire _42317 = uncoded_block[523] ^ uncoded_block[532];
  wire _42318 = _42317 ^ _1905;
  wire _42319 = _42318 ^ _37239;
  wire _42320 = _42316 ^ _42319;
  wire _42321 = _42314 ^ _42320;
  wire _42322 = _42309 ^ _42321;
  wire _42323 = _42293 ^ _42322;
  wire _42324 = _42262 ^ _42323;
  wire _42325 = _1910 ^ _31487;
  wire _42326 = _8725 ^ _1126;
  wire _42327 = _7550 ^ _3468;
  wire _42328 = _42326 ^ _42327;
  wire _42329 = _42325 ^ _42328;
  wire _42330 = _17221 ^ _262;
  wire _42331 = _19652 ^ _15247;
  wire _42332 = _42330 ^ _42331;
  wire _42333 = _3486 ^ _8152;
  wire _42334 = _20626 ^ _6325;
  wire _42335 = _42333 ^ _42334;
  wire _42336 = _42332 ^ _42335;
  wire _42337 = _42329 ^ _42336;
  wire _42338 = _1149 ^ _3494;
  wire _42339 = _3495 ^ _10418;
  wire _42340 = _42338 ^ _42339;
  wire _42341 = uncoded_block[626] ^ uncoded_block[631];
  wire _42342 = _42341 ^ _3501;
  wire _42343 = _42342 ^ _17241;
  wire _42344 = _42340 ^ _42343;
  wire _42345 = _9878 ^ _13724;
  wire _42346 = _20638 ^ _15273;
  wire _42347 = _40796 ^ _42346;
  wire _42348 = _42345 ^ _42347;
  wire _42349 = _42344 ^ _42348;
  wire _42350 = _42337 ^ _42349;
  wire _42351 = _17742 ^ _312;
  wire _42352 = uncoded_block[673] ^ uncoded_block[681];
  wire _42353 = _42352 ^ _3526;
  wire _42354 = _42351 ^ _42353;
  wire _42355 = _322 ^ _32767;
  wire _42356 = _42355 ^ _12094;
  wire _42357 = _42354 ^ _42356;
  wire _42358 = _17266 ^ _18259;
  wire _42359 = _31083 ^ _42358;
  wire _42360 = _11006 ^ _8201;
  wire _42361 = _23870 ^ _5010;
  wire _42362 = _42360 ^ _42361;
  wire _42363 = _42359 ^ _42362;
  wire _42364 = _42357 ^ _42363;
  wire _42365 = _11576 ^ _5012;
  wire _42366 = _1210 ^ _23879;
  wire _42367 = _42365 ^ _42366;
  wire _42368 = _17776 ^ _7019;
  wire _42369 = _4302 ^ _42368;
  wire _42370 = _42367 ^ _42369;
  wire _42371 = _7022 ^ _18747;
  wire _42372 = _5032 ^ _28559;
  wire _42373 = _385 ^ _3577;
  wire _42374 = _42372 ^ _42373;
  wire _42375 = _42371 ^ _42374;
  wire _42376 = _42370 ^ _42375;
  wire _42377 = _42364 ^ _42376;
  wire _42378 = _42350 ^ _42377;
  wire _42379 = _5727 ^ _392;
  wire _42380 = _393 ^ _1242;
  wire _42381 = _42379 ^ _42380;
  wire _42382 = _42381 ^ _40465;
  wire _42383 = uncoded_block[843] ^ uncoded_block[850];
  wire _42384 = _5737 ^ _42383;
  wire _42385 = _42384 ^ _30257;
  wire _42386 = _15825 ^ _41625;
  wire _42387 = _42385 ^ _42386;
  wire _42388 = _42382 ^ _42387;
  wire _42389 = _16815 ^ _2836;
  wire _42390 = _423 ^ _4354;
  wire _42391 = _42389 ^ _42390;
  wire _42392 = _21636 ^ _428;
  wire _42393 = uncoded_block[899] ^ uncoded_block[904];
  wire _42394 = _42393 ^ _3623;
  wire _42395 = _42392 ^ _42394;
  wire _42396 = _42391 ^ _42395;
  wire _42397 = uncoded_block[913] ^ uncoded_block[918];
  wire _42398 = _16312 ^ _42397;
  wire _42399 = uncoded_block[920] ^ uncoded_block[924];
  wire _42400 = uncoded_block[927] ^ uncoded_block[937];
  wire _42401 = _42399 ^ _42400;
  wire _42402 = _42398 ^ _42401;
  wire _42403 = uncoded_block[951] ^ uncoded_block[958];
  wire _42404 = _5777 ^ _42403;
  wire _42405 = _3642 ^ _42404;
  wire _42406 = _42402 ^ _42405;
  wire _42407 = _42396 ^ _42406;
  wire _42408 = _42388 ^ _42407;
  wire _42409 = _4385 ^ _10531;
  wire _42410 = _42409 ^ _7089;
  wire _42411 = _468 ^ _32425;
  wire _42412 = _7689 ^ _16338;
  wire _42413 = _42411 ^ _42412;
  wire _42414 = _42410 ^ _42413;
  wire _42415 = _13277 ^ _38517;
  wire _42416 = _22122 ^ _6459;
  wire _42417 = _42415 ^ _42416;
  wire _42418 = _491 ^ _11663;
  wire _42419 = _42418 ^ _20737;
  wire _42420 = _42417 ^ _42419;
  wire _42421 = _42414 ^ _42420;
  wire _42422 = _12199 ^ _11114;
  wire _42423 = _2909 ^ _42422;
  wire _42424 = _19295 ^ _12762;
  wire _42425 = _7117 ^ _4433;
  wire _42426 = _42424 ^ _42425;
  wire _42427 = _42423 ^ _42426;
  wire _42428 = _3685 ^ _10569;
  wire _42429 = _25773 ^ _5158;
  wire _42430 = _42428 ^ _42429;
  wire _42431 = _20251 ^ _20753;
  wire _42432 = _42431 ^ _13858;
  wire _42433 = _42430 ^ _42432;
  wire _42434 = _42427 ^ _42433;
  wire _42435 = _42421 ^ _42434;
  wire _42436 = _42408 ^ _42435;
  wire _42437 = _42378 ^ _42436;
  wire _42438 = _42324 ^ _42437;
  wire _42439 = _3698 ^ _11139;
  wire _42440 = uncoded_block[1102] ^ uncoded_block[1107];
  wire _42441 = _42440 ^ _13319;
  wire _42442 = _42439 ^ _42441;
  wire _42443 = _5175 ^ _7736;
  wire _42444 = _12789 ^ _6499;
  wire _42445 = _42443 ^ _42444;
  wire _42446 = _42442 ^ _42445;
  wire _42447 = _9494 ^ _5856;
  wire _42448 = _42447 ^ _32052;
  wire _42449 = _2956 ^ _17386;
  wire _42450 = _12239 ^ _42449;
  wire _42451 = _42448 ^ _42450;
  wire _42452 = _42446 ^ _42451;
  wire _42453 = uncoded_block[1162] ^ uncoded_block[1174];
  wire _42454 = _12243 ^ _42453;
  wire _42455 = _16898 ^ _592;
  wire _42456 = _42454 ^ _42455;
  wire _42457 = _13886 ^ _2207;
  wire _42458 = _5204 ^ _42457;
  wire _42459 = _42456 ^ _42458;
  wire _42460 = _27911 ^ _10620;
  wire _42461 = _2980 ^ _42460;
  wire _42462 = _12815 ^ _5891;
  wire _42463 = _1436 ^ _1439;
  wire _42464 = _42462 ^ _42463;
  wire _42465 = _42461 ^ _42464;
  wire _42466 = _42459 ^ _42465;
  wire _42467 = _42452 ^ _42466;
  wire _42468 = _15927 ^ _10067;
  wire _42469 = _4509 ^ _33758;
  wire _42470 = _42468 ^ _42469;
  wire _42471 = _6546 ^ _3783;
  wire _42472 = _42471 ^ _17421;
  wire _42473 = _42470 ^ _42472;
  wire _42474 = _24930 ^ _26720;
  wire _42475 = _28317 ^ _24482;
  wire _42476 = _42475 ^ _25378;
  wire _42477 = _42474 ^ _42476;
  wire _42478 = _42473 ^ _42477;
  wire _42479 = _20812 ^ _3807;
  wire _42480 = _39385 ^ _42479;
  wire _42481 = _17435 ^ _2262;
  wire _42482 = _4540 ^ _5254;
  wire _42483 = _42481 ^ _42482;
  wire _42484 = _42480 ^ _42483;
  wire _42485 = _3820 ^ _39393;
  wire _42486 = _10656 ^ _42485;
  wire _42487 = _11218 ^ _5938;
  wire _42488 = _41338 ^ _42487;
  wire _42489 = _42486 ^ _42488;
  wire _42490 = _42484 ^ _42489;
  wire _42491 = _42478 ^ _42490;
  wire _42492 = _42467 ^ _42491;
  wire _42493 = _12857 ^ _23581;
  wire _42494 = _23148 ^ _10101;
  wire _42495 = _42493 ^ _42494;
  wire _42496 = _40945 ^ _5284;
  wire _42497 = _25399 ^ _691;
  wire _42498 = _42496 ^ _42497;
  wire _42499 = _42495 ^ _42498;
  wire _42500 = _13412 ^ _7834;
  wire _42501 = uncoded_block[1399] ^ uncoded_block[1403];
  wire _42502 = _42501 ^ _701;
  wire _42503 = _42500 ^ _42502;
  wire _42504 = uncoded_block[1411] ^ uncoded_block[1414];
  wire _42505 = _8436 ^ _42504;
  wire _42506 = _10118 ^ _10683;
  wire _42507 = _42505 ^ _42506;
  wire _42508 = _42503 ^ _42507;
  wire _42509 = _42499 ^ _42508;
  wire _42510 = _1531 ^ _9595;
  wire _42511 = _12879 ^ _42510;
  wire _42512 = uncoded_block[1450] ^ uncoded_block[1452];
  wire _42513 = _2325 ^ _42512;
  wire _42514 = _5306 ^ _42513;
  wire _42515 = _42511 ^ _42514;
  wire _42516 = _2328 ^ _5309;
  wire _42517 = _3089 ^ _20361;
  wire _42518 = _42516 ^ _42517;
  wire _42519 = _3094 ^ _1550;
  wire _42520 = _18919 ^ _11255;
  wire _42521 = _42519 ^ _42520;
  wire _42522 = _42518 ^ _42521;
  wire _42523 = _42515 ^ _42522;
  wire _42524 = _42509 ^ _42523;
  wire _42525 = _733 ^ _34615;
  wire _42526 = _9042 ^ _1562;
  wire _42527 = _42525 ^ _42526;
  wire _42528 = _17489 ^ _2350;
  wire _42529 = _12899 ^ _1572;
  wire _42530 = _42528 ^ _42529;
  wire _42531 = _42527 ^ _42530;
  wire _42532 = _5334 ^ _19429;
  wire _42533 = _28370 ^ _42532;
  wire _42534 = _5337 ^ _12352;
  wire _42535 = _9059 ^ _4623;
  wire _42536 = _42534 ^ _42535;
  wire _42537 = _42533 ^ _42536;
  wire _42538 = _42531 ^ _42537;
  wire _42539 = _13461 ^ _24091;
  wire _42540 = _6008 ^ _4634;
  wire _42541 = _42540 ^ _8483;
  wire _42542 = _42539 ^ _42541;
  wire _42543 = _3914 ^ _6019;
  wire _42544 = _16997 ^ _42543;
  wire _42545 = _18949 ^ _782;
  wire _42546 = _42545 ^ _15030;
  wire _42547 = _42544 ^ _42546;
  wire _42548 = _42542 ^ _42547;
  wire _42549 = _42538 ^ _42548;
  wire _42550 = _42524 ^ _42549;
  wire _42551 = _42492 ^ _42550;
  wire _42552 = _2386 ^ _15538;
  wire _42553 = _42552 ^ _29994;
  wire _42554 = _1627 ^ _4662;
  wire _42555 = _28398 ^ _42554;
  wire _42556 = _42553 ^ _42555;
  wire _42557 = _16032 ^ _18511;
  wire _42558 = _19929 ^ _3169;
  wire _42559 = _42557 ^ _42558;
  wire _42560 = _819 ^ _4678;
  wire _42561 = _7925 ^ _20909;
  wire _42562 = _42560 ^ _42561;
  wire _42563 = _42559 ^ _42562;
  wire _42564 = _42556 ^ _42563;
  wire _42565 = _17032 ^ _6700;
  wire _42566 = _42565 ^ _41415;
  wire _42567 = _6705 ^ _7935;
  wire _42568 = _28417 ^ _42567;
  wire _42569 = _42566 ^ _42568;
  wire _42570 = _26830 ^ _20919;
  wire _42571 = _2438 ^ _3200;
  wire _42572 = _23235 ^ _42571;
  wire _42573 = _42570 ^ _42572;
  wire _42574 = _42569 ^ _42573;
  wire _42575 = _42564 ^ _42574;
  wire _42576 = _42575 ^ _37104;
  wire _42577 = _42551 ^ _42576;
  wire _42578 = _42438 ^ _42577;
  wire _42579 = uncoded_block[16] ^ uncoded_block[21];
  wire _42580 = _15075 ^ _42579;
  wire _42581 = _16562 ^ _42580;
  wire _42582 = uncoded_block[24] ^ uncoded_block[29];
  wire _42583 = _42582 ^ _18548;
  wire _42584 = uncoded_block[37] ^ uncoded_block[46];
  wire _42585 = _42584 ^ _8556;
  wire _42586 = _42583 ^ _42585;
  wire _42587 = _42581 ^ _42586;
  wire _42588 = _10806 ^ _1712;
  wire _42589 = _1714 ^ _19019;
  wire _42590 = _42588 ^ _42589;
  wire _42591 = uncoded_block[85] ^ uncoded_block[87];
  wire _42592 = _11364 ^ _42591;
  wire _42593 = _903 ^ _4741;
  wire _42594 = _42592 ^ _42593;
  wire _42595 = _42590 ^ _42594;
  wire _42596 = _42587 ^ _42595;
  wire _42597 = uncoded_block[98] ^ uncoded_block[104];
  wire _42598 = _42597 ^ _15103;
  wire _42599 = _10816 ^ _54;
  wire _42600 = _42598 ^ _42599;
  wire _42601 = _10256 ^ _38723;
  wire _42602 = uncoded_block[148] ^ uncoded_block[155];
  wire _42603 = _4046 ^ _42602;
  wire _42604 = _42601 ^ _42603;
  wire _42605 = _42600 ^ _42604;
  wire _42606 = _29208 ^ _29210;
  wire _42607 = uncoded_block[180] ^ uncoded_block[189];
  wire _42608 = _82 ^ _42607;
  wire _42609 = _42606 ^ _42608;
  wire _42610 = _7411 ^ _4070;
  wire _42611 = _42610 ^ _7416;
  wire _42612 = _42609 ^ _42611;
  wire _42613 = _42605 ^ _42612;
  wire _42614 = _42596 ^ _42613;
  wire _42615 = _24655 ^ _3299;
  wire _42616 = uncoded_block[237] ^ uncoded_block[246];
  wire _42617 = _24660 ^ _42616;
  wire _42618 = _42615 ^ _42617;
  wire _42619 = uncoded_block[252] ^ uncoded_block[265];
  wire _42620 = _8617 ^ _42619;
  wire _42621 = uncoded_block[270] ^ uncoded_block[278];
  wire _42622 = uncoded_block[282] ^ uncoded_block[292];
  wire _42623 = _42621 ^ _42622;
  wire _42624 = _42620 ^ _42623;
  wire _42625 = _42618 ^ _42624;
  wire _42626 = uncoded_block[315] ^ uncoded_block[322];
  wire _42627 = _26905 ^ _42626;
  wire _42628 = _26013 ^ _42627;
  wire _42629 = _8642 ^ _1819;
  wire _42630 = _2593 ^ _1826;
  wire _42631 = _42629 ^ _42630;
  wire _42632 = _42628 ^ _42631;
  wire _42633 = _42625 ^ _42632;
  wire _42634 = _4132 ^ _13089;
  wire _42635 = _3369 ^ _11999;
  wire _42636 = _42634 ^ _42635;
  wire _42637 = _10907 ^ _2616;
  wire _42638 = uncoded_block[397] ^ uncoded_block[403];
  wire _42639 = _42638 ^ _5564;
  wire _42640 = _42637 ^ _42639;
  wire _42641 = _42636 ^ _42640;
  wire _42642 = _40748 ^ _2637;
  wire _42643 = _201 ^ _21516;
  wire _42644 = _42642 ^ _42643;
  wire _42645 = _9275 ^ _33565;
  wire _42646 = uncoded_block[462] ^ uncoded_block[466];
  wire _42647 = _3415 ^ _42646;
  wire _42648 = _42645 ^ _42647;
  wire _42649 = _42644 ^ _42648;
  wire _42650 = _42641 ^ _42649;
  wire _42651 = _42633 ^ _42650;
  wire _42652 = _42614 ^ _42651;
  wire _42653 = uncoded_block[470] ^ uncoded_block[478];
  wire _42654 = uncoded_block[481] ^ uncoded_block[488];
  wire _42655 = _42653 ^ _42654;
  wire _42656 = _42655 ^ _13140;
  wire _42657 = _8120 ^ _6285;
  wire _42658 = _28503 ^ _33587;
  wire _42659 = _42657 ^ _42658;
  wire _42660 = _42656 ^ _42659;
  wire _42661 = uncoded_block[543] ^ uncoded_block[550];
  wire _42662 = _243 ^ _42661;
  wire _42663 = _42662 ^ _8138;
  wire _42664 = _1927 ^ _3472;
  wire _42665 = _42664 ^ _1932;
  wire _42666 = _42663 ^ _42665;
  wire _42667 = _42660 ^ _42666;
  wire _42668 = _20116 ^ _4234;
  wire _42669 = uncoded_block[600] ^ uncoded_block[605];
  wire _42670 = _6316 ^ _42669;
  wire _42671 = _42668 ^ _42670;
  wire _42672 = _4963 ^ _15261;
  wire _42673 = uncoded_block[628] ^ uncoded_block[636];
  wire _42674 = uncoded_block[639] ^ uncoded_block[648];
  wire _42675 = _42673 ^ _42674;
  wire _42676 = _42672 ^ _42675;
  wire _42677 = _42671 ^ _42676;
  wire _42678 = _12080 ^ _5671;
  wire _42679 = _303 ^ _42678;
  wire _42680 = _1180 ^ _4984;
  wire _42681 = _313 ^ _42680;
  wire _42682 = _42679 ^ _42681;
  wire _42683 = _42677 ^ _42682;
  wire _42684 = _42667 ^ _42683;
  wire _42685 = _2757 ^ _23863;
  wire _42686 = _1192 ^ _8193;
  wire _42687 = _42685 ^ _42686;
  wire _42688 = _9369 ^ _7603;
  wire _42689 = _1995 ^ _15300;
  wire _42690 = _42688 ^ _42689;
  wire _42691 = _42687 ^ _42690;
  wire _42692 = _8209 ^ _2003;
  wire _42693 = uncoded_block[756] ^ uncoded_block[771];
  wire _42694 = _42693 ^ _13219;
  wire _42695 = _42692 ^ _42694;
  wire _42696 = _25694 ^ _12675;
  wire _42697 = _374 ^ _383;
  wire _42698 = _42696 ^ _42697;
  wire _42699 = _42695 ^ _42698;
  wire _42700 = _42691 ^ _42699;
  wire _42701 = _4317 ^ _36477;
  wire _42702 = _42701 ^ _22526;
  wire _42703 = uncoded_block[836] ^ uncoded_block[842];
  wire _42704 = _1246 ^ _42703;
  wire _42705 = _42704 ^ _5061;
  wire _42706 = _42702 ^ _42705;
  wire _42707 = uncoded_block[863] ^ uncoded_block[873];
  wire _42708 = _19236 ^ _42707;
  wire _42709 = _9954 ^ _2836;
  wire _42710 = _42708 ^ _42709;
  wire _42711 = _11059 ^ _18307;
  wire _42712 = _8250 ^ _6424;
  wire _42713 = _42711 ^ _42712;
  wire _42714 = _42710 ^ _42713;
  wire _42715 = _42706 ^ _42714;
  wire _42716 = _42700 ^ _42715;
  wire _42717 = _42684 ^ _42716;
  wire _42718 = _42652 ^ _42717;
  wire _42719 = uncoded_block[914] ^ uncoded_block[922];
  wire _42720 = _42719 ^ _6435;
  wire _42721 = _7071 ^ _42720;
  wire _42722 = _13266 ^ _1308;
  wire _42723 = _8263 ^ _42722;
  wire _42724 = _42721 ^ _42723;
  wire _42725 = _36515 ^ _28233;
  wire _42726 = _42725 ^ _40859;
  wire _42727 = _19277 ^ _2114;
  wire _42728 = uncoded_block[1009] ^ uncoded_block[1016];
  wire _42729 = _42728 ^ _2893;
  wire _42730 = _42727 ^ _42729;
  wire _42731 = _42726 ^ _42730;
  wire _42732 = _42724 ^ _42731;
  wire _42733 = _498 ^ _3676;
  wire _42734 = _19777 ^ _40871;
  wire _42735 = _42733 ^ _42734;
  wire _42736 = uncoded_block[1076] ^ uncoded_block[1081];
  wire _42737 = _13851 ^ _42736;
  wire _42738 = _14356 ^ _42737;
  wire _42739 = _42735 ^ _42738;
  wire _42740 = _533 ^ _537;
  wire _42741 = uncoded_block[1099] ^ uncoded_block[1104];
  wire _42742 = _42741 ^ _3708;
  wire _42743 = _42740 ^ _42742;
  wire _42744 = uncoded_block[1112] ^ uncoded_block[1118];
  wire _42745 = _1385 ^ _42744;
  wire _42746 = uncoded_block[1123] ^ uncoded_block[1132];
  wire _42747 = _42746 ^ _10591;
  wire _42748 = _42745 ^ _42747;
  wire _42749 = _42743 ^ _42748;
  wire _42750 = _42739 ^ _42749;
  wire _42751 = _42732 ^ _42750;
  wire _42752 = _8929 ^ _574;
  wire _42753 = _4465 ^ _3728;
  wire _42754 = _42752 ^ _42753;
  wire _42755 = _2188 ^ _2964;
  wire _42756 = _42755 ^ _18844;
  wire _42757 = _42754 ^ _42756;
  wire _42758 = _3739 ^ _5200;
  wire _42759 = _23996 ^ _6522;
  wire _42760 = _42758 ^ _42759;
  wire _42761 = _40903 ^ _24456;
  wire _42762 = uncoded_block[1223] ^ uncoded_block[1229];
  wire _42763 = _42762 ^ _19827;
  wire _42764 = _42761 ^ _42763;
  wire _42765 = _42760 ^ _42764;
  wire _42766 = _42757 ^ _42765;
  wire _42767 = uncoded_block[1240] ^ uncoded_block[1248];
  wire _42768 = _42767 ^ _5902;
  wire _42769 = _7781 ^ _30361;
  wire _42770 = _42768 ^ _42769;
  wire _42771 = _26718 ^ _15455;
  wire _42772 = _1469 ^ _9547;
  wire _42773 = _42771 ^ _42772;
  wire _42774 = _42770 ^ _42773;
  wire _42775 = _7799 ^ _28665;
  wire _42776 = uncoded_block[1310] ^ uncoded_block[1315];
  wire _42777 = _42776 ^ _24942;
  wire _42778 = _42775 ^ _42777;
  wire _42779 = uncoded_block[1321] ^ uncoded_block[1327];
  wire _42780 = _42779 ^ _4550;
  wire _42781 = _9563 ^ _2277;
  wire _42782 = _42780 ^ _42781;
  wire _42783 = _42778 ^ _42782;
  wire _42784 = _42774 ^ _42783;
  wire _42785 = _42766 ^ _42784;
  wire _42786 = _42751 ^ _42785;
  wire _42787 = uncoded_block[1348] ^ uncoded_block[1354];
  wire _42788 = uncoded_block[1356] ^ uncoded_block[1364];
  wire _42789 = _42787 ^ _42788;
  wire _42790 = _10668 ^ _7823;
  wire _42791 = _42789 ^ _42790;
  wire _42792 = uncoded_block[1383] ^ uncoded_block[1395];
  wire _42793 = _4564 ^ _42792;
  wire _42794 = _30821 ^ _42504;
  wire _42795 = _42793 ^ _42794;
  wire _42796 = _42791 ^ _42795;
  wire _42797 = uncoded_block[1415] ^ uncoded_block[1425];
  wire _42798 = _42797 ^ _3075;
  wire _42799 = uncoded_block[1431] ^ uncoded_block[1436];
  wire _42800 = _42799 ^ _24521;
  wire _42801 = _42798 ^ _42800;
  wire _42802 = uncoded_block[1452] ^ uncoded_block[1464];
  wire _42803 = _42802 ^ _2338;
  wire _42804 = _40962 ^ _42803;
  wire _42805 = _42801 ^ _42804;
  wire _42806 = _42796 ^ _42805;
  wire _42807 = uncoded_block[1473] ^ uncoded_block[1477];
  wire _42808 = _42807 ^ _1556;
  wire _42809 = uncoded_block[1485] ^ uncoded_block[1494];
  wire _42810 = _9042 ^ _42809;
  wire _42811 = _42808 ^ _42810;
  wire _42812 = _30419 ^ _15515;
  wire _42813 = _16488 ^ _7265;
  wire _42814 = _42812 ^ _42813;
  wire _42815 = _42811 ^ _42814;
  wire _42816 = uncoded_block[1538] ^ uncoded_block[1559];
  wire _42817 = _36656 ^ _42816;
  wire _42818 = _5342 ^ _42817;
  wire _42819 = uncoded_block[1566] ^ uncoded_block[1572];
  wire _42820 = _3139 ^ _42819;
  wire _42821 = _40989 ^ _3927;
  wire _42822 = _42820 ^ _42821;
  wire _42823 = _42818 ^ _42822;
  wire _42824 = _42815 ^ _42823;
  wire _42825 = _42806 ^ _42824;
  wire _42826 = _4653 ^ _39062;
  wire _42827 = _11295 ^ _9088;
  wire _42828 = _42826 ^ _42827;
  wire _42829 = uncoded_block[1617] ^ uncoded_block[1626];
  wire _42830 = _42829 ^ _14525;
  wire _42831 = uncoded_block[1632] ^ uncoded_block[1639];
  wire _42832 = _42831 ^ _2411;
  wire _42833 = _42830 ^ _42832;
  wire _42834 = _42828 ^ _42833;
  wire _42835 = _12387 ^ _3958;
  wire _42836 = uncoded_block[1668] ^ uncoded_block[1674];
  wire _42837 = _5399 ^ _42836;
  wire _42838 = _42835 ^ _42837;
  wire _42839 = _41010 ^ _14543;
  wire _42840 = _9677 ^ _9120;
  wire _42841 = _42839 ^ _42840;
  wire _42842 = _42838 ^ _42841;
  wire _42843 = _42834 ^ _42842;
  wire _42844 = _3976 ^ _30908;
  wire _42845 = _42844 ^ uncoded_block[1721];
  wire _42846 = _42843 ^ _42845;
  wire _42847 = _42825 ^ _42846;
  wire _42848 = _42786 ^ _42847;
  wire _42849 = _42718 ^ _42848;
  wire _42850 = _21861 ^ _6082;
  wire _42851 = _42850 ^ _27996;
  wire _42852 = _4716 ^ _4000;
  wire _42853 = _5427 ^ _11;
  wire _42854 = _42852 ^ _42853;
  wire _42855 = _42851 ^ _42854;
  wire _42856 = _14045 ^ _2467;
  wire _42857 = _32211 ^ _1699;
  wire _42858 = uncoded_block[52] ^ uncoded_block[56];
  wire _42859 = _42858 ^ _13552;
  wire _42860 = _42857 ^ _42859;
  wire _42861 = _42856 ^ _42860;
  wire _42862 = _42855 ^ _42861;
  wire _42863 = _27254 ^ _26854;
  wire _42864 = _14061 ^ _36725;
  wire _42865 = _42863 ^ _42864;
  wire _42866 = _30933 ^ _40302;
  wire _42867 = _15101 ^ _6122;
  wire _42868 = _35506 ^ _42867;
  wire _42869 = _42866 ^ _42868;
  wire _42870 = _42865 ^ _42869;
  wire _42871 = _42862 ^ _42870;
  wire _42872 = _6763 ^ _54;
  wire _42873 = _42872 ^ _23714;
  wire _42874 = _3255 ^ _41846;
  wire _42875 = uncoded_block[131] ^ uncoded_block[135];
  wire _42876 = _923 ^ _42875;
  wire _42877 = _42874 ^ _42876;
  wire _42878 = _42873 ^ _42877;
  wire _42879 = _4760 ^ _6776;
  wire _42880 = _16600 ^ _1742;
  wire _42881 = _42879 ^ _42880;
  wire _42882 = uncoded_block[147] ^ uncoded_block[150];
  wire _42883 = _42882 ^ _3269;
  wire _42884 = _1748 ^ _933;
  wire _42885 = _42883 ^ _42884;
  wire _42886 = _42881 ^ _42885;
  wire _42887 = _42878 ^ _42886;
  wire _42888 = uncoded_block[169] ^ uncoded_block[173];
  wire _42889 = _16604 ^ _42888;
  wire _42890 = _3278 ^ _9195;
  wire _42891 = _42889 ^ _42890;
  wire _42892 = _13583 ^ _17106;
  wire _42893 = _2529 ^ _4776;
  wire _42894 = _42892 ^ _42893;
  wire _42895 = _42891 ^ _42894;
  wire _42896 = _25983 ^ _33082;
  wire _42897 = _34316 ^ _42896;
  wire _42898 = _37951 ^ _38336;
  wire _42899 = _42897 ^ _42898;
  wire _42900 = _42895 ^ _42899;
  wire _42901 = _42887 ^ _42900;
  wire _42902 = _42871 ^ _42901;
  wire _42903 = _4080 ^ _1775;
  wire _42904 = _42903 ^ _28051;
  wire _42905 = uncoded_block[246] ^ uncoded_block[254];
  wire _42906 = _42905 ^ _119;
  wire _42907 = _4798 ^ _42906;
  wire _42908 = _42904 ^ _42907;
  wire _42909 = _25108 ^ _977;
  wire _42910 = _42909 ^ _986;
  wire _42911 = _20030 ^ _27716;
  wire _42912 = _11428 ^ _15159;
  wire _42913 = _42911 ^ _42912;
  wire _42914 = _42910 ^ _42913;
  wire _42915 = _42908 ^ _42914;
  wire _42916 = uncoded_block[291] ^ uncoded_block[295];
  wire _42917 = _42916 ^ _10312;
  wire _42918 = _42917 ^ _33947;
  wire _42919 = _21017 ^ _16648;
  wire _42920 = _42919 ^ _6851;
  wire _42921 = _42918 ^ _42920;
  wire _42922 = _9780 ^ _9782;
  wire _42923 = _8063 ^ _4126;
  wire _42924 = _42922 ^ _42923;
  wire _42925 = _1825 ^ _11450;
  wire _42926 = _4845 ^ _11455;
  wire _42927 = _42925 ^ _42926;
  wire _42928 = _42924 ^ _42927;
  wire _42929 = _42921 ^ _42928;
  wire _42930 = _42915 ^ _42929;
  wire _42931 = _21497 ^ _6228;
  wire _42932 = _26032 ^ _1835;
  wire _42933 = _42931 ^ _42932;
  wire _42934 = _169 ^ _6874;
  wire _42935 = _12538 ^ _4858;
  wire _42936 = _42934 ^ _42935;
  wire _42937 = _42933 ^ _42936;
  wire _42938 = uncoded_block[386] ^ uncoded_block[393];
  wire _42939 = _42938 ^ _1847;
  wire _42940 = _10910 ^ _181;
  wire _42941 = _42939 ^ _42940;
  wire _42942 = _183 ^ _12545;
  wire _42943 = _9265 ^ _19612;
  wire _42944 = _42942 ^ _42943;
  wire _42945 = _42941 ^ _42944;
  wire _42946 = _42937 ^ _42945;
  wire _42947 = uncoded_block[425] ^ uncoded_block[433];
  wire _42948 = _42947 ^ _9820;
  wire _42949 = _31457 ^ _42948;
  wire _42950 = _1863 ^ _4174;
  wire _42951 = uncoded_block[448] ^ uncoded_block[453];
  wire _42952 = _42951 ^ _4885;
  wire _42953 = _42950 ^ _42952;
  wire _42954 = _42949 ^ _42953;
  wire _42955 = _23356 ^ _38387;
  wire _42956 = _4188 ^ _12025;
  wire _42957 = _7513 ^ _15212;
  wire _42958 = _42956 ^ _42957;
  wire _42959 = _42955 ^ _42958;
  wire _42960 = _42954 ^ _42959;
  wire _42961 = _42946 ^ _42960;
  wire _42962 = _42930 ^ _42961;
  wire _42963 = _42902 ^ _42962;
  wire _42964 = _1090 ^ _6276;
  wire _42965 = uncoded_block[492] ^ uncoded_block[498];
  wire _42966 = _42965 ^ _3434;
  wire _42967 = _42964 ^ _42966;
  wire _42968 = _5611 ^ _6925;
  wire _42969 = _18201 ^ _42968;
  wire _42970 = _42967 ^ _42969;
  wire _42971 = _236 ^ _10947;
  wire _42972 = _16709 ^ _14716;
  wire _42973 = _42971 ^ _42972;
  wire _42974 = uncoded_block[530] ^ uncoded_block[540];
  wire _42975 = _42974 ^ _25173;
  wire _42976 = _8720 ^ _25631;
  wire _42977 = _42975 ^ _42976;
  wire _42978 = _42973 ^ _42977;
  wire _42979 = _42970 ^ _42978;
  wire _42980 = _24284 ^ _3464;
  wire _42981 = _3467 ^ _6309;
  wire _42982 = _42980 ^ _42981;
  wire _42983 = _13700 ^ _15747;
  wire _42984 = _24289 ^ _20116;
  wire _42985 = _42983 ^ _42984;
  wire _42986 = _42982 ^ _42985;
  wire _42987 = uncoded_block[596] ^ uncoded_block[601];
  wire _42988 = _8148 ^ _42987;
  wire _42989 = _42988 ^ _2711;
  wire _42990 = _277 ^ _8154;
  wire _42991 = _42990 ^ _12612;
  wire _42992 = _42989 ^ _42991;
  wire _42993 = _42986 ^ _42992;
  wire _42994 = _42979 ^ _42993;
  wire _42995 = _16738 ^ _10418;
  wire _42996 = _42995 ^ _5659;
  wire _42997 = _14745 ^ _28905;
  wire _42998 = _12624 ^ _14234;
  wire _42999 = _42997 ^ _42998;
  wire _43000 = _42996 ^ _42999;
  wire _43001 = _33190 ^ _26549;
  wire _43002 = _43001 ^ _19183;
  wire _43003 = _3516 ^ _2744;
  wire _43004 = _19185 ^ _27408;
  wire _43005 = _43003 ^ _43004;
  wire _43006 = _43002 ^ _43005;
  wire _43007 = _43000 ^ _43006;
  wire _43008 = _321 ^ _18249;
  wire _43009 = _2754 ^ _6985;
  wire _43010 = _43008 ^ _43009;
  wire _43011 = _2757 ^ _4990;
  wire _43012 = _43011 ^ _30217;
  wire _43013 = _43010 ^ _43012;
  wire _43014 = uncoded_block[709] ^ uncoded_block[713];
  wire _43015 = _43014 ^ _17266;
  wire _43016 = _6998 ^ _4286;
  wire _43017 = _43015 ^ _43016;
  wire _43018 = _1991 ^ _1995;
  wire _43019 = uncoded_block[740] ^ uncoded_block[744];
  wire _43020 = _7005 ^ _43019;
  wire _43021 = _43018 ^ _43020;
  wire _43022 = _43017 ^ _43021;
  wire _43023 = _43013 ^ _43022;
  wire _43024 = _43007 ^ _43023;
  wire _43025 = _42994 ^ _43024;
  wire _43026 = uncoded_block[751] ^ uncoded_block[757];
  wire _43027 = _2775 ^ _43026;
  wire _43028 = uncoded_block[761] ^ uncoded_block[770];
  wire _43029 = _43028 ^ _12114;
  wire _43030 = _43027 ^ _43029;
  wire _43031 = uncoded_block[784] ^ uncoded_block[788];
  wire _43032 = _38464 ^ _43031;
  wire _43033 = _41207 ^ _43032;
  wire _43034 = _43030 ^ _43033;
  wire _43035 = uncoded_block[792] ^ uncoded_block[798];
  wire _43036 = _43035 ^ _7029;
  wire _43037 = _43036 ^ _20175;
  wire _43038 = _390 ^ _392;
  wire _43039 = _10483 ^ _2808;
  wire _43040 = _43038 ^ _43039;
  wire _43041 = _43037 ^ _43040;
  wire _43042 = _43034 ^ _43041;
  wire _43043 = _12131 ^ _5051;
  wire _43044 = uncoded_block[825] ^ uncoded_block[831];
  wire _43045 = _43044 ^ _4331;
  wire _43046 = _43043 ^ _43045;
  wire _43047 = _401 ^ _21159;
  wire _43048 = _14812 ^ _19725;
  wire _43049 = _43047 ^ _43048;
  wire _43050 = _43046 ^ _43049;
  wire _43051 = _30680 ^ _15824;
  wire _43052 = _17303 ^ _43051;
  wire _43053 = _416 ^ _3608;
  wire _43054 = _19240 ^ _43053;
  wire _43055 = _43052 ^ _43054;
  wire _43056 = _43050 ^ _43055;
  wire _43057 = _43042 ^ _43056;
  wire _43058 = _2053 ^ _4352;
  wire _43059 = _10506 ^ _3616;
  wire _43060 = _43058 ^ _43059;
  wire _43061 = _3617 ^ _2065;
  wire _43062 = _3623 ^ _2070;
  wire _43063 = _43061 ^ _43062;
  wire _43064 = _43060 ^ _43063;
  wire _43065 = uncoded_block[913] ^ uncoded_block[921];
  wire _43066 = _19252 ^ _43065;
  wire _43067 = _31141 ^ _5773;
  wire _43068 = _43066 ^ _43067;
  wire _43069 = _15848 ^ _453;
  wire _43070 = _8271 ^ _29387;
  wire _43071 = _43069 ^ _43070;
  wire _43072 = _43068 ^ _43071;
  wire _43073 = _43064 ^ _43072;
  wire _43074 = _1303 ^ _2869;
  wire _43075 = _27478 ^ _12179;
  wire _43076 = _43074 ^ _43075;
  wire _43077 = _12180 ^ _8847;
  wire _43078 = _5112 ^ _16841;
  wire _43079 = _43077 ^ _43078;
  wire _43080 = _43076 ^ _43079;
  wire _43081 = uncoded_block[981] ^ uncoded_block[985];
  wire _43082 = _43081 ^ _1317;
  wire _43083 = _14850 ^ _4401;
  wire _43084 = _43082 ^ _43083;
  wire _43085 = uncoded_block[1005] ^ uncoded_block[1008];
  wire _43086 = _15858 ^ _43085;
  wire _43087 = _481 ^ _43086;
  wire _43088 = _43084 ^ _43087;
  wire _43089 = _43080 ^ _43088;
  wire _43090 = _43073 ^ _43089;
  wire _43091 = _43057 ^ _43090;
  wire _43092 = _43025 ^ _43091;
  wire _43093 = _42963 ^ _43092;
  wire _43094 = _25295 ^ _2891;
  wire _43095 = _1333 ^ _9998;
  wire _43096 = _43094 ^ _43095;
  wire _43097 = _18801 ^ _2898;
  wire _43098 = _2127 ^ _1342;
  wire _43099 = _43097 ^ _43098;
  wire _43100 = _43096 ^ _43099;
  wire _43101 = uncoded_block[1039] ^ uncoded_block[1044];
  wire _43102 = _2129 ^ _43101;
  wire _43103 = uncoded_block[1050] ^ uncoded_block[1058];
  wire _43104 = _29410 ^ _43103;
  wire _43105 = _43102 ^ _43104;
  wire _43106 = _35723 ^ _42736;
  wire _43107 = _5827 ^ _43106;
  wire _43108 = _43105 ^ _43107;
  wire _43109 = _43100 ^ _43108;
  wire _43110 = _533 ^ _22149;
  wire _43111 = _2930 ^ _11139;
  wire _43112 = _43110 ^ _43111;
  wire _43113 = _18365 ^ _34943;
  wire _43114 = _4450 ^ _8337;
  wire _43115 = _43113 ^ _43114;
  wire _43116 = _43112 ^ _43115;
  wire _43117 = uncoded_block[1118] ^ uncoded_block[1124];
  wire _43118 = _43117 ^ _18832;
  wire _43119 = _560 ^ _10591;
  wire _43120 = _43118 ^ _43119;
  wire _43121 = uncoded_block[1140] ^ uncoded_block[1145];
  wire _43122 = _10593 ^ _43121;
  wire _43123 = _43122 ^ _18379;
  wire _43124 = _43120 ^ _43123;
  wire _43125 = _43116 ^ _43124;
  wire _43126 = _43109 ^ _43125;
  wire _43127 = uncoded_block[1162] ^ uncoded_block[1168];
  wire _43128 = _578 ^ _43127;
  wire _43129 = _3729 ^ _43128;
  wire _43130 = _29033 ^ _35353;
  wire _43131 = _43129 ^ _43130;
  wire _43132 = _36573 ^ _1420;
  wire _43133 = _22179 ^ _8951;
  wire _43134 = _43132 ^ _43133;
  wire _43135 = uncoded_block[1199] ^ uncoded_block[1205];
  wire _43136 = _43135 ^ _2216;
  wire _43137 = _43136 ^ _33335;
  wire _43138 = _43134 ^ _43137;
  wire _43139 = _43131 ^ _43138;
  wire _43140 = _31643 ^ _4503;
  wire _43141 = uncoded_block[1233] ^ uncoded_block[1237];
  wire _43142 = _43141 ^ _2230;
  wire _43143 = _14411 ^ _43142;
  wire _43144 = _43140 ^ _43143;
  wire _43145 = uncoded_block[1241] ^ uncoded_block[1247];
  wire _43146 = _43145 ^ _2998;
  wire _43147 = _43146 ^ _24926;
  wire _43148 = _5235 ^ _3786;
  wire _43149 = _7179 ^ _5907;
  wire _43150 = _43148 ^ _43149;
  wire _43151 = _43147 ^ _43150;
  wire _43152 = _43144 ^ _43151;
  wire _43153 = _43139 ^ _43152;
  wire _43154 = _43126 ^ _43153;
  wire _43155 = _22202 ^ _38587;
  wire _43156 = _6564 ^ _16424;
  wire _43157 = _36597 ^ _43156;
  wire _43158 = _43155 ^ _43157;
  wire _43159 = _15462 ^ _6572;
  wire _43160 = _20314 ^ _5926;
  wire _43161 = _43159 ^ _43160;
  wire _43162 = _2265 ^ _4543;
  wire _43163 = _7201 ^ _1494;
  wire _43164 = _43162 ^ _43163;
  wire _43165 = _43161 ^ _43164;
  wire _43166 = _43158 ^ _43165;
  wire _43167 = _24036 ^ _1497;
  wire _43168 = _7815 ^ _5268;
  wire _43169 = _43167 ^ _43168;
  wire _43170 = _5938 ^ _6587;
  wire _43171 = _6588 ^ _7211;
  wire _43172 = _43170 ^ _43171;
  wire _43173 = _43169 ^ _43172;
  wire _43174 = _5281 ^ _11226;
  wire _43175 = _10669 ^ _3055;
  wire _43176 = _43174 ^ _43175;
  wire _43177 = _687 ^ _7222;
  wire _43178 = _43177 ^ _693;
  wire _43179 = _43176 ^ _43178;
  wire _43180 = _43173 ^ _43179;
  wire _43181 = _43166 ^ _43180;
  wire _43182 = _2296 ^ _2299;
  wire _43183 = _4578 ^ _28344;
  wire _43184 = _43182 ^ _43183;
  wire _43185 = _17461 ^ _4583;
  wire _43186 = uncoded_block[1420] ^ uncoded_block[1425];
  wire _43187 = _43186 ^ _2311;
  wire _43188 = _43185 ^ _43187;
  wire _43189 = _43184 ^ _43188;
  wire _43190 = uncoded_block[1433] ^ uncoded_block[1443];
  wire _43191 = _5299 ^ _43190;
  wire _43192 = _43191 ^ _39809;
  wire _43193 = _719 ^ _2329;
  wire _43194 = _5313 ^ _1550;
  wire _43195 = _43193 ^ _43194;
  wire _43196 = _43192 ^ _43195;
  wire _43197 = _43189 ^ _43196;
  wire _43198 = _9608 ^ _5316;
  wire _43199 = uncoded_block[1478] ^ uncoded_block[1483];
  wire _43200 = _43199 ^ _1563;
  wire _43201 = _43198 ^ _43200;
  wire _43202 = _3891 ^ _3894;
  wire _43203 = _9615 ^ _43202;
  wire _43204 = _43201 ^ _43203;
  wire _43205 = _38638 ^ _9053;
  wire _43206 = uncoded_block[1518] ^ uncoded_block[1523];
  wire _43207 = _43206 ^ _8473;
  wire _43208 = _43205 ^ _43207;
  wire _43209 = _4623 ^ _19900;
  wire _43210 = _3906 ^ _3128;
  wire _43211 = _43209 ^ _43210;
  wire _43212 = _43208 ^ _43211;
  wire _43213 = _43204 ^ _43212;
  wire _43214 = _43197 ^ _43213;
  wire _43215 = _43181 ^ _43214;
  wire _43216 = _43154 ^ _43215;
  wire _43217 = uncoded_block[1550] ^ uncoded_block[1555];
  wire _43218 = _7274 ^ _43217;
  wire _43219 = _31732 ^ _774;
  wire _43220 = _43218 ^ _43219;
  wire _43221 = _37871 ^ _7891;
  wire _43222 = _43221 ^ _17008;
  wire _43223 = _43220 ^ _43222;
  wire _43224 = _3921 ^ _32567;
  wire _43225 = _789 ^ _791;
  wire _43226 = _43224 ^ _43225;
  wire _43227 = _4654 ^ _6674;
  wire _43228 = _20406 ^ _7906;
  wire _43229 = _43227 ^ _43228;
  wire _43230 = _43226 ^ _43229;
  wire _43231 = _43223 ^ _43230;
  wire _43232 = _7297 ^ _3160;
  wire _43233 = _2400 ^ _2404;
  wire _43234 = _43232 ^ _43233;
  wire _43235 = _30885 ^ _9104;
  wire _43236 = _43234 ^ _43235;
  wire _43237 = _11311 ^ _14530;
  wire _43238 = _12389 ^ _822;
  wire _43239 = _43237 ^ _43238;
  wire _43240 = _7927 ^ _6058;
  wire _43241 = _43240 ^ _37095;
  wire _43242 = _43239 ^ _43241;
  wire _43243 = _43236 ^ _43242;
  wire _43244 = _43231 ^ _43243;
  wire _43245 = _2427 ^ _3967;
  wire _43246 = _43245 ^ _21393;
  wire _43247 = _1669 ^ _20436;
  wire _43248 = _20437 ^ _851;
  wire _43249 = _43247 ^ _43248;
  wire _43250 = _43246 ^ _43249;
  wire _43251 = _22316 ^ _2441;
  wire _43252 = _43251 ^ _14033;
  wire _43253 = _43250 ^ _43252;
  wire _43254 = _43244 ^ _43253;
  wire _43255 = _43216 ^ _43254;
  wire _43256 = _43093 ^ _43255;
  wire _43257 = _21407 ^ _3;
  wire _43258 = _17559 ^ _871;
  wire _43259 = _43257 ^ _43258;
  wire _43260 = uncoded_block[19] ^ uncoded_block[23];
  wire _43261 = _43260 ^ _9694;
  wire _43262 = _43261 ^ _22792;
  wire _43263 = _43259 ^ _43262;
  wire _43264 = _4723 ^ _6101;
  wire _43265 = _7963 ^ _43264;
  wire _43266 = uncoded_block[52] ^ uncoded_block[57];
  wire _43267 = _43266 ^ _1705;
  wire _43268 = _34 ^ _2480;
  wire _43269 = _43267 ^ _43268;
  wire _43270 = _43265 ^ _43269;
  wire _43271 = _43263 ^ _43270;
  wire _43272 = _1712 ^ _2481;
  wire _43273 = _14586 ^ _2484;
  wire _43274 = _43272 ^ _43273;
  wire _43275 = _12447 ^ _4031;
  wire _43276 = _25066 ^ _43275;
  wire _43277 = _43274 ^ _43276;
  wire _43278 = uncoded_block[112] ^ uncoded_block[115];
  wire _43279 = _5453 ^ _43278;
  wire _43280 = _43279 ^ _11372;
  wire _43281 = _56 ^ _2502;
  wire _43282 = _43281 ^ _33065;
  wire _43283 = _43280 ^ _43282;
  wire _43284 = _43277 ^ _43283;
  wire _43285 = _43271 ^ _43284;
  wire _43286 = _17595 ^ _35892;
  wire _43287 = _73 ^ _15118;
  wire _43288 = _20489 ^ _43287;
  wire _43289 = _43286 ^ _43288;
  wire _43290 = _19536 ^ _1752;
  wire _43291 = _43290 ^ _14615;
  wire _43292 = _8009 ^ _4776;
  wire _43293 = _43292 ^ _6802;
  wire _43294 = _43291 ^ _43293;
  wire _43295 = _43289 ^ _43294;
  wire _43296 = _14622 ^ _8021;
  wire _43297 = _9750 ^ _4074;
  wire _43298 = _43296 ^ _43297;
  wire _43299 = _11409 ^ _6814;
  wire _43300 = uncoded_block[237] ^ uncoded_block[245];
  wire _43301 = _6821 ^ _43300;
  wire _43302 = _43299 ^ _43301;
  wire _43303 = _43298 ^ _43302;
  wire _43304 = _1785 ^ _3311;
  wire _43305 = _31828 ^ _43304;
  wire _43306 = _14639 ^ _10297;
  wire _43307 = uncoded_block[266] ^ uncoded_block[271];
  wire _43308 = _43307 ^ _3321;
  wire _43309 = _43306 ^ _43308;
  wire _43310 = _43305 ^ _43309;
  wire _43311 = _43303 ^ _43310;
  wire _43312 = _43295 ^ _43311;
  wire _43313 = _43285 ^ _43312;
  wire _43314 = _1795 ^ _7445;
  wire _43315 = _43314 ^ _13065;
  wire _43316 = _5522 ^ _4819;
  wire _43317 = _43316 ^ _20039;
  wire _43318 = _43315 ^ _43317;
  wire _43319 = _34745 ^ _3339;
  wire _43320 = _27726 ^ _16152;
  wire _43321 = _43319 ^ _43320;
  wire _43322 = _43318 ^ _43321;
  wire _43323 = _4125 ^ _5536;
  wire _43324 = _10320 ^ _43323;
  wire _43325 = _2592 ^ _6217;
  wire _43326 = _43325 ^ _3356;
  wire _43327 = _43324 ^ _43326;
  wire _43328 = uncoded_block[348] ^ uncoded_block[354];
  wire _43329 = _43328 ^ _15686;
  wire _43330 = _17163 ^ _1838;
  wire _43331 = _43329 ^ _43330;
  wire _43332 = _3375 ^ _1038;
  wire _43333 = _2613 ^ _4151;
  wire _43334 = _43332 ^ _43333;
  wire _43335 = _43331 ^ _43334;
  wire _43336 = _43327 ^ _43335;
  wire _43337 = _43322 ^ _43336;
  wire _43338 = _6881 ^ _5559;
  wire _43339 = uncoded_block[407] ^ uncoded_block[412];
  wire _43340 = _12545 ^ _43339;
  wire _43341 = _43338 ^ _43340;
  wire _43342 = _6250 ^ _17676;
  wire _43343 = _43341 ^ _43342;
  wire _43344 = _40377 ^ _2641;
  wire _43345 = _43344 ^ _13123;
  wire _43346 = _11486 ^ _3411;
  wire _43347 = _2650 ^ _6264;
  wire _43348 = _43346 ^ _43347;
  wire _43349 = _43345 ^ _43348;
  wire _43350 = _43343 ^ _43349;
  wire _43351 = _13662 ^ _1079;
  wire _43352 = _24721 ^ _5592;
  wire _43353 = _43351 ^ _43352;
  wire _43354 = _4194 ^ _2664;
  wire _43355 = _9831 ^ _43354;
  wire _43356 = _43353 ^ _43355;
  wire _43357 = uncoded_block[493] ^ uncoded_block[498];
  wire _43358 = _43357 ^ _6279;
  wire _43359 = _43358 ^ _13675;
  wire _43360 = _17694 ^ _13676;
  wire _43361 = _43360 ^ _42315;
  wire _43362 = _43359 ^ _43361;
  wire _43363 = _43356 ^ _43362;
  wire _43364 = _43350 ^ _43363;
  wire _43365 = _43337 ^ _43364;
  wire _43366 = _43313 ^ _43365;
  wire _43367 = _1108 ^ _38815;
  wire _43368 = _1114 ^ _21550;
  wire _43369 = _43367 ^ _43368;
  wire _43370 = _9854 ^ _1118;
  wire _43371 = _3459 ^ _25631;
  wire _43372 = _43370 ^ _43371;
  wire _43373 = _43369 ^ _43372;
  wire _43374 = _3461 ^ _258;
  wire _43375 = _18682 ^ _1130;
  wire _43376 = _43374 ^ _43375;
  wire _43377 = _19652 ^ _6947;
  wire _43378 = uncoded_block[587] ^ uncoded_block[593];
  wire _43379 = _8733 ^ _43378;
  wire _43380 = _43377 ^ _43379;
  wire _43381 = _43376 ^ _43380;
  wire _43382 = _43373 ^ _43381;
  wire _43383 = _2707 ^ _9868;
  wire _43384 = _17722 ^ _43383;
  wire _43385 = _14218 ^ _16233;
  wire _43386 = _43385 ^ _16237;
  wire _43387 = _43384 ^ _43386;
  wire _43388 = _15261 ^ _12071;
  wire _43389 = _34421 ^ _43388;
  wire _43390 = _22028 ^ _22479;
  wire _43391 = _4972 ^ _6341;
  wire _43392 = _43390 ^ _43391;
  wire _43393 = _43389 ^ _43392;
  wire _43394 = _43387 ^ _43393;
  wire _43395 = _43382 ^ _43394;
  wire _43396 = _22958 ^ _3514;
  wire _43397 = _43396 ^ _310;
  wire _43398 = _1174 ^ _16752;
  wire _43399 = _43398 ^ _21587;
  wire _43400 = _43397 ^ _43399;
  wire _43401 = _8184 ^ _8186;
  wire _43402 = _3528 ^ _43401;
  wire _43403 = _10445 ^ _3533;
  wire _43404 = uncoded_block[712] ^ uncoded_block[717];
  wire _43405 = _33204 ^ _43404;
  wire _43406 = _43403 ^ _43405;
  wire _43407 = _43402 ^ _43406;
  wire _43408 = _43400 ^ _43407;
  wire _43409 = _20147 ^ _20152;
  wire _43410 = uncoded_block[740] ^ uncoded_block[746];
  wire _43411 = _1206 ^ _43410;
  wire _43412 = _19205 ^ _43411;
  wire _43413 = _43409 ^ _43412;
  wire _43414 = uncoded_block[756] ^ uncoded_block[759];
  wire _43415 = _43414 ^ _9914;
  wire _43416 = _13210 ^ _43415;
  wire _43417 = uncoded_block[762] ^ uncoded_block[767];
  wire _43418 = _43417 ^ _1218;
  wire _43419 = _1221 ^ _19705;
  wire _43420 = _43418 ^ _43419;
  wire _43421 = _43416 ^ _43420;
  wire _43422 = _43413 ^ _43421;
  wire _43423 = _43408 ^ _43422;
  wire _43424 = _43395 ^ _43423;
  wire _43425 = uncoded_block[788] ^ uncoded_block[793];
  wire _43426 = _43425 ^ _1233;
  wire _43427 = _35262 ^ _43426;
  wire _43428 = _8224 ^ _9394;
  wire _43429 = _43428 ^ _17790;
  wire _43430 = _43427 ^ _43429;
  wire _43431 = _2029 ^ _5052;
  wire _43432 = _33655 ^ _43431;
  wire _43433 = _33659 ^ _8808;
  wire _43434 = _2820 ^ _7643;
  wire _43435 = _43433 ^ _43434;
  wire _43436 = _43432 ^ _43435;
  wire _43437 = _43430 ^ _43436;
  wire _43438 = _12146 ^ _3600;
  wire _43439 = _408 ^ _2824;
  wire _43440 = _43438 ^ _43439;
  wire _43441 = _414 ^ _416;
  wire _43442 = _6416 ^ _16815;
  wire _43443 = _43441 ^ _43442;
  wire _43444 = _43440 ^ _43443;
  wire _43445 = _3615 ^ _31575;
  wire _43446 = _18311 ^ _6428;
  wire _43447 = _3625 ^ _23917;
  wire _43448 = _43446 ^ _43447;
  wire _43449 = _43445 ^ _43448;
  wire _43450 = _43444 ^ _43449;
  wire _43451 = _43437 ^ _43450;
  wire _43452 = _17821 ^ _28972;
  wire _43453 = _448 ^ _24837;
  wire _43454 = uncoded_block[939] ^ uncoded_block[946];
  wire _43455 = _43454 ^ _9975;
  wire _43456 = _43453 ^ _43455;
  wire _43457 = _43452 ^ _43456;
  wire _43458 = _13266 ^ _5779;
  wire _43459 = _43458 ^ _34095;
  wire _43460 = _12180 ^ _11648;
  wire _43461 = _8281 ^ _43460;
  wire _43462 = _43459 ^ _43461;
  wire _43463 = _43457 ^ _43462;
  wire _43464 = _38915 ^ _28980;
  wire _43465 = _43464 ^ _22117;
  wire _43466 = _2882 ^ _17340;
  wire _43467 = _43466 ^ _28609;
  wire _43468 = _43465 ^ _43467;
  wire _43469 = uncoded_block[1006] ^ uncoded_block[1014];
  wire _43470 = _43469 ^ _7108;
  wire _43471 = _43470 ^ _2897;
  wire _43472 = _8875 ^ _499;
  wire _43473 = _2127 ^ _2129;
  wire _43474 = _43472 ^ _43473;
  wire _43475 = _43471 ^ _43474;
  wire _43476 = _43468 ^ _43475;
  wire _43477 = _43463 ^ _43476;
  wire _43478 = _43451 ^ _43477;
  wire _43479 = _43424 ^ _43478;
  wire _43480 = _43366 ^ _43479;
  wire _43481 = _1346 ^ _2910;
  wire _43482 = _43481 ^ _5815;
  wire _43483 = _4430 ^ _7117;
  wire _43484 = _36543 ^ _1366;
  wire _43485 = _43483 ^ _43484;
  wire _43486 = _43482 ^ _43485;
  wire _43487 = uncoded_block[1077] ^ uncoded_block[1084];
  wire _43488 = _11125 ^ _43487;
  wire _43489 = _12774 ^ _3698;
  wire _43490 = _43488 ^ _43489;
  wire _43491 = _5843 ^ _8910;
  wire _43492 = _8914 ^ _13319;
  wire _43493 = _43491 ^ _43492;
  wire _43494 = _43490 ^ _43493;
  wire _43495 = _43486 ^ _43494;
  wire _43496 = _32873 ^ _12789;
  wire _43497 = _15894 ^ _560;
  wire _43498 = _43496 ^ _43497;
  wire _43499 = _10591 ^ _20266;
  wire _43500 = _8930 ^ _2179;
  wire _43501 = _43499 ^ _43500;
  wire _43502 = _43498 ^ _43501;
  wire _43503 = _8351 ^ _3727;
  wire _43504 = _18379 ^ _43503;
  wire _43505 = _23988 ^ _35744;
  wire _43506 = _43504 ^ _43505;
  wire _43507 = _43502 ^ _43506;
  wire _43508 = _43495 ^ _43507;
  wire _43509 = _40155 ^ _2197;
  wire _43510 = uncoded_block[1188] ^ uncoded_block[1193];
  wire _43511 = _43510 ^ _12810;
  wire _43512 = _8370 ^ _4491;
  wire _43513 = _43511 ^ _43512;
  wire _43514 = _43509 ^ _43513;
  wire _43515 = _2217 ^ _12259;
  wire _43516 = _2219 ^ _14407;
  wire _43517 = _43515 ^ _43516;
  wire _43518 = _6532 ^ _5894;
  wire _43519 = _5219 ^ _15927;
  wire _43520 = _43518 ^ _43519;
  wire _43521 = _43517 ^ _43520;
  wire _43522 = _43514 ^ _43521;
  wire _43523 = uncoded_block[1249] ^ uncoded_block[1253];
  wire _43524 = _37796 ^ _43523;
  wire _43525 = _26706 ^ _43524;
  wire _43526 = _29054 ^ _24016;
  wire _43527 = _43525 ^ _43526;
  wire _43528 = _25826 ^ _7183;
  wire _43529 = _25824 ^ _43528;
  wire _43530 = _4525 ^ _3797;
  wire _43531 = _11195 ^ _3800;
  wire _43532 = _43530 ^ _43531;
  wire _43533 = _43529 ^ _43532;
  wire _43534 = _43527 ^ _43533;
  wire _43535 = _43522 ^ _43534;
  wire _43536 = _43508 ^ _43535;
  wire _43537 = _7193 ^ _6564;
  wire _43538 = uncoded_block[1301] ^ uncoded_block[1305];
  wire _43539 = _43538 ^ _2259;
  wire _43540 = _43537 ^ _43539;
  wire _43541 = _9552 ^ _9555;
  wire _43542 = _24033 ^ _43541;
  wire _43543 = _43540 ^ _43542;
  wire _43544 = _3814 ^ _16435;
  wire _43545 = _43544 ^ _18884;
  wire _43546 = _2277 ^ _11215;
  wire _43547 = _5268 ^ _16942;
  wire _43548 = _43546 ^ _43547;
  wire _43549 = _43545 ^ _43548;
  wire _43550 = _43543 ^ _43549;
  wire _43551 = _5940 ^ _32106;
  wire _43552 = _43551 ^ _13934;
  wire _43553 = _29496 ^ _3834;
  wire _43554 = _43553 ^ _35406;
  wire _43555 = _43552 ^ _43554;
  wire _43556 = _13412 ^ _5952;
  wire _43557 = _3065 ^ _4572;
  wire _43558 = _43556 ^ _43557;
  wire _43559 = _14968 ^ _9585;
  wire _43560 = _30395 ^ _43559;
  wire _43561 = _43558 ^ _43560;
  wire _43562 = _43555 ^ _43561;
  wire _43563 = _43550 ^ _43562;
  wire _43564 = _22237 ^ _3850;
  wire _43565 = _9022 ^ _11239;
  wire _43566 = _43564 ^ _43565;
  wire _43567 = _24065 ^ _38626;
  wire _43568 = _16963 ^ _43567;
  wire _43569 = _43566 ^ _43568;
  wire _43570 = _5976 ^ _11247;
  wire _43571 = _13437 ^ _24070;
  wire _43572 = _43570 ^ _43571;
  wire _43573 = _7247 ^ _16977;
  wire _43574 = _43573 ^ _34616;
  wire _43575 = _43572 ^ _43574;
  wire _43576 = _43569 ^ _43575;
  wire _43577 = _7861 ^ _1563;
  wire _43578 = _43577 ^ _16483;
  wire _43579 = _14484 ^ _41762;
  wire _43580 = _43579 ^ _35038;
  wire _43581 = _43578 ^ _43580;
  wire _43582 = _9621 ^ _4620;
  wire _43583 = _43582 ^ _16991;
  wire _43584 = _32975 ^ _6012;
  wire _43585 = _3907 ^ _43584;
  wire _43586 = _43583 ^ _43585;
  wire _43587 = _43581 ^ _43586;
  wire _43588 = _43576 ^ _43587;
  wire _43589 = _43563 ^ _43588;
  wire _43590 = _43536 ^ _43589;
  wire _43591 = _6013 ^ _15020;
  wire _43592 = _6016 ^ _26794;
  wire _43593 = _43591 ^ _43592;
  wire _43594 = uncoded_block[1564] ^ uncoded_block[1576];
  wire _43595 = _43594 ^ _3921;
  wire _43596 = _784 ^ _19918;
  wire _43597 = _43595 ^ _43596;
  wire _43598 = _43593 ^ _43597;
  wire _43599 = _791 ^ _3933;
  wire _43600 = _43599 ^ _15543;
  wire _43601 = _3153 ^ _1627;
  wire _43602 = _43601 ^ _2399;
  wire _43603 = _43600 ^ _43602;
  wire _43604 = _43598 ^ _43603;
  wire _43605 = _27215 ^ _10185;
  wire _43606 = _14525 ^ _6048;
  wire _43607 = _43605 ^ _43606;
  wire _43608 = _2405 ^ _5392;
  wire _43609 = _43608 ^ _36683;
  wire _43610 = _43607 ^ _43609;
  wire _43611 = _816 ^ _6691;
  wire _43612 = uncoded_block[1661] ^ uncoded_block[1669];
  wire _43613 = _820 ^ _43612;
  wire _43614 = _43611 ^ _43613;
  wire _43615 = _3182 ^ _17537;
  wire _43616 = _43615 ^ _22766;
  wire _43617 = _43614 ^ _43616;
  wire _43618 = _43610 ^ _43617;
  wire _43619 = _43604 ^ _43618;
  wire _43620 = _24130 ^ _3967;
  wire _43621 = _840 ^ _3975;
  wire _43622 = _43620 ^ _43621;
  wire _43623 = _20437 ^ _2437;
  wire _43624 = _43623 ^ _26373;
  wire _43625 = _43622 ^ _43624;
  wire _43626 = _43625 ^ uncoded_block[1722];
  wire _43627 = _43619 ^ _43626;
  wire _43628 = _43590 ^ _43627;
  wire _43629 = _43480 ^ _43628;
  wire _43630 = _17559 ^ _868;
  wire _43631 = _21408 ^ _43630;
  wire _43632 = _4000 ^ _14565;
  wire _43633 = _4718 ^ _2466;
  wire _43634 = _43632 ^ _43633;
  wire _43635 = _43631 ^ _43634;
  wire _43636 = _19503 ^ _20464;
  wire _43637 = _1703 ^ _10801;
  wire _43638 = _35 ^ _12438;
  wire _43639 = _43637 ^ _43638;
  wire _43640 = _43636 ^ _43639;
  wire _43641 = _43635 ^ _43640;
  wire _43642 = _2484 ^ _1718;
  wire _43643 = _39111 ^ _43642;
  wire _43644 = _15097 ^ _7986;
  wire _43645 = _22809 ^ _43644;
  wire _43646 = _43643 ^ _43645;
  wire _43647 = uncoded_block[110] ^ uncoded_block[114];
  wire _43648 = _911 ^ _43647;
  wire _43649 = uncoded_block[123] ^ uncoded_block[133];
  wire _43650 = _33056 ^ _43649;
  wire _43651 = _43648 ^ _43650;
  wire _43652 = _926 ^ _1736;
  wire _43653 = _39910 ^ _15114;
  wire _43654 = _43652 ^ _43653;
  wire _43655 = _43651 ^ _43654;
  wire _43656 = _43646 ^ _43655;
  wire _43657 = _43641 ^ _43656;
  wire _43658 = uncoded_block[146] ^ uncoded_block[155];
  wire _43659 = _43658 ^ _73;
  wire _43660 = _19040 ^ _1749;
  wire _43661 = _43659 ^ _43660;
  wire _43662 = _6787 ^ _42888;
  wire _43663 = _20979 ^ _7403;
  wire _43664 = _43662 ^ _43663;
  wire _43665 = _43661 ^ _43664;
  wire _43666 = _5479 ^ _945;
  wire _43667 = _19544 ^ _17112;
  wire _43668 = _43666 ^ _43667;
  wire _43669 = _1764 ^ _8600;
  wire _43670 = uncoded_block[218] ^ uncoded_block[232];
  wire _43671 = _6161 ^ _43670;
  wire _43672 = _43669 ^ _43671;
  wire _43673 = _43668 ^ _43672;
  wire _43674 = _43665 ^ _43673;
  wire _43675 = _6822 ^ _10292;
  wire _43676 = _5503 ^ _11952;
  wire _43677 = _43675 ^ _43676;
  wire _43678 = _8034 ^ _20999;
  wire _43679 = _43678 ^ _24671;
  wire _43680 = _43677 ^ _43679;
  wire _43681 = uncoded_block[276] ^ uncoded_block[280];
  wire _43682 = _3321 ^ _43681;
  wire _43683 = _7442 ^ _43682;
  wire _43684 = _33522 ^ _9772;
  wire _43685 = _994 ^ _2573;
  wire _43686 = _43684 ^ _43685;
  wire _43687 = _43683 ^ _43686;
  wire _43688 = _43680 ^ _43687;
  wire _43689 = _43674 ^ _43688;
  wire _43690 = _43657 ^ _43689;
  wire _43691 = uncoded_block[300] ^ uncoded_block[305];
  wire _43692 = _17142 ^ _43691;
  wire _43693 = _20536 ^ _3338;
  wire _43694 = _43692 ^ _43693;
  wire _43695 = _17642 ^ _6208;
  wire _43696 = _43695 ^ _21021;
  wire _43697 = _43694 ^ _43696;
  wire _43698 = _34751 ^ _7463;
  wire _43699 = _43698 ^ _22408;
  wire _43700 = _18621 ^ _14662;
  wire _43701 = _8069 ^ _3362;
  wire _43702 = _43700 ^ _43701;
  wire _43703 = _43699 ^ _43702;
  wire _43704 = _43697 ^ _43703;
  wire _43705 = uncoded_block[363] ^ uncoded_block[368];
  wire _43706 = _6228 ^ _43705;
  wire _43707 = _13094 ^ _28838;
  wire _43708 = _43706 ^ _43707;
  wire _43709 = uncoded_block[379] ^ uncoded_block[384];
  wire _43710 = _43709 ^ _18633;
  wire _43711 = _9806 ^ _181;
  wire _43712 = _43710 ^ _43711;
  wire _43713 = _43708 ^ _43712;
  wire _43714 = _6244 ^ _2629;
  wire _43715 = _3394 ^ _193;
  wire _43716 = _43714 ^ _43715;
  wire _43717 = uncoded_block[419] ^ uncoded_block[424];
  wire _43718 = _43717 ^ _8672;
  wire _43719 = _6894 ^ _13117;
  wire _43720 = _43718 ^ _43719;
  wire _43721 = _43716 ^ _43720;
  wire _43722 = _43713 ^ _43721;
  wire _43723 = _43704 ^ _43722;
  wire _43724 = _22903 ^ _26495;
  wire _43725 = _31460 ^ _43724;
  wire _43726 = _8105 ^ _23357;
  wire _43727 = _1879 ^ _2657;
  wire _43728 = _43726 ^ _43727;
  wire _43729 = _43725 ^ _43728;
  wire _43730 = _21526 ^ _39989;
  wire _43731 = _1091 ^ _34785;
  wire _43732 = _43730 ^ _43731;
  wire _43733 = _5606 ^ _2671;
  wire _43734 = _43733 ^ _27370;
  wire _43735 = _43732 ^ _43734;
  wire _43736 = _43729 ^ _43735;
  wire _43737 = _4208 ^ _1108;
  wire _43738 = _26514 ^ _1905;
  wire _43739 = _43737 ^ _43738;
  wire _43740 = _5620 ^ _1909;
  wire _43741 = uncoded_block[550] ^ uncoded_block[555];
  wire _43742 = _43741 ^ _1123;
  wire _43743 = _43740 ^ _43742;
  wire _43744 = _43739 ^ _43743;
  wire _43745 = uncoded_block[562] ^ uncoded_block[572];
  wire _43746 = _24284 ^ _43745;
  wire _43747 = _43746 ^ _8732;
  wire _43748 = uncoded_block[589] ^ uncoded_block[595];
  wire _43749 = _35220 ^ _43748;
  wire _43750 = _2706 ^ _7558;
  wire _43751 = _43749 ^ _43750;
  wire _43752 = _43747 ^ _43751;
  wire _43753 = _43744 ^ _43752;
  wire _43754 = _43736 ^ _43753;
  wire _43755 = _43723 ^ _43754;
  wire _43756 = _43690 ^ _43755;
  wire _43757 = _1146 ^ _6323;
  wire _43758 = _43757 ^ _16237;
  wire _43759 = uncoded_block[614] ^ uncoded_block[621];
  wire _43760 = _43759 ^ _10418;
  wire _43761 = uncoded_block[630] ^ uncoded_block[635];
  wire _43762 = _287 ^ _43761;
  wire _43763 = _43760 ^ _43762;
  wire _43764 = _43758 ^ _43763;
  wire _43765 = _4249 ^ _6335;
  wire _43766 = _4256 ^ _34028;
  wire _43767 = _43765 ^ _43766;
  wire _43768 = _304 ^ _8172;
  wire _43769 = _43768 ^ _2743;
  wire _43770 = _43767 ^ _43769;
  wire _43771 = _43764 ^ _43770;
  wire _43772 = uncoded_block[671] ^ uncoded_block[675];
  wire _43773 = _1174 ^ _43772;
  wire _43774 = _23410 ^ _1971;
  wire _43775 = _43773 ^ _43774;
  wire _43776 = _8767 ^ _4989;
  wire _43777 = _18721 ^ _23863;
  wire _43778 = _43776 ^ _43777;
  wire _43779 = _43775 ^ _43778;
  wire _43780 = _13742 ^ _5690;
  wire _43781 = _343 ^ _1988;
  wire _43782 = _43780 ^ _43781;
  wire _43783 = _1990 ^ _349;
  wire _43784 = _37678 ^ _4289;
  wire _43785 = _43783 ^ _43784;
  wire _43786 = _43782 ^ _43785;
  wire _43787 = _43779 ^ _43786;
  wire _43788 = _43771 ^ _43787;
  wire _43789 = _5704 ^ _40817;
  wire _43790 = _42365 ^ _43789;
  wire _43791 = _11012 ^ _17774;
  wire _43792 = uncoded_block[762] ^ uncoded_block[766];
  wire _43793 = _43792 ^ _30234;
  wire _43794 = _43791 ^ _43793;
  wire _43795 = _43790 ^ _43794;
  wire _43796 = _2792 ^ _3567;
  wire _43797 = _3568 ^ _14793;
  wire _43798 = _43796 ^ _43797;
  wire _43799 = _11024 ^ _382;
  wire _43800 = _29780 ^ _43799;
  wire _43801 = _43798 ^ _43800;
  wire _43802 = _43795 ^ _43801;
  wire _43803 = _9928 ^ _3577;
  wire _43804 = _392 ^ _11597;
  wire _43805 = _43803 ^ _43804;
  wire _43806 = _2029 ^ _14290;
  wire _43807 = _43806 ^ _16799;
  wire _43808 = _43805 ^ _43807;
  wire _43809 = _27846 ^ _2035;
  wire _43810 = _10495 ^ _3599;
  wire _43811 = _43809 ^ _43810;
  wire _43812 = _7643 ^ _2821;
  wire _43813 = _7049 ^ _6410;
  wire _43814 = _43812 ^ _43813;
  wire _43815 = _43811 ^ _43814;
  wire _43816 = _43808 ^ _43815;
  wire _43817 = _43802 ^ _43816;
  wire _43818 = _43788 ^ _43817;
  wire _43819 = _9949 ^ _5071;
  wire _43820 = uncoded_block[876] ^ uncoded_block[882];
  wire _43821 = _33671 ^ _43820;
  wire _43822 = _43819 ^ _43821;
  wire _43823 = _4352 ^ _3614;
  wire _43824 = _8826 ^ _28965;
  wire _43825 = _43823 ^ _43824;
  wire _43826 = _43822 ^ _43825;
  wire _43827 = uncoded_block[909] ^ uncoded_block[913];
  wire _43828 = _43827 ^ _17818;
  wire _43829 = _15350 ^ _39692;
  wire _43830 = _43828 ^ _43829;
  wire _43831 = _31141 ^ _1296;
  wire _43832 = _3637 ^ _452;
  wire _43833 = _43831 ^ _43832;
  wire _43834 = _43830 ^ _43833;
  wire _43835 = _43826 ^ _43834;
  wire _43836 = _2865 ^ _456;
  wire _43837 = _3643 ^ _6441;
  wire _43838 = _43836 ^ _43837;
  wire _43839 = _464 ^ _5785;
  wire _43840 = _43839 ^ _1316;
  wire _43841 = _43838 ^ _43840;
  wire _43842 = uncoded_block[975] ^ uncoded_block[979];
  wire _43843 = _43842 ^ _29832;
  wire _43844 = uncoded_block[986] ^ uncoded_block[990];
  wire _43845 = _7093 ^ _43844;
  wire _43846 = _43843 ^ _43845;
  wire _43847 = _3663 ^ _28985;
  wire _43848 = uncoded_block[999] ^ uncoded_block[1004];
  wire _43849 = _43848 ^ _43085;
  wire _43850 = _43847 ^ _43849;
  wire _43851 = _43846 ^ _43850;
  wire _43852 = _43841 ^ _43851;
  wire _43853 = _43835 ^ _43852;
  wire _43854 = _2894 ^ _8872;
  wire _43855 = _35316 ^ _43854;
  wire _43856 = _35710 ^ _1345;
  wire _43857 = _38937 ^ _23964;
  wire _43858 = _43856 ^ _43857;
  wire _43859 = _43855 ^ _43858;
  wire _43860 = _1364 ^ _2143;
  wire _43861 = _23967 ^ _43860;
  wire _43862 = _529 ^ _8895;
  wire _43863 = _40877 ^ _1374;
  wire _43864 = _43862 ^ _43863;
  wire _43865 = _43861 ^ _43864;
  wire _43866 = _43859 ^ _43865;
  wire _43867 = _10021 ^ _7129;
  wire _43868 = _43867 ^ _32869;
  wire _43869 = _15407 ^ _3713;
  wire _43870 = _8916 ^ _43869;
  wire _43871 = _43868 ^ _43870;
  wire _43872 = _16377 ^ _35737;
  wire _43873 = _5856 ^ _35343;
  wire _43874 = uncoded_block[1146] ^ uncoded_block[1151];
  wire _43875 = uncoded_block[1157] ^ uncoded_block[1163];
  wire _43876 = _43874 ^ _43875;
  wire _43877 = _43873 ^ _43876;
  wire _43878 = _43872 ^ _43877;
  wire _43879 = _43871 ^ _43878;
  wire _43880 = _43866 ^ _43879;
  wire _43881 = _43853 ^ _43880;
  wire _43882 = _43818 ^ _43881;
  wire _43883 = _43756 ^ _43882;
  wire _43884 = uncoded_block[1172] ^ uncoded_block[1177];
  wire _43885 = _30756 ^ _43884;
  wire _43886 = _6519 ^ _590;
  wire _43887 = _43885 ^ _43886;
  wire _43888 = _35354 ^ _5203;
  wire _43889 = _24910 ^ _1421;
  wire _43890 = _43888 ^ _43889;
  wire _43891 = _43887 ^ _43890;
  wire _43892 = _22183 ^ _1428;
  wire _43893 = _17901 ^ _43892;
  wire _43894 = _605 ^ _4499;
  wire _43895 = _13355 ^ _612;
  wire _43896 = _43894 ^ _43895;
  wire _43897 = _43893 ^ _43896;
  wire _43898 = _43891 ^ _43897;
  wire _43899 = _1440 ^ _15441;
  wire _43900 = _620 ^ _4511;
  wire _43901 = _43899 ^ _43900;
  wire _43902 = _8968 ^ _7780;
  wire _43903 = _43902 ^ _42769;
  wire _43904 = _43901 ^ _43903;
  wire _43905 = _1458 ^ _3008;
  wire _43906 = _628 ^ _30789;
  wire _43907 = _43905 ^ _43906;
  wire _43908 = _3794 ^ _5243;
  wire _43909 = _13380 ^ _1469;
  wire _43910 = _43908 ^ _43909;
  wire _43911 = _43907 ^ _43910;
  wire _43912 = _43904 ^ _43911;
  wire _43913 = _43898 ^ _43912;
  wire _43914 = uncoded_block[1294] ^ uncoded_block[1300];
  wire _43915 = _43914 ^ _16424;
  wire _43916 = _8992 ^ _2261;
  wire _43917 = _43915 ^ _43916;
  wire _43918 = _7201 ^ _5931;
  wire _43919 = _37012 ^ _43918;
  wire _43920 = _43917 ^ _43919;
  wire _43921 = _4551 ^ _4553;
  wire _43922 = _7815 ^ _664;
  wire _43923 = _43921 ^ _43922;
  wire _43924 = _15473 ^ _4559;
  wire _43925 = _7211 ^ _2284;
  wire _43926 = _43924 ^ _43925;
  wire _43927 = _43923 ^ _43926;
  wire _43928 = _43920 ^ _43927;
  wire _43929 = _1509 ^ _9572;
  wire _43930 = _7824 ^ _3058;
  wire _43931 = _43929 ^ _43930;
  wire _43932 = _1513 ^ _7828;
  wire _43933 = _8428 ^ _43932;
  wire _43934 = _43931 ^ _43933;
  wire _43935 = _3840 ^ _6600;
  wire _43936 = _5293 ^ _3846;
  wire _43937 = _43935 ^ _43936;
  wire _43938 = _16954 ^ _23163;
  wire _43939 = _10118 ^ _10120;
  wire _43940 = _43938 ^ _43939;
  wire _43941 = _43937 ^ _43940;
  wire _43942 = _43934 ^ _43941;
  wire _43943 = _43928 ^ _43942;
  wire _43944 = _43913 ^ _43943;
  wire _43945 = _24058 ^ _15498;
  wire _43946 = uncoded_block[1435] ^ uncoded_block[1440];
  wire _43947 = _43946 ^ _1541;
  wire _43948 = _43945 ^ _43947;
  wire _43949 = _2325 ^ _6622;
  wire _43950 = _43949 ^ _35422;
  wire _43951 = _43948 ^ _43950;
  wire _43952 = _9602 ^ _35423;
  wire _43953 = _13963 ^ _1562;
  wire _43954 = _43952 ^ _43953;
  wire _43955 = uncoded_block[1494] ^ uncoded_block[1497];
  wire _43956 = _43955 ^ _3109;
  wire _43957 = _36647 ^ _43956;
  wire _43958 = _43954 ^ _43957;
  wire _43959 = _43951 ^ _43958;
  wire _43960 = _11264 ^ _5333;
  wire _43961 = _9620 ^ _9055;
  wire _43962 = _43960 ^ _43961;
  wire _43963 = _754 ^ _3900;
  wire _43964 = _22266 ^ _12914;
  wire _43965 = _43963 ^ _43964;
  wire _43966 = _43962 ^ _43965;
  wire _43967 = uncoded_block[1542] ^ uncoded_block[1545];
  wire _43968 = _15009 ^ _43967;
  wire _43969 = _13471 ^ _9070;
  wire _43970 = _43968 ^ _43969;
  wire _43971 = _37871 ^ _7285;
  wire _43972 = _40236 ^ _43971;
  wire _43973 = _43970 ^ _43972;
  wire _43974 = _43966 ^ _43973;
  wire _43975 = _43959 ^ _43974;
  wire _43976 = _42545 ^ _24105;
  wire _43977 = _3927 ^ _3146;
  wire _43978 = _15541 ^ _1621;
  wire _43979 = _43977 ^ _43978;
  wire _43980 = _43976 ^ _43979;
  wire _43981 = uncoded_block[1601] ^ uncoded_block[1605];
  wire _43982 = _43981 ^ _3154;
  wire _43983 = _43982 ^ _10182;
  wire _43984 = _7911 ^ _6684;
  wire _43985 = _5386 ^ _1636;
  wire _43986 = _43984 ^ _43985;
  wire _43987 = _43983 ^ _43986;
  wire _43988 = _43980 ^ _43987;
  wire _43989 = _1646 ^ _816;
  wire _43990 = _38670 ^ _43989;
  wire _43991 = _1649 ^ _17529;
  wire _43992 = _7925 ^ _10196;
  wire _43993 = _43991 ^ _43992;
  wire _43994 = _43990 ^ _43993;
  wire _43995 = uncoded_block[1666] ^ uncoded_block[1672];
  wire _43996 = _3179 ^ _43995;
  wire _43997 = _43996 ^ _29158;
  wire _43998 = _7933 ^ _9675;
  wire _43999 = _3972 ^ _11327;
  wire _44000 = _43998 ^ _43999;
  wire _44001 = _43997 ^ _44000;
  wire _44002 = _43994 ^ _44001;
  wire _44003 = _43988 ^ _44002;
  wire _44004 = _43975 ^ _44003;
  wire _44005 = _43944 ^ _44004;
  wire _44006 = _16551 ^ _851;
  wire _44007 = _9126 ^ _12976;
  wire _44008 = _44006 ^ _44007;
  wire _44009 = _44008 ^ uncoded_block[1722];
  wire _44010 = _44005 ^ _44009;
  wire _44011 = _43883 ^ _44010;
  wire _44012 = _2 ^ _21409;
  wire _44013 = _43260 ^ _22790;
  wire _44014 = _40284 ^ _44013;
  wire _44015 = _44012 ^ _44014;
  wire _44016 = _21412 ^ _3225;
  wire _44017 = _44016 ^ _24610;
  wire _44018 = _4008 ^ _7359;
  wire _44019 = _44018 ^ _39105;
  wire _44020 = _44017 ^ _44019;
  wire _44021 = _44015 ^ _44020;
  wire _44022 = _7365 ^ _11357;
  wire _44023 = _44022 ^ _13557;
  wire _44024 = _6749 ^ _6754;
  wire _44025 = _6755 ^ _8566;
  wire _44026 = _44024 ^ _44025;
  wire _44027 = _44023 ^ _44026;
  wire _44028 = _4026 ^ _4745;
  wire _44029 = _19025 ^ _911;
  wire _44030 = _44028 ^ _44029;
  wire _44031 = _37537 ^ _13014;
  wire _44032 = _44031 ^ _23714;
  wire _44033 = _44030 ^ _44032;
  wire _44034 = _44027 ^ _44033;
  wire _44035 = _44021 ^ _44034;
  wire _44036 = _38721 ^ _38723;
  wire _44037 = _8581 ^ _6776;
  wire _44038 = _44036 ^ _44037;
  wire _44039 = _6138 ^ _6780;
  wire _44040 = _44039 ^ _1746;
  wire _44041 = _44038 ^ _44040;
  wire _44042 = _4049 ^ _29208;
  wire _44043 = _7398 ^ _44042;
  wire _44044 = _6788 ^ _938;
  wire _44045 = _3278 ^ _41855;
  wire _44046 = _44044 ^ _44045;
  wire _44047 = _44043 ^ _44046;
  wire _44048 = _44041 ^ _44047;
  wire _44049 = _2525 ^ _29628;
  wire _44050 = _44049 ^ _11401;
  wire _44051 = _6805 ^ _12479;
  wire _44052 = _28043 ^ _3292;
  wire _44053 = _44051 ^ _44052;
  wire _44054 = _44050 ^ _44053;
  wire _44055 = _960 ^ _102;
  wire _44056 = uncoded_block[223] ^ uncoded_block[227];
  wire _44057 = _44056 ^ _4791;
  wire _44058 = _44055 ^ _44057;
  wire _44059 = _22380 ^ _968;
  wire _44060 = _7423 ^ _7425;
  wire _44061 = _44059 ^ _44060;
  wire _44062 = _44058 ^ _44061;
  wire _44063 = _44054 ^ _44062;
  wire _44064 = _44048 ^ _44063;
  wire _44065 = _44035 ^ _44064;
  wire _44066 = _13053 ^ _14117;
  wire _44067 = _26433 ^ _44066;
  wire _44068 = _1786 ^ _7438;
  wire _44069 = _44068 ^ _6189;
  wire _44070 = _44067 ^ _44069;
  wire _44071 = uncoded_block[269] ^ uncoded_block[275];
  wire _44072 = _7440 ^ _44071;
  wire _44073 = _44072 ^ _21011;
  wire _44074 = _4105 ^ _11429;
  wire _44075 = _8633 ^ _13615;
  wire _44076 = _44074 ^ _44075;
  wire _44077 = _44073 ^ _44076;
  wire _44078 = _44070 ^ _44077;
  wire _44079 = _28067 ^ _145;
  wire _44080 = _35934 ^ _44079;
  wire _44081 = _1818 ^ _152;
  wire _44082 = _12518 ^ _44081;
  wire _44083 = _44080 ^ _44082;
  wire _44084 = _11444 ^ _9240;
  wire _44085 = _5536 ^ _1825;
  wire _44086 = _44084 ^ _44085;
  wire _44087 = _11987 ^ _7465;
  wire _44088 = _5541 ^ _15179;
  wire _44089 = _44087 ^ _44088;
  wire _44090 = _44086 ^ _44089;
  wire _44091 = _44083 ^ _44090;
  wire _44092 = _44078 ^ _44091;
  wire _44093 = _2602 ^ _3365;
  wire _44094 = _26032 ^ _17165;
  wire _44095 = _44093 ^ _44094;
  wire _44096 = _13094 ^ _10899;
  wire _44097 = _1841 ^ _19599;
  wire _44098 = _44096 ^ _44097;
  wire _44099 = _44095 ^ _44098;
  wire _44100 = _18633 ^ _42286;
  wire _44101 = _26042 ^ _17668;
  wire _44102 = _44100 ^ _44101;
  wire _44103 = _1055 ^ _4872;
  wire _44104 = _24244 ^ _44103;
  wire _44105 = _44102 ^ _44104;
  wire _44106 = _44099 ^ _44105;
  wire _44107 = _6889 ^ _6254;
  wire _44108 = _7497 ^ _5577;
  wire _44109 = _44107 ^ _44108;
  wire _44110 = _5578 ^ _24716;
  wire _44111 = uncoded_block[451] ^ uncoded_block[462];
  wire _44112 = _3411 ^ _44111;
  wire _44113 = _44110 ^ _44112;
  wire _44114 = _44109 ^ _44113;
  wire _44115 = _34776 ^ _9284;
  wire _44116 = _24723 ^ _8110;
  wire _44117 = _21982 ^ _44116;
  wire _44118 = _44115 ^ _44117;
  wire _44119 = _44114 ^ _44118;
  wire _44120 = _44106 ^ _44119;
  wire _44121 = _44092 ^ _44120;
  wire _44122 = _44065 ^ _44121;
  wire _44123 = _35592 ^ _8698;
  wire _44124 = _16697 ^ _44123;
  wire _44125 = _37227 ^ _19137;
  wire _44126 = _44124 ^ _44125;
  wire _44127 = _4918 ^ _20099;
  wire _44128 = _14709 ^ _44127;
  wire _44129 = _4925 ^ _6932;
  wire _44130 = _24279 ^ _6298;
  wire _44131 = _44129 ^ _44130;
  wire _44132 = _44128 ^ _44131;
  wire _44133 = _44126 ^ _44132;
  wire _44134 = uncoded_block[546] ^ uncoded_block[554];
  wire _44135 = _44134 ^ _12051;
  wire _44136 = _44135 ^ _9321;
  wire _44137 = _3467 ^ _4941;
  wire _44138 = _1132 ^ _10400;
  wire _44139 = _44137 ^ _44138;
  wire _44140 = _44136 ^ _44139;
  wire _44141 = _4946 ^ _266;
  wire _44142 = _20116 ^ _20618;
  wire _44143 = _44141 ^ _44142;
  wire _44144 = _1939 ^ _2710;
  wire _44145 = _278 ^ _7563;
  wire _44146 = _44144 ^ _44145;
  wire _44147 = _44143 ^ _44146;
  wire _44148 = _44140 ^ _44147;
  wire _44149 = _44133 ^ _44148;
  wire _44150 = _6960 ^ _12618;
  wire _44151 = _36844 ^ _44150;
  wire _44152 = _12620 ^ _3501;
  wire _44153 = _4249 ^ _6336;
  wire _44154 = _44152 ^ _44153;
  wire _44155 = _44151 ^ _44154;
  wire _44156 = _36853 ^ _4261;
  wire _44157 = _28530 ^ _44156;
  wire _44158 = _4262 ^ _9886;
  wire _44159 = uncoded_block[672] ^ uncoded_block[677];
  wire _44160 = uncoded_block[678] ^ uncoded_block[684];
  wire _44161 = _44159 ^ _44160;
  wire _44162 = _44158 ^ _44161;
  wire _44163 = _44157 ^ _44162;
  wire _44164 = _44155 ^ _44163;
  wire _44165 = _15281 ^ _4271;
  wire _44166 = _44165 ^ _20142;
  wire _44167 = _33204 ^ _2762;
  wire _44168 = _6993 ^ _44167;
  wire _44169 = _44166 ^ _44168;
  wire _44170 = _1194 ^ _5002;
  wire _44171 = uncoded_block[721] ^ uncoded_block[724];
  wire _44172 = _6367 ^ _44171;
  wire _44173 = _44170 ^ _44172;
  wire _44174 = _344 ^ _7603;
  wire _44175 = _44174 ^ _23426;
  wire _44176 = _44173 ^ _44175;
  wire _44177 = _44169 ^ _44176;
  wire _44178 = _44164 ^ _44177;
  wire _44179 = _44149 ^ _44178;
  wire _44180 = _352 ^ _11576;
  wire _44181 = _5012 ^ _2002;
  wire _44182 = _44180 ^ _44181;
  wire _44183 = _5019 ^ _5709;
  wire _44184 = _5711 ^ _34862;
  wire _44185 = _44183 ^ _44184;
  wire _44186 = _44182 ^ _44185;
  wire _44187 = _12675 ^ _1233;
  wire _44188 = _18747 ^ _44187;
  wire _44189 = _383 ^ _26589;
  wire _44190 = _5727 ^ _8228;
  wire _44191 = _44189 ^ _44190;
  wire _44192 = _44188 ^ _44191;
  wire _44193 = _44186 ^ _44192;
  wire _44194 = _5046 ^ _3584;
  wire _44195 = _31114 ^ _44194;
  wire _44196 = _44195 ^ _3592;
  wire _44197 = _16293 ^ _10495;
  wire _44198 = _44197 ^ _36895;
  wire _44199 = uncoded_block[858] ^ uncoded_block[863];
  wire _44200 = _44199 ^ _5071;
  wire _44201 = _13243 ^ _44200;
  wire _44202 = _44198 ^ _44201;
  wire _44203 = _44196 ^ _44202;
  wire _44204 = _44193 ^ _44203;
  wire _44205 = _5753 ^ _8820;
  wire _44206 = _4348 ^ _44205;
  wire _44207 = _2058 ^ _1273;
  wire _44208 = uncoded_block[894] ^ uncoded_block[901];
  wire _44209 = _12704 ^ _44208;
  wire _44210 = _44207 ^ _44209;
  wire _44211 = _44206 ^ _44210;
  wire _44212 = _1280 ^ _5761;
  wire _44213 = _2071 ^ _7665;
  wire _44214 = _44212 ^ _44213;
  wire _44215 = _17818 ^ _438;
  wire _44216 = _15840 ^ _8260;
  wire _44217 = _44215 ^ _44216;
  wire _44218 = _44214 ^ _44217;
  wire _44219 = _44211 ^ _44218;
  wire _44220 = _5096 ^ _25736;
  wire _44221 = _26189 ^ _23926;
  wire _44222 = _44220 ^ _44221;
  wire _44223 = _5779 ^ _9437;
  wire _44224 = _44223 ^ _12729;
  wire _44225 = _44222 ^ _44224;
  wire _44226 = _17334 ^ _1316;
  wire _44227 = _5114 ^ _11094;
  wire _44228 = _3659 ^ _12186;
  wire _44229 = _44227 ^ _44228;
  wire _44230 = _44226 ^ _44229;
  wire _44231 = _44225 ^ _44230;
  wire _44232 = _44219 ^ _44231;
  wire _44233 = _44204 ^ _44232;
  wire _44234 = _44179 ^ _44233;
  wire _44235 = _44122 ^ _44234;
  wire _44236 = _15369 ^ _2882;
  wire _44237 = _22575 ^ _13277;
  wire _44238 = _44236 ^ _44237;
  wire _44239 = _35704 ^ _20730;
  wire _44240 = uncoded_block[1011] ^ uncoded_block[1020];
  wire _44241 = _1327 ^ _44240;
  wire _44242 = _44239 ^ _44241;
  wire _44243 = _44238 ^ _44242;
  wire _44244 = _495 ^ _1339;
  wire _44245 = _21208 ^ _44244;
  wire _44246 = _499 ^ _501;
  wire _44247 = _44246 ^ _16351;
  wire _44248 = _44245 ^ _44247;
  wire _44249 = _44243 ^ _44248;
  wire _44250 = _512 ^ _2133;
  wire _44251 = _10011 ^ _4430;
  wire _44252 = _44250 ^ _44251;
  wire _44253 = _12764 ^ _2921;
  wire _44254 = _44253 ^ _11123;
  wire _44255 = _44252 ^ _44254;
  wire _44256 = _3692 ^ _15883;
  wire _44257 = _5839 ^ _10021;
  wire _44258 = _44256 ^ _44257;
  wire _44259 = uncoded_block[1097] ^ uncoded_block[1102];
  wire _44260 = _44259 ^ _39734;
  wire _44261 = _33727 ^ _44260;
  wire _44262 = _44258 ^ _44261;
  wire _44263 = _44255 ^ _44262;
  wire _44264 = _44249 ^ _44263;
  wire _44265 = _8918 ^ _13323;
  wire _44266 = _7736 ^ _3718;
  wire _44267 = uncoded_block[1128] ^ uncoded_block[1133];
  wire _44268 = _4459 ^ _44267;
  wire _44269 = _44266 ^ _44268;
  wire _44270 = _44265 ^ _44269;
  wire _44271 = _5856 ^ _20266;
  wire _44272 = _36139 ^ _8932;
  wire _44273 = _44271 ^ _44272;
  wire _44274 = _27532 ^ _11711;
  wire _44275 = _2958 ^ _2964;
  wire _44276 = _44274 ^ _44275;
  wire _44277 = _44273 ^ _44276;
  wire _44278 = _44270 ^ _44277;
  wire _44279 = _36971 ^ _12250;
  wire _44280 = _16898 ^ _590;
  wire _44281 = _6520 ^ _2200;
  wire _44282 = _44280 ^ _44281;
  wire _44283 = _44279 ^ _44282;
  wire _44284 = _33330 ^ _14398;
  wire _44285 = _7758 ^ _7763;
  wire _44286 = _44284 ^ _44285;
  wire _44287 = _1425 ^ _2216;
  wire _44288 = _12259 ^ _14914;
  wire _44289 = _44287 ^ _44288;
  wire _44290 = _44286 ^ _44289;
  wire _44291 = _44283 ^ _44290;
  wire _44292 = _44278 ^ _44291;
  wire _44293 = _44264 ^ _44292;
  wire _44294 = _13355 ^ _4504;
  wire _44295 = _18400 ^ _1442;
  wire _44296 = _44294 ^ _44295;
  wire _44297 = _7774 ^ _4509;
  wire _44298 = _44297 ^ _13366;
  wire _44299 = _44296 ^ _44298;
  wire _44300 = uncoded_block[1253] ^ uncoded_block[1257];
  wire _44301 = _5901 ^ _44300;
  wire _44302 = _5234 ^ _7178;
  wire _44303 = _44301 ^ _44302;
  wire _44304 = _33763 ^ _21738;
  wire _44305 = _44303 ^ _44304;
  wire _44306 = _44299 ^ _44305;
  wire _44307 = _21280 ^ _3794;
  wire _44308 = _16924 ^ _13380;
  wire _44309 = _44307 ^ _44308;
  wire _44310 = _9545 ^ _3801;
  wire _44311 = _17927 ^ _1472;
  wire _44312 = _44310 ^ _44311;
  wire _44313 = _44309 ^ _44312;
  wire _44314 = _8407 ^ _4540;
  wire _44315 = _23570 ^ _44314;
  wire _44316 = uncoded_block[1326] ^ uncoded_block[1330];
  wire _44317 = _44316 ^ _5931;
  wire _44318 = _32098 ^ _44317;
  wire _44319 = _44315 ^ _44318;
  wire _44320 = _44313 ^ _44319;
  wire _44321 = _44306 ^ _44320;
  wire _44322 = _10092 ^ _17938;
  wire _44323 = _35781 ^ _44322;
  wire _44324 = _11771 ^ _3041;
  wire _44325 = _44324 ^ _22222;
  wire _44326 = _44323 ^ _44325;
  wire _44327 = _5273 ^ _25393;
  wire _44328 = _44327 ^ _33367;
  wire _44329 = _11227 ^ _18443;
  wire _44330 = _44328 ^ _44329;
  wire _44331 = _44326 ^ _44330;
  wire _44332 = uncoded_block[1388] ^ uncoded_block[1391];
  wire _44333 = _44332 ^ _1516;
  wire _44334 = _25851 ^ _44333;
  wire _44335 = _16458 ^ _3847;
  wire _44336 = _5957 ^ _5961;
  wire _44337 = _44335 ^ _44336;
  wire _44338 = _44334 ^ _44337;
  wire _44339 = _5962 ^ _2306;
  wire _44340 = _17960 ^ _2308;
  wire _44341 = _44339 ^ _44340;
  wire _44342 = _24521 ^ _2319;
  wire _44343 = _44342 ^ _4592;
  wire _44344 = _44341 ^ _44343;
  wire _44345 = _44338 ^ _44344;
  wire _44346 = _44331 ^ _44345;
  wire _44347 = _44321 ^ _44346;
  wire _44348 = _44293 ^ _44347;
  wire _44349 = _35806 ^ _7854;
  wire _44350 = _20361 ^ _3094;
  wire _44351 = _1550 ^ _20367;
  wire _44352 = _44350 ^ _44351;
  wire _44353 = _44349 ^ _44352;
  wire _44354 = _9610 ^ _15994;
  wire _44355 = _2349 ^ _9044;
  wire _44356 = _44354 ^ _44355;
  wire _44357 = uncoded_block[1497] ^ uncoded_block[1504];
  wire _44358 = _3890 ^ _44357;
  wire _44359 = _19421 ^ _5336;
  wire _44360 = _44358 ^ _44359;
  wire _44361 = _44356 ^ _44360;
  wire _44362 = _44353 ^ _44361;
  wire _44363 = _6643 ^ _1579;
  wire _44364 = uncoded_block[1527] ^ uncoded_block[1531];
  wire _44365 = _8473 ^ _44364;
  wire _44366 = _44363 ^ _44365;
  wire _44367 = _36235 ^ _34228;
  wire _44368 = _44366 ^ _44367;
  wire _44369 = _3128 ^ _30858;
  wire _44370 = _14496 ^ _5358;
  wire _44371 = _44369 ^ _44370;
  wire _44372 = uncoded_block[1560] ^ uncoded_block[1564];
  wire _44373 = _44372 ^ _11284;
  wire _44374 = _44373 ^ _30444;
  wire _44375 = _44371 ^ _44374;
  wire _44376 = _44368 ^ _44375;
  wire _44377 = _44362 ^ _44376;
  wire _44378 = _4648 ^ _1609;
  wire _44379 = _44378 ^ _42552;
  wire _44380 = _6673 ^ _792;
  wire _44381 = _3934 ^ _3936;
  wire _44382 = _44380 ^ _44381;
  wire _44383 = _44379 ^ _44382;
  wire _44384 = _1625 ^ _42166;
  wire _44385 = _44384 ^ _21374;
  wire _44386 = _18020 ^ _18023;
  wire _44387 = uncoded_block[1627] ^ uncoded_block[1632];
  wire _44388 = _10185 ^ _44387;
  wire _44389 = _44386 ^ _44388;
  wire _44390 = _44385 ^ _44389;
  wire _44391 = _44383 ^ _44390;
  wire _44392 = _7914 ^ _7306;
  wire _44393 = uncoded_block[1640] ^ uncoded_block[1646];
  wire _44394 = uncoded_block[1655] ^ uncoded_block[1659];
  wire _44395 = _44393 ^ _44394;
  wire _44396 = _44392 ^ _44395;
  wire _44397 = _41801 ^ _4687;
  wire _44398 = _44397 ^ _7324;
  wire _44399 = _44396 ^ _44398;
  wire _44400 = _5401 ^ _25480;
  wire _44401 = _44400 ^ _30021;
  wire _44402 = _20436 ^ _1672;
  wire _44403 = _43999 ^ _44402;
  wire _44404 = _44401 ^ _44403;
  wire _44405 = _44399 ^ _44404;
  wire _44406 = _44391 ^ _44405;
  wire _44407 = _44377 ^ _44406;
  wire _44408 = uncoded_block[1708] ^ uncoded_block[1711];
  wire _44409 = _44408 ^ _11333;
  wire _44410 = _44409 ^ _38689;
  wire _44411 = _44410 ^ uncoded_block[1722];
  wire _44412 = _44407 ^ _44411;
  wire _44413 = _44348 ^ _44412;
  wire _44414 = _44235 ^ _44413;
  wire _44415 = _10226 ^ _20453;
  wire _44416 = _7959 ^ _1693;
  wire _44417 = _44415 ^ _44416;
  wire _44418 = _41028 ^ _44417;
  wire _44419 = _18 ^ _20941;
  wire _44420 = _41033 ^ _44419;
  wire _44421 = uncoded_block[47] ^ uncoded_block[53];
  wire _44422 = _12425 ^ _44421;
  wire _44423 = _16572 ^ _13553;
  wire _44424 = _44422 ^ _44423;
  wire _44425 = _44420 ^ _44424;
  wire _44426 = _44418 ^ _44425;
  wire _44427 = _10806 ^ _34;
  wire _44428 = _6745 ^ _21881;
  wire _44429 = _44427 ^ _44428;
  wire _44430 = uncoded_block[87] ^ uncoded_block[94];
  wire _44431 = _11364 ^ _44430;
  wire _44432 = _6751 ^ _44431;
  wire _44433 = _44429 ^ _44432;
  wire _44434 = _47 ^ _15097;
  wire _44435 = _15101 ^ _33056;
  wire _44436 = _44434 ^ _44435;
  wire _44437 = _13016 ^ _917;
  wire _44438 = _4042 ^ _8581;
  wire _44439 = _44437 ^ _44438;
  wire _44440 = _44436 ^ _44439;
  wire _44441 = _44433 ^ _44440;
  wire _44442 = _44426 ^ _44441;
  wire _44443 = _64 ^ _9730;
  wire _44444 = _67 ^ _1744;
  wire _44445 = _44443 ^ _44444;
  wire _44446 = _5469 ^ _23281;
  wire _44447 = _44446 ^ _4055;
  wire _44448 = _44445 ^ _44447;
  wire _44449 = _41061 ^ _940;
  wire _44450 = _33491 ^ _44449;
  wire _44451 = _4062 ^ _13588;
  wire _44452 = _20981 ^ _44451;
  wire _44453 = _44450 ^ _44452;
  wire _44454 = _44448 ^ _44453;
  wire _44455 = _25983 ^ _35908;
  wire _44456 = _33496 ^ _44455;
  wire _44457 = _14101 ^ _19549;
  wire _44458 = _44457 ^ _8607;
  wire _44459 = _44456 ^ _44458;
  wire _44460 = _25990 ^ _22380;
  wire _44461 = _6822 ^ _970;
  wire _44462 = _44460 ^ _44461;
  wire _44463 = _5503 ^ _4085;
  wire _44464 = _44463 ^ _37568;
  wire _44465 = _44462 ^ _44464;
  wire _44466 = _44459 ^ _44465;
  wire _44467 = _44454 ^ _44466;
  wire _44468 = _44442 ^ _44467;
  wire _44469 = _9761 ^ _20520;
  wire _44470 = _44469 ^ _26443;
  wire _44471 = _6192 ^ _36768;
  wire _44472 = _44471 ^ _9773;
  wire _44473 = _44470 ^ _44472;
  wire _44474 = _2571 ^ _995;
  wire _44475 = _44474 ^ _41092;
  wire _44476 = _18142 ^ _27319;
  wire _44477 = _44475 ^ _44476;
  wire _44478 = _44473 ^ _44477;
  wire _44479 = _3346 ^ _2583;
  wire _44480 = _11444 ^ _26461;
  wire _44481 = _44479 ^ _44480;
  wire _44482 = uncoded_block[336] ^ uncoded_block[342];
  wire _44483 = _44482 ^ _4841;
  wire _44484 = _11454 ^ _20554;
  wire _44485 = _44483 ^ _44484;
  wire _44486 = _44481 ^ _44485;
  wire _44487 = _7470 ^ _17165;
  wire _44488 = _44487 ^ _35947;
  wire _44489 = _4857 ^ _3377;
  wire _44490 = _2613 ^ _12005;
  wire _44491 = _44489 ^ _44490;
  wire _44492 = _44488 ^ _44491;
  wire _44493 = _44486 ^ _44492;
  wire _44494 = _44478 ^ _44493;
  wire _44495 = _5559 ^ _5561;
  wire _44496 = _41114 ^ _44495;
  wire _44497 = _3391 ^ _24243;
  wire _44498 = _13110 ^ _13112;
  wire _44499 = _44497 ^ _44498;
  wire _44500 = _44496 ^ _44499;
  wire _44501 = uncoded_block[423] ^ uncoded_block[431];
  wire _44502 = _14160 ^ _44501;
  wire _44503 = _10352 ^ _25601;
  wire _44504 = _44502 ^ _44503;
  wire _44505 = _206 ^ _27756;
  wire _44506 = _14173 ^ _5586;
  wire _44507 = _44505 ^ _44506;
  wire _44508 = _44504 ^ _44507;
  wire _44509 = _44500 ^ _44508;
  wire _44510 = _4185 ^ _23357;
  wire _44511 = _3418 ^ _13132;
  wire _44512 = _44510 ^ _44511;
  wire _44513 = _7516 ^ _5604;
  wire _44514 = _1087 ^ _44513;
  wire _44515 = _44512 ^ _44514;
  wire _44516 = _27369 ^ _9298;
  wire _44517 = _14185 ^ _44516;
  wire _44518 = _19638 ^ _1107;
  wire _44519 = _1108 ^ _7534;
  wire _44520 = _44518 ^ _44519;
  wire _44521 = _44517 ^ _44520;
  wire _44522 = _44515 ^ _44521;
  wire _44523 = _44509 ^ _44522;
  wire _44524 = _44494 ^ _44523;
  wire _44525 = _44468 ^ _44524;
  wire _44526 = _2683 ^ _6293;
  wire _44527 = _44526 ^ _1910;
  wire _44528 = _4933 ^ _1122;
  wire _44529 = _44528 ^ _3462;
  wire _44530 = _44527 ^ _44529;
  wire _44531 = _3464 ^ _8727;
  wire _44532 = _44531 ^ _33597;
  wire _44533 = _3474 ^ _9325;
  wire _44534 = _266 ^ _270;
  wire _44535 = _44533 ^ _44534;
  wire _44536 = _44532 ^ _44535;
  wire _44537 = _44530 ^ _44536;
  wire _44538 = _33602 ^ _34809;
  wire _44539 = _41162 ^ _5653;
  wire _44540 = _43383 ^ _44539;
  wire _44541 = _44538 ^ _44540;
  wire _44542 = _4243 ^ _16738;
  wire _44543 = _4964 ^ _17238;
  wire _44544 = _44542 ^ _44543;
  wire _44545 = _14745 ^ _6330;
  wire _44546 = _44545 ^ _25203;
  wire _44547 = _44544 ^ _44546;
  wire _44548 = _44541 ^ _44547;
  wire _44549 = _44537 ^ _44548;
  wire _44550 = uncoded_block[641] ^ uncoded_block[645];
  wire _44551 = _4255 ^ _44550;
  wire _44552 = _6338 ^ _34028;
  wire _44553 = _44551 ^ _44552;
  wire _44554 = _14755 ^ _9352;
  wire _44555 = _44554 ^ _36024;
  wire _44556 = _44553 ^ _44555;
  wire _44557 = _6349 ^ _6352;
  wire _44558 = _26993 ^ _44557;
  wire _44559 = uncoded_block[686] ^ uncoded_block[692];
  wire _44560 = _5678 ^ _44559;
  wire _44561 = _44560 ^ _19685;
  wire _44562 = _44558 ^ _44561;
  wire _44563 = _44556 ^ _44562;
  wire _44564 = _4989 ^ _10447;
  wire _44565 = _4995 ^ _10452;
  wire _44566 = _44564 ^ _44565;
  wire _44567 = _1988 ^ _13749;
  wire _44568 = _35645 ^ _44567;
  wire _44569 = _44566 ^ _44568;
  wire _44570 = _25224 ^ _44180;
  wire _44571 = _5013 ^ _1210;
  wire _44572 = _21605 ^ _7015;
  wire _44573 = _44571 ^ _44572;
  wire _44574 = _44570 ^ _44573;
  wire _44575 = _44569 ^ _44574;
  wire _44576 = _44563 ^ _44575;
  wire _44577 = _44549 ^ _44576;
  wire _44578 = _4301 ^ _12113;
  wire _44579 = _36465 ^ _44578;
  wire _44580 = _9382 ^ _17284;
  wire _44581 = _14790 ^ _44580;
  wire _44582 = _44579 ^ _44581;
  wire _44583 = _1232 ^ _6391;
  wire _44584 = _18279 ^ _44583;
  wire _44585 = _44584 ^ _41216;
  wire _44586 = _44582 ^ _44585;
  wire _44587 = _393 ^ _14290;
  wire _44588 = _37697 ^ _44587;
  wire _44589 = uncoded_block[824] ^ uncoded_block[833];
  wire _44590 = _44589 ^ _22532;
  wire _44591 = _10495 ^ _1257;
  wire _44592 = _44590 ^ _44591;
  wire _44593 = _44588 ^ _44592;
  wire _44594 = _5741 ^ _15330;
  wire _44595 = _5066 ^ _13244;
  wire _44596 = _44594 ^ _44595;
  wire _44597 = _6415 ^ _15826;
  wire _44598 = _32811 ^ _44597;
  wire _44599 = _44596 ^ _44598;
  wire _44600 = _44593 ^ _44599;
  wire _44601 = _44586 ^ _44600;
  wire _44602 = _2835 ^ _423;
  wire _44603 = uncoded_block[890] ^ uncoded_block[896];
  wire _44604 = _5082 ^ _44603;
  wire _44605 = _44602 ^ _44604;
  wire _44606 = _1278 ^ _8254;
  wire _44607 = _3623 ^ _432;
  wire _44608 = _44606 ^ _44607;
  wire _44609 = _44605 ^ _44608;
  wire _44610 = uncoded_block[913] ^ uncoded_block[917];
  wire _44611 = _12708 ^ _44610;
  wire _44612 = _41238 ^ _2076;
  wire _44613 = _44611 ^ _44612;
  wire _44614 = _11076 ^ _455;
  wire _44615 = _8263 ^ _44614;
  wire _44616 = _44613 ^ _44615;
  wire _44617 = _44609 ^ _44616;
  wire _44618 = _456 ^ _460;
  wire _44619 = _44618 ^ _27479;
  wire _44620 = uncoded_block[971] ^ uncoded_block[980];
  wire _44621 = _2093 ^ _44620;
  wire _44622 = _5792 ^ _8856;
  wire _44623 = _44621 ^ _44622;
  wire _44624 = _44619 ^ _44623;
  wire _44625 = _2882 ^ _479;
  wire _44626 = _44625 ^ _42415;
  wire _44627 = _25757 ^ _9994;
  wire _44628 = _44626 ^ _44627;
  wire _44629 = _44624 ^ _44628;
  wire _44630 = _44617 ^ _44629;
  wire _44631 = _44601 ^ _44630;
  wire _44632 = _44577 ^ _44631;
  wire _44633 = _44525 ^ _44632;
  wire _44634 = _28989 ^ _19766;
  wire _44635 = uncoded_block[1026] ^ uncoded_block[1030];
  wire _44636 = _44635 ^ _2907;
  wire _44637 = _44634 ^ _44636;
  wire _44638 = _502 ^ _43101;
  wire _44639 = _44638 ^ _24418;
  wire _44640 = _44637 ^ _44639;
  wire _44641 = _4430 ^ _12764;
  wire _44642 = _521 ^ _2917;
  wire _44643 = _44641 ^ _44642;
  wire _44644 = _8889 ^ _11122;
  wire _44645 = _15396 ^ _2146;
  wire _44646 = _44644 ^ _44645;
  wire _44647 = _44643 ^ _44646;
  wire _44648 = _44640 ^ _44647;
  wire _44649 = _2147 ^ _530;
  wire _44650 = _20753 ^ _3696;
  wire _44651 = _44649 ^ _44650;
  wire _44652 = _30740 ^ _33305;
  wire _44653 = _13316 ^ _549;
  wire _44654 = _44652 ^ _44653;
  wire _44655 = _44651 ^ _44654;
  wire _44656 = _2938 ^ _7736;
  wire _44657 = _4452 ^ _44656;
  wire _44658 = uncoded_block[1122] ^ uncoded_block[1126];
  wire _44659 = _44658 ^ _23523;
  wire _44660 = _44659 ^ _22621;
  wire _44661 = _44657 ^ _44660;
  wire _44662 = _44655 ^ _44661;
  wire _44663 = _44648 ^ _44662;
  wire _44664 = uncoded_block[1144] ^ uncoded_block[1153];
  wire _44665 = _568 ^ _44664;
  wire _44666 = _44665 ^ _24901;
  wire _44667 = _27537 ^ _27902;
  wire _44668 = _44667 ^ _591;
  wire _44669 = _44666 ^ _44668;
  wire _44670 = uncoded_block[1184] ^ uncoded_block[1188];
  wire _44671 = _44670 ^ _5203;
  wire _44672 = _14398 ^ _23999;
  wire _44673 = _44671 ^ _44672;
  wire _44674 = uncoded_block[1205] ^ uncoded_block[1209];
  wire _44675 = _2207 ^ _44674;
  wire _44676 = _1427 ^ _5213;
  wire _44677 = _44675 ^ _44676;
  wire _44678 = _44673 ^ _44677;
  wire _44679 = _44669 ^ _44678;
  wire _44680 = _3769 ^ _3771;
  wire _44681 = _27555 ^ _44680;
  wire _44682 = _15442 ^ _25815;
  wire _44683 = _44681 ^ _44682;
  wire _44684 = _621 ^ _8388;
  wire _44685 = _3001 ^ _5234;
  wire _44686 = _44684 ^ _44685;
  wire _44687 = _26712 ^ _6550;
  wire _44688 = _3008 ^ _11746;
  wire _44689 = _44687 ^ _44688;
  wire _44690 = _44686 ^ _44689;
  wire _44691 = _44683 ^ _44690;
  wire _44692 = _44679 ^ _44691;
  wire _44693 = _44663 ^ _44692;
  wire _44694 = _16419 ^ _3793;
  wire _44695 = _44694 ^ _34569;
  wire _44696 = _3798 ^ _2252;
  wire _44697 = _44696 ^ _41327;
  wire _44698 = _44695 ^ _44697;
  wire _44699 = _21748 ^ _4540;
  wire _44700 = _18878 ^ _44699;
  wire _44701 = _5254 ^ _13395;
  wire _44702 = _16435 ^ _21753;
  wire _44703 = _44701 ^ _44702;
  wire _44704 = _44700 ^ _44703;
  wire _44705 = _44698 ^ _44704;
  wire _44706 = _14949 ^ _39006;
  wire _44707 = _3042 ^ _10097;
  wire _44708 = _42114 ^ _44707;
  wire _44709 = _44706 ^ _44708;
  wire _44710 = _5273 ^ _23148;
  wire _44711 = _2284 ^ _41346;
  wire _44712 = _44710 ^ _44711;
  wire _44713 = _19861 ^ _16952;
  wire _44714 = _16452 ^ _44713;
  wire _44715 = _44712 ^ _44714;
  wire _44716 = _44709 ^ _44715;
  wire _44717 = _44705 ^ _44716;
  wire _44718 = _30393 ^ _31694;
  wire _44719 = _10113 ^ _17461;
  wire _44720 = _6607 ^ _9588;
  wire _44721 = _44719 ^ _44720;
  wire _44722 = _44718 ^ _44721;
  wire _44723 = _709 ^ _10684;
  wire _44724 = _1533 ^ _22242;
  wire _44725 = _44723 ^ _44724;
  wire _44726 = _24065 ^ _1541;
  wire _44727 = uncoded_block[1451] ^ uncoded_block[1456];
  wire _44728 = _16473 ^ _44727;
  wire _44729 = _44726 ^ _44728;
  wire _44730 = _44725 ^ _44729;
  wire _44731 = _44722 ^ _44730;
  wire _44732 = _3089 ^ _9602;
  wire _44733 = _44732 ^ _20857;
  wire _44734 = _2344 ^ _19887;
  wire _44735 = _44734 ^ _41370;
  wire _44736 = _44733 ^ _44735;
  wire _44737 = uncoded_block[1498] ^ uncoded_block[1507];
  wire _44738 = _44737 ^ _38638;
  wire _44739 = _44738 ^ _39049;
  wire _44740 = uncoded_block[1520] ^ uncoded_block[1525];
  wire _44741 = _7265 ^ _44740;
  wire _44742 = _13459 ^ _24549;
  wire _44743 = _44741 ^ _44742;
  wire _44744 = _44739 ^ _44743;
  wire _44745 = _44736 ^ _44744;
  wire _44746 = _44731 ^ _44745;
  wire _44747 = _44717 ^ _44746;
  wire _44748 = _44693 ^ _44747;
  wire _44749 = _6651 ^ _4634;
  wire _44750 = _44749 ^ _13473;
  wire _44751 = _769 ^ _1596;
  wire _44752 = uncoded_block[1563] ^ uncoded_block[1570];
  wire _44753 = _1597 ^ _44752;
  wire _44754 = _44751 ^ _44753;
  wire _44755 = _44750 ^ _44754;
  wire _44756 = _4647 ^ _15535;
  wire _44757 = uncoded_block[1586] ^ uncoded_block[1591];
  wire _44758 = _44757 ^ _21827;
  wire _44759 = _44756 ^ _44758;
  wire _44760 = _6040 ^ _4662;
  wire _44761 = _15037 ^ _44760;
  wire _44762 = _44759 ^ _44761;
  wire _44763 = _44755 ^ _44762;
  wire _44764 = _9095 ^ _31746;
  wire _44765 = _1634 ^ _44764;
  wire _44766 = _812 ^ _7306;
  wire _44767 = _41400 ^ _44766;
  wire _44768 = _44765 ^ _44767;
  wire _44769 = _27652 ^ _41405;
  wire _44770 = _820 ^ _10761;
  wire _44771 = _7927 ^ _12395;
  wire _44772 = _44770 ^ _44771;
  wire _44773 = _44769 ^ _44772;
  wire _44774 = _44768 ^ _44773;
  wire _44775 = _44763 ^ _44774;
  wire _44776 = _30014 ^ _5401;
  wire _44777 = _16541 ^ _39083;
  wire _44778 = _44776 ^ _44777;
  wire _44779 = _26365 ^ _1669;
  wire _44780 = _3973 ^ _21400;
  wire _44781 = _44779 ^ _44780;
  wire _44782 = _44778 ^ _44781;
  wire _44783 = _7337 ^ _30908;
  wire _44784 = _44783 ^ uncoded_block[1717];
  wire _44785 = _44782 ^ _44784;
  wire _44786 = _44775 ^ _44785;
  wire _44787 = _44748 ^ _44786;
  wire _44788 = _44633 ^ _44787;
  wire _44789 = _4710 ^ _3995;
  wire _44790 = uncoded_block[14] ^ uncoded_block[19];
  wire _44791 = _19001 ^ _44790;
  wire _44792 = _44789 ^ _44791;
  wire _44793 = _3220 ^ _25941;
  wire _44794 = _882 ^ _6736;
  wire _44795 = _44793 ^ _44794;
  wire _44796 = _44792 ^ _44795;
  wire _44797 = _12429 ^ _23256;
  wire _44798 = uncoded_block[61] ^ uncoded_block[67];
  wire _44799 = _44798 ^ _35;
  wire _44800 = _44797 ^ _44799;
  wire _44801 = _3241 ^ _1714;
  wire _44802 = _41 ^ _17578;
  wire _44803 = _44801 ^ _44802;
  wire _44804 = _44800 ^ _44803;
  wire _44805 = _44796 ^ _44804;
  wire _44806 = uncoded_block[93] ^ uncoded_block[98];
  wire _44807 = _14065 ^ _44806;
  wire _44808 = _44807 ^ _28442;
  wire _44809 = _1722 ^ _54;
  wire _44810 = _9721 ^ _13016;
  wire _44811 = _44809 ^ _44810;
  wire _44812 = _44808 ^ _44811;
  wire _44813 = _3262 ^ _9177;
  wire _44814 = _9729 ^ _5461;
  wire _44815 = _44813 ^ _44814;
  wire _44816 = _2511 ^ _1744;
  wire _44817 = uncoded_block[151] ^ uncoded_block[154];
  wire _44818 = uncoded_block[160] ^ uncoded_block[167];
  wire _44819 = _44817 ^ _44818;
  wire _44820 = _44816 ^ _44819;
  wire _44821 = _44815 ^ _44820;
  wire _44822 = _44812 ^ _44821;
  wire _44823 = _44805 ^ _44822;
  wire _44824 = uncoded_block[169] ^ uncoded_block[175];
  wire _44825 = _44824 ^ _941;
  wire _44826 = _2528 ^ _18111;
  wire _44827 = _44825 ^ _44826;
  wire _44828 = _18113 ^ _1763;
  wire _44829 = _44828 ^ _32247;
  wire _44830 = _44827 ^ _44829;
  wire _44831 = _953 ^ _4071;
  wire _44832 = _44831 ^ _21461;
  wire _44833 = _3299 ^ _16125;
  wire _44834 = _35533 ^ _44833;
  wire _44835 = _44832 ^ _44834;
  wire _44836 = _44830 ^ _44835;
  wire _44837 = uncoded_block[238] ^ uncoded_block[243];
  wire _44838 = _24660 ^ _44837;
  wire _44839 = _11952 ^ _7432;
  wire _44840 = _44838 ^ _44839;
  wire _44841 = _6182 ^ _1789;
  wire _44842 = uncoded_block[271] ^ uncoded_block[276];
  wire _44843 = _985 ^ _44842;
  wire _44844 = _44841 ^ _44843;
  wire _44845 = _44840 ^ _44844;
  wire _44846 = _10303 ^ _6194;
  wire _44847 = _11424 ^ _9226;
  wire _44848 = _44846 ^ _44847;
  wire _44849 = _15665 ^ _10312;
  wire _44850 = _14133 ^ _13074;
  wire _44851 = _44849 ^ _44850;
  wire _44852 = _44848 ^ _44851;
  wire _44853 = _44845 ^ _44852;
  wire _44854 = _44836 ^ _44853;
  wire _44855 = _44823 ^ _44854;
  wire _44856 = uncoded_block[319] ^ uncoded_block[324];
  wire _44857 = _1006 ^ _44856;
  wire _44858 = _152 ^ _5534;
  wire _44859 = _44857 ^ _44858;
  wire _44860 = _8063 ^ _3352;
  wire _44861 = _44860 ^ _8647;
  wire _44862 = _44859 ^ _44861;
  wire _44863 = _2596 ^ _2599;
  wire _44864 = _162 ^ _3361;
  wire _44865 = _44863 ^ _44864;
  wire _44866 = _3362 ^ _5548;
  wire _44867 = _14144 ^ _39961;
  wire _44868 = _44866 ^ _44867;
  wire _44869 = _44865 ^ _44868;
  wire _44870 = _44862 ^ _44869;
  wire _44871 = _23779 ^ _5554;
  wire _44872 = uncoded_block[404] ^ uncoded_block[410];
  wire _44873 = _17668 ^ _44872;
  wire _44874 = _44871 ^ _44873;
  wire _44875 = _2630 ^ _6249;
  wire _44876 = uncoded_block[423] ^ uncoded_block[428];
  wire _44877 = _44876 ^ _201;
  wire _44878 = _44875 ^ _44877;
  wire _44879 = _44874 ^ _44878;
  wire _44880 = _10356 ^ _19621;
  wire _44881 = _16681 ^ _44880;
  wire _44882 = uncoded_block[458] ^ uncoded_block[462];
  wire _44883 = _1870 ^ _44882;
  wire _44884 = _4185 ^ _1874;
  wire _44885 = _44883 ^ _44884;
  wire _44886 = _44881 ^ _44885;
  wire _44887 = _44879 ^ _44886;
  wire _44888 = _44870 ^ _44887;
  wire _44889 = _11494 ^ _19128;
  wire _44890 = _1880 ^ _44889;
  wire _44891 = _21528 ^ _7515;
  wire _44892 = _225 ^ _9292;
  wire _44893 = _44891 ^ _44892;
  wire _44894 = _44890 ^ _44893;
  wire _44895 = _229 ^ _10375;
  wire _44896 = _27369 ^ _3440;
  wire _44897 = _44895 ^ _44896;
  wire _44898 = _3444 ^ _1898;
  wire _44899 = _9301 ^ _16215;
  wire _44900 = _44898 ^ _44899;
  wire _44901 = _44897 ^ _44900;
  wire _44902 = _44894 ^ _44901;
  wire _44903 = uncoded_block[535] ^ uncoded_block[540];
  wire _44904 = _44903 ^ _8132;
  wire _44905 = _7541 ^ _6301;
  wire _44906 = _44904 ^ _44905;
  wire _44907 = uncoded_block[562] ^ uncoded_block[570];
  wire _44908 = _44907 ^ _11526;
  wire _44909 = _34407 ^ _44908;
  wire _44910 = _44906 ^ _44909;
  wire _44911 = _8733 ^ _9864;
  wire _44912 = _2700 ^ _7556;
  wire _44913 = _44911 ^ _44912;
  wire _44914 = _7558 ^ _6954;
  wire _44915 = _44914 ^ _44145;
  wire _44916 = _44913 ^ _44915;
  wire _44917 = _44910 ^ _44916;
  wire _44918 = _44902 ^ _44917;
  wire _44919 = _44888 ^ _44918;
  wire _44920 = _44855 ^ _44919;
  wire _44921 = _24299 ^ _3495;
  wire _44922 = _12618 ^ _18235;
  wire _44923 = _44921 ^ _44922;
  wire _44924 = uncoded_block[632] ^ uncoded_block[638];
  wire _44925 = _44924 ^ _8751;
  wire _44926 = _26112 ^ _28908;
  wire _44927 = _44925 ^ _44926;
  wire _44928 = _44923 ^ _44927;
  wire _44929 = uncoded_block[654] ^ uncoded_block[661];
  wire _44930 = _44929 ^ _22960;
  wire _44931 = _44930 ^ _313;
  wire _44932 = uncoded_block[674] ^ uncoded_block[693];
  wire _44933 = uncoded_block[695] ^ uncoded_block[698];
  wire _44934 = _44932 ^ _44933;
  wire _44935 = _3532 ^ _5685;
  wire _44936 = _44934 ^ _44935;
  wire _44937 = _44931 ^ _44936;
  wire _44938 = _44928 ^ _44937;
  wire _44939 = _337 ^ _4999;
  wire _44940 = _341 ^ _15292;
  wire _44941 = _44939 ^ _44940;
  wire _44942 = _26566 ^ _1995;
  wire _44943 = _7005 ^ _5010;
  wire _44944 = _44942 ^ _44943;
  wire _44945 = _44941 ^ _44944;
  wire _44946 = _4293 ^ _15795;
  wire _44947 = _1217 ^ _2011;
  wire _44948 = _44946 ^ _44947;
  wire _44949 = _3568 ^ _25694;
  wire _44950 = _36051 ^ _44949;
  wire _44951 = _44948 ^ _44950;
  wire _44952 = _44945 ^ _44951;
  wire _44953 = _44938 ^ _44952;
  wire _44954 = uncoded_block[797] ^ uncoded_block[804];
  wire _44955 = _44954 ^ _12127;
  wire _44956 = _33650 ^ _44955;
  wire _44957 = _14287 ^ _15318;
  wire _44958 = _5046 ^ _2028;
  wire _44959 = _44957 ^ _44958;
  wire _44960 = _44956 ^ _44959;
  wire _44961 = _5051 ^ _4330;
  wire _44962 = _44961 ^ _35272;
  wire _44963 = uncoded_block[846] ^ uncoded_block[852];
  wire _44964 = _44963 ^ _29368;
  wire _44965 = _11052 ^ _11618;
  wire _44966 = _44964 ^ _44965;
  wire _44967 = _44962 ^ _44966;
  wire _44968 = _44960 ^ _44967;
  wire _44969 = _9953 ^ _3608;
  wire _44970 = _4351 ^ _13797;
  wire _44971 = _44969 ^ _44970;
  wire _44972 = _16819 ^ _34081;
  wire _44973 = _2070 ^ _9424;
  wire _44974 = _44972 ^ _44973;
  wire _44975 = _44971 ^ _44974;
  wire _44976 = _23917 ^ _39692;
  wire _44977 = _44976 ^ _8263;
  wire _44978 = _7673 ^ _12723;
  wire _44979 = uncoded_block[947] ^ uncoded_block[954];
  wire _44980 = _44979 ^ _4384;
  wire _44981 = _44978 ^ _44980;
  wire _44982 = _44977 ^ _44981;
  wire _44983 = _44975 ^ _44982;
  wire _44984 = _44968 ^ _44983;
  wire _44985 = _44953 ^ _44984;
  wire _44986 = _9979 ^ _10531;
  wire _44987 = _468 ^ _4390;
  wire _44988 = _44986 ^ _44987;
  wire _44989 = _24853 ^ _16338;
  wire _44990 = _8854 ^ _44989;
  wire _44991 = _44988 ^ _44990;
  wire _44992 = _1323 ^ _15372;
  wire _44993 = _15373 ^ _17840;
  wire _44994 = _44992 ^ _44993;
  wire _44995 = uncoded_block[1015] ^ uncoded_block[1020];
  wire _44996 = _8296 ^ _44995;
  wire _44997 = _27494 ^ _13288;
  wire _44998 = _44996 ^ _44997;
  wire _44999 = _44994 ^ _44998;
  wire _45000 = _44991 ^ _44999;
  wire _45001 = uncoded_block[1031] ^ uncoded_block[1034];
  wire _45002 = _45001 ^ _1342;
  wire _45003 = _5810 ^ _19777;
  wire _45004 = _45002 ^ _45003;
  wire _45005 = uncoded_block[1047] ^ uncoded_block[1052];
  wire _45006 = _45005 ^ _1360;
  wire _45007 = uncoded_block[1068] ^ uncoded_block[1072];
  wire _45008 = _1363 ^ _45007;
  wire _45009 = _45006 ^ _45008;
  wire _45010 = _45004 ^ _45009;
  wire _45011 = _5831 ^ _17362;
  wire _45012 = _10575 ^ _22149;
  wire _45013 = _45011 ^ _45012;
  wire _45014 = _34942 ^ _18825;
  wire _45015 = _45013 ^ _45014;
  wire _45016 = _45010 ^ _45015;
  wire _45017 = _45000 ^ _45016;
  wire _45018 = _2164 ^ _26671;
  wire _45019 = uncoded_block[1127] ^ uncoded_block[1131];
  wire _45020 = _29427 ^ _45019;
  wire _45021 = _45018 ^ _45020;
  wire _45022 = uncoded_block[1138] ^ uncoded_block[1144];
  wire _45023 = _564 ^ _45022;
  wire _45024 = _26240 ^ _3728;
  wire _45025 = _45023 ^ _45024;
  wire _45026 = _45021 ^ _45025;
  wire _45027 = _22627 ^ _30756;
  wire _45028 = _584 ^ _27113;
  wire _45029 = _45027 ^ _45028;
  wire _45030 = _15428 ^ _11719;
  wire _45031 = _11721 ^ _44674;
  wire _45032 = _45030 ^ _45031;
  wire _45033 = _45029 ^ _45032;
  wire _45034 = _45026 ^ _45033;
  wire _45035 = _1428 ^ _14407;
  wire _45036 = uncoded_block[1222] ^ uncoded_block[1225];
  wire _45037 = uncoded_block[1227] ^ uncoded_block[1235];
  wire _45038 = _45036 ^ _45037;
  wire _45039 = _45035 ^ _45038;
  wire _45040 = _1443 ^ _17910;
  wire _45041 = _37796 ^ _6546;
  wire _45042 = _45040 ^ _45041;
  wire _45043 = _45039 ^ _45042;
  wire _45044 = _1455 ^ _30361;
  wire _45045 = _34567 ^ _9539;
  wire _45046 = _45044 ^ _45045;
  wire _45047 = _3793 ^ _28317;
  wire _45048 = uncoded_block[1303] ^ uncoded_block[1310];
  wire _45049 = _21741 ^ _45048;
  wire _45050 = _45047 ^ _45049;
  wire _45051 = _45046 ^ _45050;
  wire _45052 = _45043 ^ _45051;
  wire _45053 = _45034 ^ _45052;
  wire _45054 = _45017 ^ _45053;
  wire _45055 = _44985 ^ _45054;
  wire _45056 = _44920 ^ _45055;
  wire _45057 = uncoded_block[1315] ^ uncoded_block[1324];
  wire _45058 = _20314 ^ _45057;
  wire _45059 = _656 ^ _13922;
  wire _45060 = _45058 ^ _45059;
  wire _45061 = _8413 ^ _4553;
  wire _45062 = _45061 ^ _23143;
  wire _45063 = _45060 ^ _45062;
  wire _45064 = _11218 ^ _3042;
  wire _45065 = uncoded_block[1354] ^ uncoded_block[1357];
  wire _45066 = uncoded_block[1358] ^ uncoded_block[1364];
  wire _45067 = _45065 ^ _45066;
  wire _45068 = _45064 ^ _45067;
  wire _45069 = _10665 ^ _29934;
  wire _45070 = _7823 ^ _26743;
  wire _45071 = _45069 ^ _45070;
  wire _45072 = _45068 ^ _45071;
  wire _45073 = _45063 ^ _45072;
  wire _45074 = uncoded_block[1384] ^ uncoded_block[1390];
  wire _45075 = _3059 ^ _45074;
  wire _45076 = _45075 ^ _27164;
  wire _45077 = _3066 ^ _5293;
  wire _45078 = uncoded_block[1409] ^ uncoded_block[1417];
  wire _45079 = _3847 ^ _45078;
  wire _45080 = _45077 ^ _45079;
  wire _45081 = _45076 ^ _45080;
  wire _45082 = _16463 ^ _10683;
  wire _45083 = _5968 ^ _3081;
  wire _45084 = _45082 ^ _45083;
  wire _45085 = uncoded_block[1441] ^ uncoded_block[1444];
  wire _45086 = _45085 ^ _33385;
  wire _45087 = _28352 ^ _45086;
  wire _45088 = _45084 ^ _45087;
  wire _45089 = _45081 ^ _45088;
  wire _45090 = _45073 ^ _45089;
  wire _45091 = _18465 ^ _3088;
  wire _45092 = _18469 ^ _3097;
  wire _45093 = _45091 ^ _45092;
  wire _45094 = _4604 ^ _3884;
  wire _45095 = _5988 ^ _14995;
  wire _45096 = _45094 ^ _45095;
  wire _45097 = _45093 ^ _45096;
  wire _45098 = _9614 ^ _3890;
  wire _45099 = _6634 ^ _1571;
  wire _45100 = _45098 ^ _45099;
  wire _45101 = _18478 ^ _24539;
  wire _45102 = _45101 ^ _38235;
  wire _45103 = _45100 ^ _45102;
  wire _45104 = _45097 ^ _45103;
  wire _45105 = _15004 ^ _8473;
  wire _45106 = _8474 ^ _3905;
  wire _45107 = _45105 ^ _45106;
  wire _45108 = uncoded_block[1542] ^ uncoded_block[1550];
  wire _45109 = _6648 ^ _45108;
  wire _45110 = uncoded_block[1557] ^ uncoded_block[1565];
  wire _45111 = _15020 ^ _45110;
  wire _45112 = _45109 ^ _45111;
  wire _45113 = _45107 ^ _45112;
  wire _45114 = _777 ^ _30870;
  wire _45115 = _45114 ^ _7288;
  wire _45116 = _12369 ^ _2386;
  wire _45117 = uncoded_block[1589] ^ uncoded_block[1597];
  wire _45118 = _5368 ^ _45117;
  wire _45119 = _45116 ^ _45118;
  wire _45120 = _45115 ^ _45119;
  wire _45121 = _45113 ^ _45120;
  wire _45122 = _45104 ^ _45121;
  wire _45123 = _45090 ^ _45122;
  wire _45124 = _3936 ^ _800;
  wire _45125 = _801 ^ _25905;
  wire _45126 = _45124 ^ _45125;
  wire _45127 = _7298 ^ _38668;
  wire _45128 = uncoded_block[1632] ^ uncoded_block[1638];
  wire _45129 = _4667 ^ _45128;
  wire _45130 = _45127 ^ _45129;
  wire _45131 = _45126 ^ _45130;
  wire _45132 = _12383 ^ _5394;
  wire _45133 = _1649 ^ _24578;
  wire _45134 = _45132 ^ _45133;
  wire _45135 = _37891 ^ _9110;
  wire _45136 = _45134 ^ _45135;
  wire _45137 = _45131 ^ _45136;
  wire _45138 = _833 ^ _3190;
  wire _45139 = _9118 ^ _847;
  wire _45140 = _45138 ^ _45139;
  wire _45141 = _852 ^ _17553;
  wire _45142 = _45141 ^ uncoded_block[1722];
  wire _45143 = _45140 ^ _45142;
  wire _45144 = _45137 ^ _45143;
  wire _45145 = _45123 ^ _45144;
  wire _45146 = _45056 ^ _45145;
  wire _45147 = _18057 ^ _7;
  wire _45148 = _21862 ^ _45147;
  wire _45149 = _10226 ^ _27998;
  wire _45150 = _19961 ^ _45149;
  wire _45151 = _45148 ^ _45150;
  wire _45152 = uncoded_block[40] ^ uncoded_block[44];
  wire _45153 = _18 ^ _45152;
  wire _45154 = _31364 ^ _45153;
  wire _45155 = _6099 ^ _7364;
  wire _45156 = _1705 ^ _9705;
  wire _45157 = _45155 ^ _45156;
  wire _45158 = _45154 ^ _45157;
  wire _45159 = _45151 ^ _45158;
  wire _45160 = _39 ^ _14585;
  wire _45161 = _10245 ^ _45160;
  wire _45162 = _11364 ^ _17578;
  wire _45163 = _6755 ^ _19515;
  wire _45164 = _45162 ^ _45163;
  wire _45165 = _45161 ^ _45164;
  wire _45166 = _6758 ^ _9718;
  wire _45167 = _45166 ^ _17083;
  wire _45168 = _2491 ^ _6769;
  wire _45169 = _45168 ^ _15613;
  wire _45170 = _45167 ^ _45169;
  wire _45171 = _45165 ^ _45170;
  wire _45172 = _45159 ^ _45171;
  wire _45173 = _6774 ^ _37141;
  wire _45174 = _12459 ^ _6138;
  wire _45175 = _45173 ^ _45174;
  wire _45176 = uncoded_block[151] ^ uncoded_block[156];
  wire _45177 = _45176 ^ _19040;
  wire _45178 = _45177 ^ _11929;
  wire _45179 = _45175 ^ _45178;
  wire _45180 = _8591 ^ _10270;
  wire _45181 = uncoded_block[180] ^ uncoded_block[192];
  wire _45182 = _45181 ^ _3284;
  wire _45183 = _45180 ^ _45182;
  wire _45184 = _16116 ^ _95;
  wire _45185 = _14101 ^ _7415;
  wire _45186 = _45184 ^ _45185;
  wire _45187 = _45183 ^ _45186;
  wire _45188 = _45179 ^ _45187;
  wire _45189 = _1767 ^ _17613;
  wire _45190 = _15644 ^ _2545;
  wire _45191 = _45189 ^ _45190;
  wire _45192 = _4791 ^ _4081;
  wire _45193 = _8029 ^ _7423;
  wire _45194 = _45192 ^ _45193;
  wire _45195 = _45191 ^ _45194;
  wire _45196 = _1780 ^ _4085;
  wire _45197 = _45196 ^ _31828;
  wire _45198 = _13053 ^ _23746;
  wire _45199 = _1788 ^ _6831;
  wire _45200 = _45198 ^ _45199;
  wire _45201 = _45197 ^ _45200;
  wire _45202 = _45195 ^ _45201;
  wire _45203 = _45188 ^ _45202;
  wire _45204 = _45172 ^ _45203;
  wire _45205 = _22392 ^ _3321;
  wire _45206 = _3324 ^ _6194;
  wire _45207 = _45205 ^ _45206;
  wire _45208 = _988 ^ _1803;
  wire _45209 = _3327 ^ _9226;
  wire _45210 = _45208 ^ _45209;
  wire _45211 = _45207 ^ _45210;
  wire _45212 = uncoded_block[293] ^ uncoded_block[300];
  wire _45213 = _45212 ^ _8052;
  wire _45214 = _1002 ^ _6206;
  wire _45215 = _45213 ^ _45214;
  wire _45216 = _20539 ^ _6852;
  wire _45217 = _45216 ^ _5535;
  wire _45218 = _45215 ^ _45217;
  wire _45219 = _45211 ^ _45218;
  wire _45220 = _1017 ^ _2593;
  wire _45221 = uncoded_block[345] ^ uncoded_block[350];
  wire _45222 = _11450 ^ _45221;
  wire _45223 = _45220 ^ _45222;
  wire _45224 = uncoded_block[356] ^ uncoded_block[362];
  wire _45225 = _45224 ^ _5548;
  wire _45226 = _17163 ^ _17658;
  wire _45227 = _45225 ^ _45226;
  wire _45228 = _45223 ^ _45227;
  wire _45229 = _10895 ^ _10898;
  wire _45230 = _45229 ^ _29679;
  wire _45231 = _5552 ^ _18633;
  wire _45232 = _3383 ^ _1048;
  wire _45233 = _45231 ^ _45232;
  wire _45234 = _45230 ^ _45233;
  wire _45235 = _45228 ^ _45234;
  wire _45236 = _45219 ^ _45235;
  wire _45237 = _4867 ^ _8091;
  wire _45238 = _41115 ^ _45237;
  wire _45239 = _11477 ^ _8672;
  wire _45240 = _39193 ^ _45239;
  wire _45241 = _45238 ^ _45240;
  wire _45242 = _1857 ^ _7497;
  wire _45243 = _1863 ^ _206;
  wire _45244 = _45242 ^ _45243;
  wire _45245 = _4883 ^ _209;
  wire _45246 = _1870 ^ _8681;
  wire _45247 = _45245 ^ _45246;
  wire _45248 = _45244 ^ _45247;
  wire _45249 = _45241 ^ _45248;
  wire _45250 = uncoded_block[468] ^ uncoded_block[473];
  wire _45251 = uncoded_block[477] ^ uncoded_block[482];
  wire _45252 = _45250 ^ _45251;
  wire _45253 = _27763 ^ _45252;
  wire _45254 = _8694 ^ _9291;
  wire _45255 = _1093 ^ _8698;
  wire _45256 = _45254 ^ _45255;
  wire _45257 = _45253 ^ _45256;
  wire _45258 = _229 ^ _9294;
  wire _45259 = _3439 ^ _14193;
  wire _45260 = _45258 ^ _45259;
  wire _45261 = _20097 ^ _1900;
  wire _45262 = _3447 ^ _2683;
  wire _45263 = _45261 ^ _45262;
  wire _45264 = _45260 ^ _45263;
  wire _45265 = _45257 ^ _45264;
  wire _45266 = _45249 ^ _45265;
  wire _45267 = _45236 ^ _45266;
  wire _45268 = _45204 ^ _45267;
  wire _45269 = _24279 ^ _28882;
  wire _45270 = _4931 ^ _8720;
  wire _45271 = _45269 ^ _45270;
  wire _45272 = _25182 ^ _1916;
  wire _45273 = _45272 ^ _38413;
  wire _45274 = _45271 ^ _45273;
  wire _45275 = _262 ^ _18684;
  wire _45276 = _6943 ^ _45275;
  wire _45277 = _9325 ^ _26096;
  wire _45278 = _34013 ^ _6952;
  wire _45279 = _45277 ^ _45278;
  wire _45280 = _45276 ^ _45279;
  wire _45281 = _45274 ^ _45280;
  wire _45282 = _5646 ^ _277;
  wire _45283 = _6323 ^ _6325;
  wire _45284 = _45282 ^ _45283;
  wire _45285 = _5653 ^ _4243;
  wire _45286 = _14224 ^ _1156;
  wire _45287 = _45285 ^ _45286;
  wire _45288 = _45284 ^ _45287;
  wire _45289 = _30199 ^ _38046;
  wire _45290 = _6969 ^ _6336;
  wire _45291 = _45289 ^ _45290;
  wire _45292 = _15766 ^ _3507;
  wire _45293 = _45292 ^ _36021;
  wire _45294 = _45291 ^ _45293;
  wire _45295 = _45288 ^ _45294;
  wire _45296 = _45281 ^ _45295;
  wire _45297 = _15270 ^ _1174;
  wire _45298 = _43772 ^ _8177;
  wire _45299 = _45297 ^ _45298;
  wire _45300 = _44160 ^ _18249;
  wire _45301 = _2754 ^ _8186;
  wire _45302 = _45300 ^ _45301;
  wire _45303 = _45299 ^ _45302;
  wire _45304 = uncoded_block[699] ^ uncoded_block[704];
  wire _45305 = _19195 ^ _45304;
  wire _45306 = _6364 ^ _8190;
  wire _45307 = _45305 ^ _45306;
  wire _45308 = _40044 ^ _5002;
  wire _45309 = _12648 ^ _14774;
  wire _45310 = _45308 ^ _45309;
  wire _45311 = _45307 ^ _45310;
  wire _45312 = _45303 ^ _45311;
  wire _45313 = _7605 ^ _23870;
  wire _45314 = _8202 ^ _45313;
  wire _45315 = _2774 ^ _5012;
  wire _45316 = _5013 ^ _35254;
  wire _45317 = _45315 ^ _45316;
  wire _45318 = _45314 ^ _45317;
  wire _45319 = _4301 ^ _14788;
  wire _45320 = _17775 ^ _45319;
  wire _45321 = _5711 ^ _2015;
  wire _45322 = _45321 ^ _32378;
  wire _45323 = _45320 ^ _45322;
  wire _45324 = _45318 ^ _45323;
  wire _45325 = _45312 ^ _45324;
  wire _45326 = _45296 ^ _45325;
  wire _45327 = _18283 ^ _375;
  wire _45328 = _7628 ^ _385;
  wire _45329 = _45327 ^ _45328;
  wire _45330 = uncoded_block[809] ^ uncoded_block[814];
  wire _45331 = _32381 ^ _45330;
  wire _45332 = uncoded_block[819] ^ uncoded_block[821];
  wire _45333 = _2808 ^ _45332;
  wire _45334 = _45331 ^ _45333;
  wire _45335 = _45329 ^ _45334;
  wire _45336 = uncoded_block[831] ^ uncoded_block[836];
  wire _45337 = _5052 ^ _45336;
  wire _45338 = uncoded_block[843] ^ uncoded_block[849];
  wire _45339 = _22532 ^ _45338;
  wire _45340 = _45337 ^ _45339;
  wire _45341 = _14814 ^ _24357;
  wire _45342 = _5066 ^ _7649;
  wire _45343 = _45341 ^ _45342;
  wire _45344 = _45340 ^ _45343;
  wire _45345 = _45335 ^ _45344;
  wire _45346 = uncoded_block[866] ^ uncoded_block[870];
  wire _45347 = _5069 ^ _45346;
  wire _45348 = _12696 ^ _2831;
  wire _45349 = _45347 ^ _45348;
  wire _45350 = _2053 ^ _2836;
  wire _45351 = _1272 ^ _9416;
  wire _45352 = _45350 ^ _45351;
  wire _45353 = _45349 ^ _45352;
  wire _45354 = _20701 ^ _19735;
  wire _45355 = uncoded_block[898] ^ uncoded_block[903];
  wire _45356 = _45355 ^ _9421;
  wire _45357 = _45354 ^ _45356;
  wire _45358 = _2071 ^ _6430;
  wire _45359 = _3629 ^ _4368;
  wire _45360 = _45358 ^ _45359;
  wire _45361 = _45357 ^ _45360;
  wire _45362 = _45353 ^ _45361;
  wire _45363 = _45345 ^ _45362;
  wire _45364 = uncoded_block[932] ^ uncoded_block[937];
  wire _45365 = _1296 ^ _45364;
  wire _45366 = _6439 ^ _8271;
  wire _45367 = _45365 ^ _45366;
  wire _45368 = _5777 ^ _4381;
  wire _45369 = _5779 ^ _10529;
  wire _45370 = _45368 ^ _45369;
  wire _45371 = _45367 ^ _45370;
  wire _45372 = _22112 ^ _25283;
  wire _45373 = _32425 ^ _17836;
  wire _45374 = _45372 ^ _45373;
  wire _45375 = _4397 ^ _15369;
  wire _45376 = _2882 ^ _4401;
  wire _45377 = _45375 ^ _45376;
  wire _45378 = _45374 ^ _45377;
  wire _45379 = _45371 ^ _45378;
  wire _45380 = uncoded_block[1003] ^ uncoded_block[1007];
  wire _45381 = _9449 ^ _45380;
  wire _45382 = _19759 ^ _45381;
  wire _45383 = _5132 ^ _38127;
  wire _45384 = _45382 ^ _45383;
  wire _45385 = _495 ^ _13288;
  wire _45386 = _2907 ^ _7707;
  wire _45387 = _45385 ^ _45386;
  wire _45388 = _2133 ^ _19295;
  wire _45389 = _1347 ^ _45388;
  wire _45390 = _45387 ^ _45389;
  wire _45391 = _45384 ^ _45390;
  wire _45392 = _45379 ^ _45391;
  wire _45393 = _45363 ^ _45392;
  wire _45394 = _45326 ^ _45393;
  wire _45395 = _45268 ^ _45394;
  wire _45396 = uncoded_block[1052] ^ uncoded_block[1058];
  wire _45397 = _45396 ^ _13849;
  wire _45398 = _1366 ^ _13307;
  wire _45399 = _45397 ^ _45398;
  wire _45400 = _5834 ^ _21687;
  wire _45401 = _5839 ^ _537;
  wire _45402 = _45400 ^ _45401;
  wire _45403 = _45399 ^ _45402;
  wire _45404 = _5169 ^ _3707;
  wire _45405 = _34942 ^ _45404;
  wire _45406 = _26231 ^ _7735;
  wire _45407 = _45405 ^ _45406;
  wire _45408 = _45403 ^ _45407;
  wire _45409 = _11147 ^ _10587;
  wire _45410 = _2172 ^ _4459;
  wire _45411 = _45409 ^ _45410;
  wire _45412 = _8343 ^ _14887;
  wire _45413 = _8346 ^ _5859;
  wire _45414 = _45412 ^ _45413;
  wire _45415 = _45411 ^ _45414;
  wire _45416 = _3736 ^ _7154;
  wire _45417 = _45416 ^ _7753;
  wire _45418 = _27545 ^ _35749;
  wire _45419 = _24910 ^ _7160;
  wire _45420 = _45418 ^ _45419;
  wire _45421 = _45417 ^ _45420;
  wire _45422 = _45415 ^ _45421;
  wire _45423 = _45408 ^ _45422;
  wire _45424 = _7162 ^ _5207;
  wire _45425 = _6530 ^ _33750;
  wire _45426 = _45424 ^ _45425;
  wire _45427 = _45036 ^ _5894;
  wire _45428 = _43516 ^ _45427;
  wire _45429 = _45426 ^ _45428;
  wire _45430 = _33758 ^ _1451;
  wire _45431 = _45430 ^ _18862;
  wire _45432 = _30781 ^ _45431;
  wire _45433 = _45429 ^ _45432;
  wire _45434 = _20801 ^ _3003;
  wire _45435 = _11188 ^ _628;
  wire _45436 = _45434 ^ _45435;
  wire _45437 = _2247 ^ _4525;
  wire _45438 = _45437 ^ _19368;
  wire _45439 = _45436 ^ _45438;
  wire _45440 = uncoded_block[1295] ^ uncoded_block[1301];
  wire _45441 = _10646 ^ _45440;
  wire _45442 = _45441 ^ _15948;
  wire _45443 = _14430 ^ _654;
  wire _45444 = uncoded_block[1323] ^ uncoded_block[1330];
  wire _45445 = _45444 ^ _4550;
  wire _45446 = _45443 ^ _45445;
  wire _45447 = _45442 ^ _45446;
  wire _45448 = _45439 ^ _45447;
  wire _45449 = _45433 ^ _45448;
  wire _45450 = _45423 ^ _45449;
  wire _45451 = _4553 ^ _5262;
  wire _45452 = _45451 ^ _25842;
  wire _45453 = _29930 ^ _5273;
  wire _45454 = _27157 ^ _11224;
  wire _45455 = _45453 ^ _45454;
  wire _45456 = _45452 ^ _45455;
  wire _45457 = _3832 ^ _20334;
  wire _45458 = uncoded_block[1385] ^ uncoded_block[1395];
  wire _45459 = _687 ^ _45458;
  wire _45460 = _45457 ^ _45459;
  wire _45461 = _5955 ^ _1517;
  wire _45462 = _14457 ^ _701;
  wire _45463 = _45461 ^ _45462;
  wire _45464 = _45460 ^ _45463;
  wire _45465 = _45456 ^ _45464;
  wire _45466 = _5964 ^ _2308;
  wire _45467 = _38617 ^ _45466;
  wire _45468 = _9590 ^ _3856;
  wire _45469 = _45468 ^ _39026;
  wire _45470 = _45467 ^ _45469;
  wire _45471 = _5304 ^ _2321;
  wire _45472 = _9033 ^ _3865;
  wire _45473 = _45471 ^ _45472;
  wire _45474 = _12332 ^ _22252;
  wire _45475 = _45474 ^ _2337;
  wire _45476 = _45473 ^ _45475;
  wire _45477 = _45470 ^ _45476;
  wire _45478 = _45465 ^ _45477;
  wire _45479 = _3094 ^ _1551;
  wire _45480 = uncoded_block[1473] ^ uncoded_block[1480];
  wire _45481 = _45480 ^ _10706;
  wire _45482 = _45479 ^ _45481;
  wire _45483 = _3103 ^ _6631;
  wire _45484 = _45483 ^ _23189;
  wire _45485 = _45482 ^ _45484;
  wire _45486 = uncoded_block[1510] ^ uncoded_block[1516];
  wire _45487 = _45486 ^ _9624;
  wire _45488 = _9049 ^ _45487;
  wire _45489 = _2360 ^ _16008;
  wire _45490 = _42535 ^ _45489;
  wire _45491 = _45488 ^ _45490;
  wire _45492 = _45485 ^ _45491;
  wire _45493 = _5348 ^ _29125;
  wire _45494 = _45493 ^ _35440;
  wire _45495 = _6015 ^ _4638;
  wire _45496 = uncoded_block[1561] ^ uncoded_block[1566];
  wire _45497 = _45496 ^ _17007;
  wire _45498 = _45495 ^ _45497;
  wire _45499 = _45494 ^ _45498;
  wire _45500 = _784 ^ _17009;
  wire _45501 = _12928 ^ _45500;
  wire _45502 = uncoded_block[1592] ^ uncoded_block[1597];
  wire _45503 = _45502 ^ _1621;
  wire _45504 = _17012 ^ _45503;
  wire _45505 = _45501 ^ _45504;
  wire _45506 = _45499 ^ _45505;
  wire _45507 = _45492 ^ _45506;
  wire _45508 = _45478 ^ _45507;
  wire _45509 = _45450 ^ _45508;
  wire _45510 = uncoded_block[1608] ^ uncoded_block[1613];
  wire _45511 = _14517 ^ _45510;
  wire _45512 = _45511 ^ _18508;
  wire _45513 = uncoded_block[1622] ^ uncoded_block[1625];
  wire _45514 = _45513 ^ _12947;
  wire _45515 = _1636 ^ _9659;
  wire _45516 = _45514 ^ _45515;
  wire _45517 = _45512 ^ _45516;
  wire _45518 = _3948 ^ _27651;
  wire _45519 = _45518 ^ _42182;
  wire _45520 = _29569 ^ _5399;
  wire _45521 = _26824 ^ _45520;
  wire _45522 = _45519 ^ _45521;
  wire _45523 = _45517 ^ _45522;
  wire _45524 = _7928 ^ _830;
  wire _45525 = uncoded_block[1679] ^ uncoded_block[1685];
  wire _45526 = _832 ^ _45525;
  wire _45527 = _45524 ^ _45526;
  wire _45528 = _1665 ^ _11325;
  wire _45529 = _45528 ^ _35476;
  wire _45530 = _45527 ^ _45529;
  wire _45531 = _4700 ^ _2435;
  wire _45532 = _45531 ^ _30905;
  wire _45533 = _14553 ^ _18992;
  wire _45534 = _45532 ^ _45533;
  wire _45535 = _45530 ^ _45534;
  wire _45536 = _45523 ^ _45535;
  wire _45537 = _45536 ^ uncoded_block[1722];
  wire _45538 = _45509 ^ _45537;
  wire _45539 = _45395 ^ _45538;
  wire _45540 = _3209 ^ _3993;
  wire _45541 = uncoded_block[10] ^ uncoded_block[15];
  wire _45542 = _3995 ^ _45541;
  wire _45543 = _45540 ^ _45542;
  wire _45544 = _39881 ^ _11345;
  wire _45545 = _45543 ^ _45544;
  wire _45546 = _21871 ^ _15591;
  wire _45547 = _11891 ^ _45546;
  wire _45548 = _23 ^ _3233;
  wire _45549 = _42858 ^ _7364;
  wire _45550 = _45548 ^ _45549;
  wire _45551 = _45547 ^ _45550;
  wire _45552 = _45545 ^ _45551;
  wire _45553 = _901 ^ _19019;
  wire _45554 = _41443 ^ _45553;
  wire _45555 = _11364 ^ _6755;
  wire _45556 = uncoded_block[89] ^ uncoded_block[95];
  wire _45557 = _45556 ^ _9718;
  wire _45558 = _45555 ^ _45557;
  wire _45559 = _45554 ^ _45558;
  wire _45560 = _19025 ^ _14595;
  wire _45561 = _2491 ^ _3253;
  wire _45562 = _45560 ^ _45561;
  wire _45563 = _16592 ^ _56;
  wire _45564 = _2502 ^ _4753;
  wire _45565 = _45563 ^ _45564;
  wire _45566 = _45562 ^ _45565;
  wire _45567 = _45559 ^ _45566;
  wire _45568 = _45552 ^ _45567;
  wire _45569 = _3263 ^ _9729;
  wire _45570 = _39124 ^ _45569;
  wire _45571 = _11918 ^ _17097;
  wire _45572 = _1744 ^ _73;
  wire _45573 = _45571 ^ _45572;
  wire _45574 = _45570 ^ _45573;
  wire _45575 = _19536 ^ _81;
  wire _45576 = _23726 ^ _45575;
  wire _45577 = _14093 ^ _33076;
  wire _45578 = _45576 ^ _45577;
  wire _45579 = _45574 ^ _45578;
  wire _45580 = _14616 ^ _33077;
  wire _45581 = _13590 ^ _12479;
  wire _45582 = _45580 ^ _45581;
  wire _45583 = _955 ^ _19549;
  wire _45584 = _27295 ^ _10854;
  wire _45585 = _45583 ^ _45584;
  wire _45586 = _45582 ^ _45585;
  wire _45587 = uncoded_block[226] ^ uncoded_block[229];
  wire _45588 = _45587 ^ _30087;
  wire _45589 = _45588 ^ _22852;
  wire _45590 = _5505 ^ _7434;
  wire _45591 = _14117 ^ _14639;
  wire _45592 = _45590 ^ _45591;
  wire _45593 = _45589 ^ _45592;
  wire _45594 = _45586 ^ _45593;
  wire _45595 = _45579 ^ _45594;
  wire _45596 = _45568 ^ _45595;
  wire _45597 = _25108 ^ _20523;
  wire _45598 = _985 ^ _10872;
  wire _45599 = _45597 ^ _45598;
  wire _45600 = _27716 ^ _24212;
  wire _45601 = _11965 ^ _45600;
  wire _45602 = _45599 ^ _45601;
  wire _45603 = _9226 ^ _3328;
  wire _45604 = _17142 ^ _17144;
  wire _45605 = _45603 ^ _45604;
  wire _45606 = _3337 ^ _14654;
  wire _45607 = _10314 ^ _45606;
  wire _45608 = _45605 ^ _45607;
  wire _45609 = _45602 ^ _45608;
  wire _45610 = _4830 ^ _1009;
  wire _45611 = _12521 ^ _1822;
  wire _45612 = _45610 ^ _45611;
  wire _45613 = _1825 ^ _1021;
  wire _45614 = _6218 ^ _4844;
  wire _45615 = _45613 ^ _45614;
  wire _45616 = _45612 ^ _45615;
  wire _45617 = _31437 ^ _27737;
  wire _45618 = _5548 ^ _7470;
  wire _45619 = uncoded_block[371] ^ uncoded_block[377];
  wire _45620 = _1835 ^ _45619;
  wire _45621 = _45618 ^ _45620;
  wire _45622 = _45617 ^ _45621;
  wire _45623 = _45616 ^ _45622;
  wire _45624 = _45609 ^ _45623;
  wire _45625 = _10901 ^ _4149;
  wire _45626 = _3381 ^ _19604;
  wire _45627 = _45625 ^ _45626;
  wire _45628 = _7487 ^ _13106;
  wire _45629 = _41114 ^ _45628;
  wire _45630 = _45627 ^ _45629;
  wire _45631 = _19612 ^ _7492;
  wire _45632 = _8664 ^ _45631;
  wire _45633 = _2639 ^ _42297;
  wire _45634 = _45632 ^ _45633;
  wire _45635 = _45630 ^ _45634;
  wire _45636 = _4882 ^ _209;
  wire _45637 = _212 ^ _13127;
  wire _45638 = _45636 ^ _45637;
  wire _45639 = _23356 ^ _34384;
  wire _45640 = _45638 ^ _45639;
  wire _45641 = uncoded_block[471] ^ uncoded_block[477];
  wire _45642 = _45641 ^ _1085;
  wire _45643 = _8694 ^ _6276;
  wire _45644 = _45642 ^ _45643;
  wire _45645 = _10937 ^ _8698;
  wire _45646 = _229 ^ _1892;
  wire _45647 = _45645 ^ _45646;
  wire _45648 = _45644 ^ _45647;
  wire _45649 = _45640 ^ _45648;
  wire _45650 = _45635 ^ _45649;
  wire _45651 = _45624 ^ _45650;
  wire _45652 = _45596 ^ _45651;
  wire _45653 = _19137 ^ _26511;
  wire _45654 = _3444 ^ _4921;
  wire _45655 = _6929 ^ _3450;
  wire _45656 = _45654 ^ _45655;
  wire _45657 = _45653 ^ _45656;
  wire _45658 = _4217 ^ _8132;
  wire _45659 = _1117 ^ _6300;
  wire _45660 = _45658 ^ _45659;
  wire _45661 = _24284 ^ _32736;
  wire _45662 = _16719 ^ _45661;
  wire _45663 = _45660 ^ _45662;
  wire _45664 = _45657 ^ _45663;
  wire _45665 = _13165 ^ _13168;
  wire _45666 = _1132 ^ _9325;
  wire _45667 = _45665 ^ _45666;
  wire _45668 = _20116 ^ _34013;
  wire _45669 = _45668 ^ _20620;
  wire _45670 = _45667 ^ _45669;
  wire _45671 = _17232 ^ _1149;
  wire _45672 = _43757 ^ _45671;
  wire _45673 = _281 ^ _16738;
  wire _45674 = _45673 ^ _14746;
  wire _45675 = _45672 ^ _45674;
  wire _45676 = _45670 ^ _45675;
  wire _45677 = _45664 ^ _45676;
  wire _45678 = _290 ^ _293;
  wire _45679 = _45678 ^ _12077;
  wire _45680 = _9350 ^ _21111;
  wire _45681 = _6339 ^ _45680;
  wire _45682 = _45679 ^ _45681;
  wire _45683 = _20638 ^ _21113;
  wire _45684 = _28158 ^ _1178;
  wire _45685 = _45683 ^ _45684;
  wire _45686 = _8760 ^ _1971;
  wire _45687 = _45686 ^ _38443;
  wire _45688 = _45685 ^ _45687;
  wire _45689 = _45682 ^ _45688;
  wire _45690 = _41966 ^ _5682;
  wire _45691 = uncoded_block[700] ^ uncoded_block[703];
  wire _45692 = _6360 ^ _45691;
  wire _45693 = _11564 ^ _4996;
  wire _45694 = _45692 ^ _45693;
  wire _45695 = _45690 ^ _45694;
  wire _45696 = _4998 ^ _5002;
  wire _45697 = _30221 ^ _3544;
  wire _45698 = _45696 ^ _45697;
  wire _45699 = _344 ^ _7001;
  wire _45700 = _12653 ^ _7005;
  wire _45701 = _45699 ^ _45700;
  wire _45702 = _45698 ^ _45701;
  wire _45703 = _45695 ^ _45702;
  wire _45704 = _45689 ^ _45703;
  wire _45705 = _45677 ^ _45704;
  wire _45706 = _41195 ^ _15794;
  wire _45707 = _4299 ^ _364;
  wire _45708 = _44572 ^ _45707;
  wire _45709 = _45706 ^ _45708;
  wire _45710 = _14271 ^ _13216;
  wire _45711 = _8786 ^ _45710;
  wire _45712 = _31106 ^ _1224;
  wire _45713 = _20166 ^ _45712;
  wire _45714 = _45711 ^ _45713;
  wire _45715 = _45709 ^ _45714;
  wire _45716 = uncoded_block[793] ^ uncoded_block[800];
  wire _45717 = _5033 ^ _45716;
  wire _45718 = _9394 ^ _392;
  wire _45719 = _45717 ^ _45718;
  wire _45720 = _2806 ^ _14291;
  wire _45721 = _400 ^ _9402;
  wire _45722 = _45720 ^ _45721;
  wire _45723 = _45719 ^ _45722;
  wire _45724 = uncoded_block[836] ^ uncoded_block[839];
  wire _45725 = _45724 ^ _1256;
  wire _45726 = _33239 ^ _6406;
  wire _45727 = _45725 ^ _45726;
  wire _45728 = _4343 ^ _5066;
  wire _45729 = _6412 ^ _5071;
  wire _45730 = _45728 ^ _45729;
  wire _45731 = _45727 ^ _45730;
  wire _45732 = _45723 ^ _45731;
  wire _45733 = _45715 ^ _45732;
  wire _45734 = _4346 ^ _12151;
  wire _45735 = _16304 ^ _2836;
  wire _45736 = _45734 ^ _45735;
  wire _45737 = _14821 ^ _9416;
  wire _45738 = uncoded_block[891] ^ uncoded_block[895];
  wire _45739 = _45738 ^ _5758;
  wire _45740 = _45737 ^ _45739;
  wire _45741 = _45736 ^ _45740;
  wire _45742 = _3617 ^ _5090;
  wire _45743 = _12708 ^ _3629;
  wire _45744 = _45742 ^ _45743;
  wire _45745 = _446 ^ _448;
  wire _45746 = _3633 ^ _45745;
  wire _45747 = _45744 ^ _45746;
  wire _45748 = _45741 ^ _45747;
  wire _45749 = _8262 ^ _2862;
  wire _45750 = _2083 ^ _453;
  wire _45751 = _45749 ^ _45750;
  wire _45752 = uncoded_block[951] ^ uncoded_block[957];
  wire _45753 = uncoded_block[958] ^ uncoded_block[961];
  wire _45754 = _45752 ^ _45753;
  wire _45755 = _24385 ^ _45754;
  wire _45756 = _45751 ^ _45755;
  wire _45757 = uncoded_block[968] ^ uncoded_block[973];
  wire _45758 = _12180 ^ _45757;
  wire _45759 = _5114 ^ _5790;
  wire _45760 = _45758 ^ _45759;
  wire _45761 = uncoded_block[989] ^ uncoded_block[997];
  wire _45762 = _8287 ^ _45761;
  wire _45763 = _45762 ^ _16849;
  wire _45764 = _45760 ^ _45763;
  wire _45765 = _45756 ^ _45764;
  wire _45766 = _45748 ^ _45765;
  wire _45767 = _45733 ^ _45766;
  wire _45768 = _45705 ^ _45767;
  wire _45769 = _45652 ^ _45768;
  wire _45770 = _9996 ^ _5135;
  wire _45771 = _15861 ^ _45770;
  wire _45772 = _4417 ^ _22595;
  wire _45773 = _12195 ^ _45772;
  wire _45774 = _45771 ^ _45773;
  wire _45775 = _1346 ^ _512;
  wire _45776 = _45775 ^ _13293;
  wire _45777 = _13844 ^ _11116;
  wire _45778 = _45777 ^ _40129;
  wire _45779 = _45776 ^ _45778;
  wire _45780 = _45774 ^ _45779;
  wire _45781 = _526 ^ _12217;
  wire _45782 = _2924 ^ _3695;
  wire _45783 = _45781 ^ _45782;
  wire _45784 = _11687 ^ _30740;
  wire _45785 = _45784 ^ _34527;
  wire _45786 = _45783 ^ _45785;
  wire _45787 = _4444 ^ _9484;
  wire _45788 = _4450 ^ _25323;
  wire _45789 = _45787 ^ _45788;
  wire _45790 = uncoded_block[1119] ^ uncoded_block[1123];
  wire _45791 = _1388 ^ _45790;
  wire _45792 = uncoded_block[1130] ^ uncoded_block[1140];
  wire _45793 = _12791 ^ _45792;
  wire _45794 = _45791 ^ _45793;
  wire _45795 = _45789 ^ _45794;
  wire _45796 = _45786 ^ _45795;
  wire _45797 = _45780 ^ _45796;
  wire _45798 = _40893 ^ _14384;
  wire _45799 = _11711 ^ _17389;
  wire _45800 = _17390 ^ _10602;
  wire _45801 = _45799 ^ _45800;
  wire _45802 = _45798 ^ _45801;
  wire _45803 = _16901 ^ _5201;
  wire _45804 = _36572 ^ _45803;
  wire _45805 = _12808 ^ _3749;
  wire _45806 = _45805 ^ _27908;
  wire _45807 = _45804 ^ _45806;
  wire _45808 = _45802 ^ _45807;
  wire _45809 = _24001 ^ _2982;
  wire _45810 = _2211 ^ _45809;
  wire _45811 = _43894 ^ _42463;
  wire _45812 = _45810 ^ _45811;
  wire _45813 = _2989 ^ _17910;
  wire _45814 = _6538 ^ _1451;
  wire _45815 = _45813 ^ _45814;
  wire _45816 = _7778 ^ _11739;
  wire _45817 = _45816 ^ _29466;
  wire _45818 = _45815 ^ _45817;
  wire _45819 = _45812 ^ _45818;
  wire _45820 = _45808 ^ _45819;
  wire _45821 = _45797 ^ _45820;
  wire _45822 = uncoded_block[1273] ^ uncoded_block[1278];
  wire _45823 = uncoded_block[1279] ^ uncoded_block[1284];
  wire _45824 = _45822 ^ _45823;
  wire _45825 = _44688 ^ _45824;
  wire _45826 = uncoded_block[1289] ^ uncoded_block[1292];
  wire _45827 = _45826 ^ _7194;
  wire _45828 = _37808 ^ _45827;
  wire _45829 = _45825 ^ _45828;
  wire _45830 = _2254 ^ _7196;
  wire _45831 = _37813 ^ _656;
  wire _45832 = _45830 ^ _45831;
  wire _45833 = _6579 ^ _8414;
  wire _45834 = _45832 ^ _45833;
  wire _45835 = _45829 ^ _45834;
  wire _45836 = _3041 ^ _1502;
  wire _45837 = _22677 ^ _45836;
  wire _45838 = _6587 ^ _27157;
  wire _45839 = _11224 ^ _22224;
  wire _45840 = _45838 ^ _45839;
  wire _45841 = _45837 ^ _45840;
  wire _45842 = _5284 ^ _32935;
  wire _45843 = _6596 ^ _5950;
  wire _45844 = _45842 ^ _45843;
  wire _45845 = uncoded_block[1394] ^ uncoded_block[1402];
  wire _45846 = _5952 ^ _45845;
  wire _45847 = _4578 ^ _8436;
  wire _45848 = _45846 ^ _45847;
  wire _45849 = _45844 ^ _45848;
  wire _45850 = _45841 ^ _45849;
  wire _45851 = _45835 ^ _45850;
  wire _45852 = _702 ^ _13422;
  wire _45853 = _10118 ^ _9021;
  wire _45854 = _45852 ^ _45853;
  wire _45855 = uncoded_block[1423] ^ uncoded_block[1429];
  wire _45856 = _45855 ^ _1531;
  wire _45857 = _8443 ^ _2318;
  wire _45858 = _45856 ^ _45857;
  wire _45859 = _45854 ^ _45858;
  wire _45860 = _6614 ^ _43570;
  wire _45861 = uncoded_block[1467] ^ uncoded_block[1473];
  wire _45862 = _3094 ^ _45861;
  wire _45863 = _37454 ^ _45862;
  wire _45864 = _45860 ^ _45863;
  wire _45865 = _45859 ^ _45864;
  wire _45866 = _32135 ^ _23621;
  wire _45867 = _9044 ^ _3890;
  wire _45868 = uncoded_block[1501] ^ uncoded_block[1509];
  wire _45869 = _3109 ^ _45868;
  wire _45870 = _45867 ^ _45869;
  wire _45871 = _45866 ^ _45870;
  wire _45872 = _7264 ^ _2357;
  wire _45873 = _3900 ^ _11820;
  wire _45874 = _45872 ^ _45873;
  wire _45875 = _5347 ^ _6650;
  wire _45876 = _758 ^ _4634;
  wire _45877 = _45875 ^ _45876;
  wire _45878 = _45874 ^ _45877;
  wire _45879 = _45871 ^ _45878;
  wire _45880 = _45865 ^ _45879;
  wire _45881 = _45851 ^ _45880;
  wire _45882 = _45821 ^ _45881;
  wire _45883 = _35439 ^ _7277;
  wire _45884 = _9070 ^ _6016;
  wire _45885 = _45883 ^ _45884;
  wire _45886 = uncoded_block[1561] ^ uncoded_block[1565];
  wire _45887 = _45886 ^ _11284;
  wire _45888 = _26337 ^ _4648;
  wire _45889 = _45887 ^ _45888;
  wire _45890 = _45885 ^ _45889;
  wire _45891 = _2386 ^ _14511;
  wire _45892 = _27640 ^ _45891;
  wire _45893 = _11294 ^ _797;
  wire _45894 = _41782 ^ _45893;
  wire _45895 = _45892 ^ _45894;
  wire _45896 = _45890 ^ _45895;
  wire _45897 = _8502 ^ _6677;
  wire _45898 = _3937 ^ _6679;
  wire _45899 = _45897 ^ _45898;
  wire _45900 = _5383 ^ _29557;
  wire _45901 = _45900 ^ _40640;
  wire _45902 = _45899 ^ _45901;
  wire _45903 = _10754 ^ _12383;
  wire _45904 = _4673 ^ _1649;
  wire _45905 = _45903 ^ _45904;
  wire _45906 = _3172 ^ _820;
  wire _45907 = _3174 ^ _29569;
  wire _45908 = _45906 ^ _45907;
  wire _45909 = _45905 ^ _45908;
  wire _45910 = _45902 ^ _45909;
  wire _45911 = _45896 ^ _45910;
  wire _45912 = _2419 ^ _19466;
  wire _45913 = uncoded_block[1671] ^ uncoded_block[1677];
  wire _45914 = _6058 ^ _45913;
  wire _45915 = _45912 ^ _45914;
  wire _45916 = _836 ^ _3190;
  wire _45917 = _20428 ^ _45916;
  wire _45918 = _45915 ^ _45917;
  wire _45919 = _42840 ^ _27233;
  wire _45920 = _44408 ^ _2441;
  wire _45921 = _45920 ^ _7947;
  wire _45922 = _45919 ^ _45921;
  wire _45923 = _45918 ^ _45922;
  wire _45924 = _45911 ^ _45923;
  wire _45925 = _45882 ^ _45924;
  wire _45926 = _45769 ^ _45925;
  wire _45927 = _9688 ^ _8545;
  wire _45928 = _3217 ^ _2462;
  wire _45929 = _45927 ^ _45928;
  wire _45930 = _12994 ^ _31790;
  wire _45931 = uncoded_block[64] ^ uncoded_block[75];
  wire _45932 = _45931 ^ _25957;
  wire _45933 = _45930 ^ _45932;
  wire _45934 = _45929 ^ _45933;
  wire _45935 = uncoded_block[93] ^ uncoded_block[110];
  wire _45936 = _45935 ^ _56;
  wire _45937 = uncoded_block[130] ^ uncoded_block[141];
  wire _45938 = uncoded_block[149] ^ uncoded_block[160];
  wire _45939 = _45937 ^ _45938;
  wire _45940 = _45936 ^ _45939;
  wire _45941 = _6787 ^ _4770;
  wire _45942 = uncoded_block[187] ^ uncoded_block[193];
  wire _45943 = uncoded_block[194] ^ uncoded_block[200];
  wire _45944 = _45942 ^ _45943;
  wire _45945 = _45941 ^ _45944;
  wire _45946 = _45940 ^ _45945;
  wire _45947 = _45934 ^ _45946;
  wire _45948 = uncoded_block[207] ^ uncoded_block[216];
  wire _45949 = _1764 ^ _45948;
  wire _45950 = uncoded_block[226] ^ uncoded_block[235];
  wire _45951 = _14105 ^ _45950;
  wire _45952 = _45949 ^ _45951;
  wire _45953 = _6180 ^ _10297;
  wire _45954 = uncoded_block[263] ^ uncoded_block[276];
  wire _45955 = _45954 ^ _30104;
  wire _45956 = _45953 ^ _45955;
  wire _45957 = _45952 ^ _45956;
  wire _45958 = uncoded_block[291] ^ uncoded_block[303];
  wire _45959 = _9226 ^ _45958;
  wire _45960 = uncoded_block[320] ^ uncoded_block[331];
  wire _45961 = _15671 ^ _45960;
  wire _45962 = _45959 ^ _45961;
  wire _45963 = uncoded_block[338] ^ uncoded_block[349];
  wire _45964 = _11446 ^ _45963;
  wire _45965 = uncoded_block[355] ^ uncoded_block[361];
  wire _45966 = _1028 ^ _45965;
  wire _45967 = _45964 ^ _45966;
  wire _45968 = _45962 ^ _45967;
  wire _45969 = _45957 ^ _45968;
  wire _45970 = _45947 ^ _45969;
  wire _45971 = _8076 ^ _4858;
  wire _45972 = uncoded_block[397] ^ uncoded_block[402];
  wire _45973 = _2616 ^ _45972;
  wire _45974 = _45971 ^ _45973;
  wire _45975 = uncoded_block[418] ^ uncoded_block[431];
  wire _45976 = _36796 ^ _45975;
  wire _45977 = _10352 ^ _1076;
  wire _45978 = _45976 ^ _45977;
  wire _45979 = _45974 ^ _45978;
  wire _45980 = uncoded_block[466] ^ uncoded_block[471];
  wire _45981 = _11491 ^ _45980;
  wire _45982 = uncoded_block[488] ^ uncoded_block[495];
  wire _45983 = _4188 ^ _45982;
  wire _45984 = _45981 ^ _45983;
  wire _45985 = uncoded_block[507] ^ uncoded_block[512];
  wire _45986 = _1097 ^ _45985;
  wire _45987 = uncoded_block[520] ^ uncoded_block[525];
  wire _45988 = uncoded_block[535] ^ uncoded_block[541];
  wire _45989 = _45987 ^ _45988;
  wire _45990 = _45986 ^ _45989;
  wire _45991 = _45984 ^ _45990;
  wire _45992 = _45979 ^ _45991;
  wire _45993 = uncoded_block[548] ^ uncoded_block[554];
  wire _45994 = _45993 ^ _12051;
  wire _45995 = _7545 ^ _3468;
  wire _45996 = _45994 ^ _45995;
  wire _45997 = _10969 ^ _2701;
  wire _45998 = uncoded_block[599] ^ uncoded_block[614];
  wire _45999 = uncoded_block[627] ^ uncoded_block[635];
  wire _46000 = _45998 ^ _45999;
  wire _46001 = _45997 ^ _46000;
  wire _46002 = _45996 ^ _46001;
  wire _46003 = uncoded_block[653] ^ uncoded_block[666];
  wire _46004 = uncoded_block[669] ^ uncoded_block[678];
  wire _46005 = _46003 ^ _46004;
  wire _46006 = _7579 ^ _46005;
  wire _46007 = uncoded_block[692] ^ uncoded_block[706];
  wire _46008 = _15281 ^ _46007;
  wire _46009 = _33205 ^ _12647;
  wire _46010 = _46008 ^ _46009;
  wire _46011 = _46006 ^ _46010;
  wire _46012 = _46002 ^ _46011;
  wire _46013 = _45992 ^ _46012;
  wire _46014 = _45970 ^ _46013;
  wire _46015 = uncoded_block[734] ^ uncoded_block[744];
  wire _46016 = uncoded_block[747] ^ uncoded_block[758];
  wire _46017 = _46015 ^ _46016;
  wire _46018 = _1992 ^ _46017;
  wire _46019 = uncoded_block[780] ^ uncoded_block[787];
  wire _46020 = _2784 ^ _46019;
  wire _46021 = _2021 ^ _7029;
  wire _46022 = _46020 ^ _46021;
  wire _46023 = _46018 ^ _46022;
  wire _46024 = _32381 ^ _2028;
  wire _46025 = _27843 ^ _27846;
  wire _46026 = _46024 ^ _46025;
  wire _46027 = uncoded_block[862] ^ uncoded_block[868];
  wire _46028 = _8809 ^ _46027;
  wire _46029 = uncoded_block[877] ^ uncoded_block[883];
  wire _46030 = _11620 ^ _46029;
  wire _46031 = _46028 ^ _46030;
  wire _46032 = _46026 ^ _46031;
  wire _46033 = _46023 ^ _46032;
  wire _46034 = _4352 ^ _45738;
  wire _46035 = uncoded_block[900] ^ uncoded_block[904];
  wire _46036 = _8826 ^ _46035;
  wire _46037 = _46034 ^ _46036;
  wire _46038 = uncoded_block[910] ^ uncoded_block[924];
  wire _46039 = uncoded_block[925] ^ uncoded_block[945];
  wire _46040 = _46038 ^ _46039;
  wire _46041 = uncoded_block[960] ^ uncoded_block[971];
  wire _46042 = uncoded_block[978] ^ uncoded_block[986];
  wire _46043 = _46041 ^ _46042;
  wire _46044 = _46040 ^ _46043;
  wire _46045 = _46037 ^ _46044;
  wire _46046 = uncoded_block[1000] ^ uncoded_block[1006];
  wire _46047 = _4398 ^ _46046;
  wire _46048 = uncoded_block[1010] ^ uncoded_block[1016];
  wire _46049 = _46048 ^ _2894;
  wire _46050 = _46047 ^ _46049;
  wire _46051 = uncoded_block[1037] ^ uncoded_block[1046];
  wire _46052 = _9454 ^ _46051;
  wire _46053 = uncoded_block[1047] ^ uncoded_block[1062];
  wire _46054 = _46053 ^ _12217;
  wire _46055 = _46052 ^ _46054;
  wire _46056 = _46050 ^ _46055;
  wire _46057 = _46045 ^ _46056;
  wire _46058 = _46033 ^ _46057;
  wire _46059 = uncoded_block[1076] ^ uncoded_block[1082];
  wire _46060 = uncoded_block[1087] ^ uncoded_block[1097];
  wire _46061 = _46059 ^ _46060;
  wire _46062 = uncoded_block[1098] ^ uncoded_block[1102];
  wire _46063 = uncoded_block[1106] ^ uncoded_block[1109];
  wire _46064 = _46062 ^ _46063;
  wire _46065 = _46061 ^ _46064;
  wire _46066 = uncoded_block[1117] ^ uncoded_block[1120];
  wire _46067 = _10585 ^ _46066;
  wire _46068 = _5178 ^ _14887;
  wire _46069 = _46067 ^ _46068;
  wire _46070 = _46065 ^ _46069;
  wire _46071 = uncoded_block[1136] ^ uncoded_block[1149];
  wire _46072 = uncoded_block[1153] ^ uncoded_block[1163];
  wire _46073 = _46071 ^ _46072;
  wire _46074 = uncoded_block[1165] ^ uncoded_block[1170];
  wire _46075 = uncoded_block[1172] ^ uncoded_block[1184];
  wire _46076 = _46074 ^ _46075;
  wire _46077 = _46073 ^ _46076;
  wire _46078 = uncoded_block[1198] ^ uncoded_block[1203];
  wire _46079 = _13346 ^ _46078;
  wire _46080 = _608 ^ _1436;
  wire _46081 = _46079 ^ _46080;
  wire _46082 = _46077 ^ _46081;
  wire _46083 = _46070 ^ _46082;
  wire _46084 = uncoded_block[1231] ^ uncoded_block[1236];
  wire _46085 = _46084 ^ _23550;
  wire _46086 = _2232 ^ _11739;
  wire _46087 = _46085 ^ _46086;
  wire _46088 = uncoded_block[1259] ^ uncoded_block[1275];
  wire _46089 = uncoded_block[1282] ^ uncoded_block[1295];
  wire _46090 = _46088 ^ _46089;
  wire _46091 = uncoded_block[1300] ^ uncoded_block[1305];
  wire _46092 = _46091 ^ _14430;
  wire _46093 = _46090 ^ _46092;
  wire _46094 = _46087 ^ _46093;
  wire _46095 = _13395 ^ _657;
  wire _46096 = uncoded_block[1342] ^ uncoded_block[1347];
  wire _46097 = _46096 ^ _10097;
  wire _46098 = _46095 ^ _46097;
  wire _46099 = _2284 ^ _10668;
  wire _46100 = _15966 ^ _11781;
  wire _46101 = _46099 ^ _46100;
  wire _46102 = _46098 ^ _46101;
  wire _46103 = _46094 ^ _46102;
  wire _46104 = _46083 ^ _46103;
  wire _46105 = _46058 ^ _46104;
  wire _46106 = _46014 ^ _46105;
  wire _46107 = uncoded_block[1399] ^ uncoded_block[1405];
  wire _46108 = _46107 ^ _8436;
  wire _46109 = uncoded_block[1418] ^ uncoded_block[1425];
  wire _46110 = _10681 ^ _46109;
  wire _46111 = _46108 ^ _46110;
  wire _46112 = _9025 ^ _14469;
  wire _46113 = _3084 ^ _23176;
  wire _46114 = _46112 ^ _46113;
  wire _46115 = _46111 ^ _46114;
  wire _46116 = uncoded_block[1478] ^ uncoded_block[1485];
  wire _46117 = _1555 ^ _46116;
  wire _46118 = uncoded_block[1494] ^ uncoded_block[1501];
  wire _46119 = _5990 ^ _46118;
  wire _46120 = _46117 ^ _46119;
  wire _46121 = uncoded_block[1510] ^ uncoded_block[1515];
  wire _46122 = _46121 ^ _5343;
  wire _46123 = uncoded_block[1538] ^ uncoded_block[1547];
  wire _46124 = _46123 ^ _15026;
  wire _46125 = _46122 ^ _46124;
  wire _46126 = _46120 ^ _46125;
  wire _46127 = _46115 ^ _46126;
  wire _46128 = uncoded_block[1582] ^ uncoded_block[1589];
  wire _46129 = _13478 ^ _46128;
  wire _46130 = uncoded_block[1595] ^ uncoded_block[1604];
  wire _46131 = uncoded_block[1605] ^ uncoded_block[1611];
  wire _46132 = _46130 ^ _46131;
  wire _46133 = _46129 ^ _46132;
  wire _46134 = _6684 ^ _19931;
  wire _46135 = _17529 ^ _3174;
  wire _46136 = _46134 ^ _46135;
  wire _46137 = _46133 ^ _46136;
  wire _46138 = uncoded_block[1678] ^ uncoded_block[1688];
  wire _46139 = _2422 ^ _46138;
  wire _46140 = _31335 ^ _46139;
  wire _46141 = uncoded_block[1695] ^ uncoded_block[1709];
  wire _46142 = _42191 ^ _46141;
  wire _46143 = _46142 ^ uncoded_block[1712];
  wire _46144 = _46140 ^ _46143;
  wire _46145 = _46137 ^ _46144;
  wire _46146 = _46127 ^ _46145;
  wire _46147 = _46106 ^ _46146;
  wire _46148 = _1683 ^ _3212;
  wire _46149 = _46148 ^ _10789;
  wire _46150 = uncoded_block[14] ^ uncoded_block[18];
  wire _46151 = _46150 ^ _19963;
  wire _46152 = _11344 ^ _15;
  wire _46153 = _46151 ^ _46152;
  wire _46154 = _46149 ^ _46153;
  wire _46155 = _16 ^ _10796;
  wire _46156 = _20457 ^ _886;
  wire _46157 = _46155 ^ _46156;
  wire _46158 = _10238 ^ _11355;
  wire _46159 = uncoded_block[70] ^ uncoded_block[77];
  wire _46160 = _9705 ^ _46159;
  wire _46161 = _46158 ^ _46160;
  wire _46162 = _46157 ^ _46161;
  wire _46163 = _46154 ^ _46162;
  wire _46164 = _11363 ^ _41;
  wire _46165 = _4025 ^ _9713;
  wire _46166 = _46164 ^ _46165;
  wire _46167 = _6758 ^ _12447;
  wire _46168 = _1721 ^ _20957;
  wire _46169 = _46167 ^ _46168;
  wire _46170 = _46166 ^ _46169;
  wire _46171 = uncoded_block[114] ^ uncoded_block[120];
  wire _46172 = _46171 ^ _13017;
  wire _46173 = uncoded_block[133] ^ uncoded_block[136];
  wire _46174 = _4042 ^ _46173;
  wire _46175 = _46172 ^ _46174;
  wire _46176 = _6136 ^ _33909;
  wire _46177 = _4764 ^ _1749;
  wire _46178 = _46176 ^ _46177;
  wire _46179 = _46175 ^ _46178;
  wire _46180 = _46170 ^ _46179;
  wire _46181 = _46163 ^ _46180;
  wire _46182 = uncoded_block[165] ^ uncoded_block[170];
  wire _46183 = _46182 ^ _2521;
  wire _46184 = _46183 ^ _34715;
  wire _46185 = _3284 ^ _16116;
  wire _46186 = _4063 ^ _46185;
  wire _46187 = _46184 ^ _46186;
  wire _46188 = _10849 ^ _10278;
  wire _46189 = uncoded_block[209] ^ uncoded_block[215];
  wire _46190 = _1764 ^ _46189;
  wire _46191 = _46188 ^ _46190;
  wire _46192 = _35136 ^ _17118;
  wire _46193 = _46192 ^ _1776;
  wire _46194 = _46191 ^ _46193;
  wire _46195 = _46187 ^ _46194;
  wire _46196 = _6822 ^ _10860;
  wire _46197 = _46196 ^ _32258;
  wire _46198 = _31834 ^ _1786;
  wire _46199 = _120 ^ _7440;
  wire _46200 = _46198 ^ _46199;
  wire _46201 = _46197 ^ _46200;
  wire _46202 = uncoded_block[269] ^ uncoded_block[276];
  wire _46203 = _46202 ^ _7445;
  wire _46204 = _46203 ^ _20529;
  wire _46205 = _135 ^ _17635;
  wire _46206 = _1807 ^ _4824;
  wire _46207 = _46205 ^ _46206;
  wire _46208 = _46204 ^ _46207;
  wire _46209 = _46201 ^ _46208;
  wire _46210 = _46195 ^ _46209;
  wire _46211 = _46181 ^ _46210;
  wire _46212 = _3337 ^ _145;
  wire _46213 = _13618 ^ _46212;
  wire _46214 = _30116 ^ _8642;
  wire _46215 = _46214 ^ _41505;
  wire _46216 = _46213 ^ _46215;
  wire _46217 = _7463 ^ _9242;
  wire _46218 = _35556 ^ _46217;
  wire _46219 = _1021 ^ _8652;
  wire _46220 = _13089 ^ _15686;
  wire _46221 = _46219 ^ _46220;
  wire _46222 = _46218 ^ _46221;
  wire _46223 = _46216 ^ _46222;
  wire _46224 = _40360 ^ _3369;
  wire _46225 = uncoded_block[373] ^ uncoded_block[383];
  wire _46226 = _1838 ^ _46225;
  wire _46227 = _46224 ^ _46226;
  wire _46228 = _19599 ^ _3381;
  wire _46229 = _12005 ^ _180;
  wire _46230 = _46228 ^ _46229;
  wire _46231 = _46227 ^ _46230;
  wire _46232 = _9808 ^ _27747;
  wire _46233 = _19613 ^ _8671;
  wire _46234 = _14163 ^ _6254;
  wire _46235 = _46233 ^ _46234;
  wire _46236 = _46232 ^ _46235;
  wire _46237 = _46231 ^ _46236;
  wire _46238 = _46223 ^ _46237;
  wire _46239 = _1069 ^ _2650;
  wire _46240 = _35578 ^ _46239;
  wire _46241 = _26495 ^ _4181;
  wire _46242 = _11491 ^ _1878;
  wire _46243 = _46241 ^ _46242;
  wire _46244 = _46240 ^ _46243;
  wire _46245 = _8686 ^ _1083;
  wire _46246 = _4895 ^ _8694;
  wire _46247 = _46245 ^ _46246;
  wire _46248 = _24728 ^ _4906;
  wire _46249 = _46247 ^ _46248;
  wire _46250 = _46244 ^ _46249;
  wire _46251 = _14707 ^ _13148;
  wire _46252 = _4208 ^ _3444;
  wire _46253 = _46251 ^ _46252;
  wire _46254 = _6289 ^ _4921;
  wire _46255 = _46254 ^ _15231;
  wire _46256 = _46253 ^ _46255;
  wire _46257 = _6293 ^ _2684;
  wire _46258 = _5628 ^ _1913;
  wire _46259 = _46257 ^ _46258;
  wire _46260 = _4934 ^ _4937;
  wire _46261 = _3465 ^ _39617;
  wire _46262 = _46260 ^ _46261;
  wire _46263 = _46259 ^ _46262;
  wire _46264 = _46256 ^ _46263;
  wire _46265 = _46250 ^ _46264;
  wire _46266 = _46238 ^ _46265;
  wire _46267 = _46211 ^ _46266;
  wire _46268 = _4941 ^ _11526;
  wire _46269 = _46268 ^ _41939;
  wire _46270 = _36835 ^ _3481;
  wire _46271 = _46269 ^ _46270;
  wire _46272 = _4953 ^ _2709;
  wire _46273 = _46272 ^ _37256;
  wire _46274 = _4242 ^ _7564;
  wire _46275 = _15261 ^ _8749;
  wire _46276 = _46274 ^ _46275;
  wire _46277 = _46273 ^ _46276;
  wire _46278 = _46271 ^ _46277;
  wire _46279 = _4249 ^ _16241;
  wire _46280 = _2729 ^ _10425;
  wire _46281 = _46279 ^ _46280;
  wire _46282 = _6341 ^ _40030;
  wire _46283 = _4261 ^ _2742;
  wire _46284 = _46282 ^ _46283;
  wire _46285 = _46281 ^ _46284;
  wire _46286 = _9886 ^ _3519;
  wire _46287 = _32764 ^ _2751;
  wire _46288 = _46286 ^ _46287;
  wire _46289 = _14766 ^ _6361;
  wire _46290 = _15283 ^ _46289;
  wire _46291 = _46288 ^ _46290;
  wire _46292 = _46285 ^ _46291;
  wire _46293 = _46278 ^ _46292;
  wire _46294 = uncoded_block[707] ^ uncoded_block[711];
  wire _46295 = _46294 ^ _3536;
  wire _46296 = uncoded_block[714] ^ uncoded_block[719];
  wire _46297 = uncoded_block[720] ^ uncoded_block[725];
  wire _46298 = _46296 ^ _46297;
  wire _46299 = _46295 ^ _46298;
  wire _46300 = uncoded_block[731] ^ uncoded_block[736];
  wire _46301 = _14774 ^ _46300;
  wire _46302 = _7005 ^ _4289;
  wire _46303 = _46301 ^ _46302;
  wire _46304 = _46299 ^ _46303;
  wire _46305 = _21600 ^ _356;
  wire _46306 = _24331 ^ _4298;
  wire _46307 = _46305 ^ _46306;
  wire _46308 = _5019 ^ _17776;
  wire _46309 = _6382 ^ _7620;
  wire _46310 = _46308 ^ _46309;
  wire _46311 = _46307 ^ _46310;
  wire _46312 = _46304 ^ _46311;
  wire _46313 = _368 ^ _12673;
  wire _46314 = _46313 ^ _5722;
  wire _46315 = _34062 ^ _5041;
  wire _46316 = _2023 ^ _46315;
  wire _46317 = _46314 ^ _46316;
  wire _46318 = _11030 ^ _22525;
  wire _46319 = uncoded_block[824] ^ uncoded_block[836];
  wire _46320 = _397 ^ _46319;
  wire _46321 = _46318 ^ _46320;
  wire _46322 = _2035 ^ _5737;
  wire _46323 = _8808 ^ _1257;
  wire _46324 = _46322 ^ _46323;
  wire _46325 = _46321 ^ _46324;
  wire _46326 = _46317 ^ _46325;
  wire _46327 = _46312 ^ _46326;
  wire _46328 = _46293 ^ _46327;
  wire _46329 = _14814 ^ _2046;
  wire _46330 = _46329 ^ _5067;
  wire _46331 = _9949 ^ _1266;
  wire _46332 = _12150 ^ _11620;
  wire _46333 = _46331 ^ _46332;
  wire _46334 = _46330 ^ _46333;
  wire _46335 = _16815 ^ _11056;
  wire _46336 = _3613 ^ _14827;
  wire _46337 = _46335 ^ _46336;
  wire _46338 = _5083 ^ _5085;
  wire _46339 = _46338 ^ _33680;
  wire _46340 = _46337 ^ _46339;
  wire _46341 = _46334 ^ _46340;
  wire _46342 = _37717 ^ _44215;
  wire _46343 = uncoded_block[922] ^ uncoded_block[929];
  wire _46344 = uncoded_block[933] ^ uncoded_block[941];
  wire _46345 = _46343 ^ _46344;
  wire _46346 = _46345 ^ _24385;
  wire _46347 = _46342 ^ _46346;
  wire _46348 = _5105 ^ _5783;
  wire _46349 = _4383 ^ _46348;
  wire _46350 = _11646 ^ _8847;
  wire _46351 = _13821 ^ _471;
  wire _46352 = _46350 ^ _46351;
  wire _46353 = _46349 ^ _46352;
  wire _46354 = _46347 ^ _46353;
  wire _46355 = _46341 ^ _46354;
  wire _46356 = _10538 ^ _1319;
  wire _46357 = _40109 ^ _1327;
  wire _46358 = _33277 ^ _46357;
  wire _46359 = _46356 ^ _46358;
  wire _46360 = _1330 ^ _5131;
  wire _46361 = _11663 ^ _8872;
  wire _46362 = _46360 ^ _46361;
  wire _46363 = _27496 ^ _3678;
  wire _46364 = uncoded_block[1045] ^ uncoded_block[1049];
  wire _46365 = _2130 ^ _46364;
  wire _46366 = _46363 ^ _46365;
  wire _46367 = _46362 ^ _46366;
  wire _46368 = _46359 ^ _46367;
  wire _46369 = _13847 ^ _34932;
  wire _46370 = _8888 ^ _3689;
  wire _46371 = _21685 ^ _2147;
  wire _46372 = _46370 ^ _46371;
  wire _46373 = _46369 ^ _46372;
  wire _46374 = uncoded_block[1080] ^ uncoded_block[1085];
  wire _46375 = _46374 ^ _3696;
  wire _46376 = _46375 ^ _23070;
  wire _46377 = _5166 ^ _5169;
  wire _46378 = _8910 ^ _20761;
  wire _46379 = _46377 ^ _46378;
  wire _46380 = _46376 ^ _46379;
  wire _46381 = _46373 ^ _46380;
  wire _46382 = _46368 ^ _46381;
  wire _46383 = _46355 ^ _46382;
  wire _46384 = _46328 ^ _46383;
  wire _46385 = _46267 ^ _46384;
  wire _46386 = uncoded_block[1125] ^ uncoded_block[1134];
  wire _46387 = _46386 ^ _9496;
  wire _46388 = _23980 ^ _46387;
  wire _46389 = uncoded_block[1145] ^ uncoded_block[1149];
  wire _46390 = _46389 ^ _4468;
  wire _46391 = uncoded_block[1154] ^ uncoded_block[1157];
  wire _46392 = _46391 ^ _3733;
  wire _46393 = _46390 ^ _46392;
  wire _46394 = _46388 ^ _46393;
  wire _46395 = _22627 ^ _13335;
  wire _46396 = _9506 ^ _585;
  wire _46397 = _46395 ^ _46396;
  wire _46398 = _2193 ^ _592;
  wire _46399 = _2196 ^ _10612;
  wire _46400 = _46398 ^ _46399;
  wire _46401 = _46397 ^ _46400;
  wire _46402 = _46394 ^ _46401;
  wire _46403 = _14398 ^ _17400;
  wire _46404 = _16399 ^ _1427;
  wire _46405 = _46403 ^ _46404;
  wire _46406 = _3765 ^ _6532;
  wire _46407 = _21720 ^ _46406;
  wire _46408 = _46405 ^ _46407;
  wire _46409 = _12819 ^ _1439;
  wire _46410 = _31228 ^ _7774;
  wire _46411 = _46409 ^ _46410;
  wire _46412 = _4509 ^ _11734;
  wire _46413 = _46412 ^ _13367;
  wire _46414 = _46411 ^ _46413;
  wire _46415 = _46408 ^ _46414;
  wire _46416 = _46402 ^ _46415;
  wire _46417 = _3784 ^ _627;
  wire _46418 = _35373 ^ _46417;
  wire _46419 = uncoded_block[1267] ^ uncoded_block[1271];
  wire _46420 = _46419 ^ _1463;
  wire _46421 = _7183 ^ _16924;
  wire _46422 = _46420 ^ _46421;
  wire _46423 = _46418 ^ _46422;
  wire _46424 = _18866 ^ _1469;
  wire _46425 = _46424 ^ _23130;
  wire _46426 = _16431 ^ _7802;
  wire _46427 = _14430 ^ _21293;
  wire _46428 = _46426 ^ _46427;
  wire _46429 = _46425 ^ _46428;
  wire _46430 = _46423 ^ _46429;
  wire _46431 = _19848 ^ _28672;
  wire _46432 = _3034 ^ _14440;
  wire _46433 = uncoded_block[1343] ^ uncoded_block[1347];
  wire _46434 = _46433 ^ _3041;
  wire _46435 = _46432 ^ _46434;
  wire _46436 = _46431 ^ _46435;
  wire _46437 = _10097 ^ _6588;
  wire _46438 = _25393 ^ _2283;
  wire _46439 = _46437 ^ _46438;
  wire _46440 = _29939 ^ _10108;
  wire _46441 = _36195 ^ _46440;
  wire _46442 = _46439 ^ _46441;
  wire _46443 = _46436 ^ _46442;
  wire _46444 = _46430 ^ _46443;
  wire _46445 = _46416 ^ _46444;
  wire _46446 = _11782 ^ _2293;
  wire _46447 = _694 ^ _13938;
  wire _46448 = _46446 ^ _46447;
  wire _46449 = _29090 ^ _3846;
  wire _46450 = _18452 ^ _702;
  wire _46451 = _46449 ^ _46450;
  wire _46452 = _46448 ^ _46451;
  wire _46453 = _7843 ^ _3082;
  wire _46454 = _4590 ^ _2322;
  wire _46455 = _37038 ^ _46454;
  wire _46456 = _46453 ^ _46455;
  wire _46457 = _46452 ^ _46456;
  wire _46458 = _3865 ^ _16474;
  wire _46459 = _46458 ^ _23612;
  wire _46460 = _10136 ^ _40603;
  wire _46461 = _13963 ^ _19887;
  wire _46462 = _46460 ^ _46461;
  wire _46463 = _46459 ^ _46462;
  wire _46464 = _2349 ^ _15996;
  wire _46465 = _46464 ^ _15512;
  wire _46466 = _747 ^ _3894;
  wire _46467 = _4616 ^ _8467;
  wire _46468 = _46466 ^ _46467;
  wire _46469 = _46465 ^ _46468;
  wire _46470 = _46463 ^ _46469;
  wire _46471 = _46457 ^ _46470;
  wire _46472 = _7265 ^ _15004;
  wire _46473 = _46472 ^ _29122;
  wire _46474 = uncoded_block[1536] ^ uncoded_block[1541];
  wire _46475 = _6005 ^ _46474;
  wire _46476 = _23198 ^ _46475;
  wire _46477 = _46473 ^ _46476;
  wire _46478 = _13472 ^ _22731;
  wire _46479 = _13988 ^ _46478;
  wire _46480 = _4638 ^ _7889;
  wire _46481 = _24102 ^ _30870;
  wire _46482 = _46480 ^ _46481;
  wire _46483 = _46479 ^ _46482;
  wire _46484 = _46477 ^ _46483;
  wire _46485 = uncoded_block[1574] ^ uncoded_block[1578];
  wire _46486 = _46485 ^ _1609;
  wire _46487 = uncoded_block[1582] ^ uncoded_block[1586];
  wire _46488 = _46487 ^ _20401;
  wire _46489 = _46486 ^ _46488;
  wire _46490 = _2394 ^ _13486;
  wire _46491 = _5373 ^ _3153;
  wire _46492 = _46490 ^ _46491;
  wire _46493 = _46489 ^ _46492;
  wire _46494 = _6677 ^ _4662;
  wire _46495 = _12940 ^ _804;
  wire _46496 = _46494 ^ _46495;
  wire _46497 = uncoded_block[1625] ^ uncoded_block[1630];
  wire _46498 = _805 ^ _46497;
  wire _46499 = _19929 ^ _7308;
  wire _46500 = _46498 ^ _46499;
  wire _46501 = _46496 ^ _46500;
  wire _46502 = _46493 ^ _46501;
  wire _46503 = _46484 ^ _46502;
  wire _46504 = _46471 ^ _46503;
  wire _46505 = _46445 ^ _46504;
  wire _46506 = _7309 ^ _7921;
  wire _46507 = _46506 ^ _18031;
  wire _46508 = uncoded_block[1666] ^ uncoded_block[1671];
  wire _46509 = _12960 ^ _46508;
  wire _46510 = _39076 ^ _46509;
  wire _46511 = _46507 ^ _46510;
  wire _46512 = _31339 ^ _35081;
  wire _46513 = _46512 ^ _3191;
  wire _46514 = _6066 ^ _29162;
  wire _46515 = _6068 ^ _15063;
  wire _46516 = _46514 ^ _46515;
  wire _46517 = _46513 ^ _46516;
  wire _46518 = _46511 ^ _46517;
  wire _46519 = _7335 ^ _854;
  wire _46520 = _46519 ^ _21402;
  wire _46521 = _46518 ^ _46520;
  wire _46522 = _46505 ^ _46521;
  wire _46523 = _46385 ^ _46522;
  wire _46524 = _32201 ^ _6724;
  wire _46525 = _3211 ^ _46524;
  wire _46526 = _3213 ^ _4713;
  wire _46527 = _868 ^ _7351;
  wire _46528 = _46526 ^ _46527;
  wire _46529 = _46525 ^ _46528;
  wire _46530 = _37113 ^ _15589;
  wire _46531 = _19501 ^ _2466;
  wire _46532 = _882 ^ _8554;
  wire _46533 = _46531 ^ _46532;
  wire _46534 = _46530 ^ _46533;
  wire _46535 = _46529 ^ _46534;
  wire _46536 = _888 ^ _20465;
  wire _46537 = _14050 ^ _46536;
  wire _46538 = _35 ^ _10244;
  wire _46539 = _44427 ^ _46538;
  wire _46540 = _46537 ^ _46539;
  wire _46541 = uncoded_block[79] ^ uncoded_block[87];
  wire _46542 = _901 ^ _46541;
  wire _46543 = _903 ^ _20952;
  wire _46544 = _46542 ^ _46543;
  wire _46545 = _3249 ^ _15097;
  wire _46546 = uncoded_block[106] ^ uncoded_block[110];
  wire _46547 = _19025 ^ _46546;
  wire _46548 = _46545 ^ _46547;
  wire _46549 = _46544 ^ _46548;
  wire _46550 = _46540 ^ _46549;
  wire _46551 = _46535 ^ _46550;
  wire _46552 = _18090 ^ _12451;
  wire _46553 = _10817 ^ _46552;
  wire _46554 = uncoded_block[132] ^ uncoded_block[135];
  wire _46555 = _46554 ^ _2510;
  wire _46556 = _17589 ^ _46555;
  wire _46557 = _46553 ^ _46556;
  wire _46558 = _24178 ^ _15622;
  wire _46559 = _31391 ^ _46558;
  wire _46560 = _74 ^ _16604;
  wire _46561 = _36325 ^ _46560;
  wire _46562 = _46559 ^ _46561;
  wire _46563 = _46557 ^ _46562;
  wire _46564 = _5473 ^ _2521;
  wire _46565 = _20979 ^ _4770;
  wire _46566 = _46564 ^ _46565;
  wire _46567 = _6798 ^ _32248;
  wire _46568 = _31404 ^ _46567;
  wire _46569 = _46566 ^ _46568;
  wire _46570 = _6806 ^ _959;
  wire _46571 = _46570 ^ _30086;
  wire _46572 = uncoded_block[232] ^ uncoded_block[240];
  wire _46573 = _4080 ^ _46572;
  wire _46574 = _6172 ^ _1781;
  wire _46575 = _46573 ^ _46574;
  wire _46576 = _46571 ^ _46575;
  wire _46577 = _46569 ^ _46576;
  wire _46578 = _46563 ^ _46577;
  wire _46579 = _46551 ^ _46578;
  wire _46580 = uncoded_block[250] ^ uncoded_block[256];
  wire _46581 = _7432 ^ _46580;
  wire _46582 = _8041 ^ _6185;
  wire _46583 = _46581 ^ _46582;
  wire _46584 = _6188 ^ _14642;
  wire _46585 = _4102 ^ _5512;
  wire _46586 = _46584 ^ _46585;
  wire _46587 = _46583 ^ _46586;
  wire _46588 = _4103 ^ _988;
  wire _46589 = _46588 ^ _23757;
  wire _46590 = uncoded_block[295] ^ uncoded_block[303];
  wire _46591 = _994 ^ _46590;
  wire _46592 = _25569 ^ _15168;
  wire _46593 = _46591 ^ _46592;
  wire _46594 = _46589 ^ _46593;
  wire _46595 = _46587 ^ _46594;
  wire _46596 = _44856 ^ _18617;
  wire _46597 = uncoded_block[336] ^ uncoded_block[341];
  wire _46598 = _3352 ^ _46597;
  wire _46599 = _46596 ^ _46598;
  wire _46600 = _159 ^ _3359;
  wire _46601 = _46600 ^ _14666;
  wire _46602 = _46599 ^ _46601;
  wire _46603 = _1029 ^ _21030;
  wire _46604 = _8655 ^ _6232;
  wire _46605 = _46603 ^ _46604;
  wire _46606 = _7474 ^ _6235;
  wire _46607 = uncoded_block[383] ^ uncoded_block[386];
  wire _46608 = _46607 ^ _21504;
  wire _46609 = _46606 ^ _46608;
  wire _46610 = _46605 ^ _46609;
  wire _46611 = _46602 ^ _46610;
  wire _46612 = _46595 ^ _46611;
  wire _46613 = _1847 ^ _1849;
  wire _46614 = _46613 ^ _12546;
  wire _46615 = _15197 ^ _35576;
  wire _46616 = _21509 ^ _46615;
  wire _46617 = _46614 ^ _46616;
  wire _46618 = _14689 ^ _25601;
  wire _46619 = _46618 ^ _36389;
  wire _46620 = uncoded_block[446] ^ uncoded_block[450];
  wire _46621 = _46620 ^ _12562;
  wire _46622 = uncoded_block[458] ^ uncoded_block[463];
  wire _46623 = _6261 ^ _46622;
  wire _46624 = _46621 ^ _46623;
  wire _46625 = _46619 ^ _46624;
  wire _46626 = _46617 ^ _46625;
  wire _46627 = _4890 ^ _23357;
  wire _46628 = _26944 ^ _12025;
  wire _46629 = _46627 ^ _46628;
  wire _46630 = _7515 ^ _4903;
  wire _46631 = _21062 ^ _46630;
  wire _46632 = _46629 ^ _46631;
  wire _46633 = _4905 ^ _8120;
  wire _46634 = _13674 ^ _17694;
  wire _46635 = _46633 ^ _46634;
  wire _46636 = _232 ^ _9841;
  wire _46637 = _46636 ^ _9849;
  wire _46638 = _46635 ^ _46637;
  wire _46639 = _46632 ^ _46638;
  wire _46640 = _46626 ^ _46639;
  wire _46641 = _46612 ^ _46640;
  wire _46642 = _46579 ^ _46641;
  wire _46643 = uncoded_block[537] ^ uncoded_block[544];
  wire _46644 = _5617 ^ _46643;
  wire _46645 = _13686 ^ _46644;
  wire _46646 = _1909 ^ _6300;
  wire _46647 = _20107 ^ _1916;
  wire _46648 = _46646 ^ _46647;
  wire _46649 = _46645 ^ _46648;
  wire _46650 = _3461 ^ _3464;
  wire _46651 = _46650 ^ _16722;
  wire _46652 = _17221 ^ _28136;
  wire _46653 = _6947 ^ _28891;
  wire _46654 = _46652 ^ _46653;
  wire _46655 = _46651 ^ _46654;
  wire _46656 = _46649 ^ _46655;
  wire _46657 = uncoded_block[595] ^ uncoded_block[601];
  wire _46658 = _2700 ^ _46657;
  wire _46659 = _46658 ^ _9335;
  wire _46660 = _41570 ^ _16238;
  wire _46661 = _1946 ^ _12618;
  wire _46662 = _46660 ^ _46661;
  wire _46663 = _46659 ^ _46662;
  wire _46664 = _6966 ^ _289;
  wire _46665 = _46664 ^ _25203;
  wire _46666 = _9343 ^ _4972;
  wire _46667 = _46666 ^ _39633;
  wire _46668 = _46665 ^ _46667;
  wire _46669 = _46663 ^ _46668;
  wire _46670 = _46656 ^ _46669;
  wire _46671 = _3508 ^ _3513;
  wire _46672 = _46671 ^ _16750;
  wire _46673 = _1173 ^ _311;
  wire _46674 = _46673 ^ _11553;
  wire _46675 = _46672 ^ _46674;
  wire _46676 = _1968 ^ _6353;
  wire _46677 = _26557 ^ _32767;
  wire _46678 = _46676 ^ _46677;
  wire _46679 = uncoded_block[705] ^ uncoded_block[711];
  wire _46680 = _17258 ^ _46679;
  wire _46681 = _22969 ^ _46680;
  wire _46682 = _46678 ^ _46681;
  wire _46683 = _46675 ^ _46682;
  wire _46684 = _337 ^ _6367;
  wire _46685 = _46684 ^ _28548;
  wire _46686 = _7001 ^ _46300;
  wire _46687 = _46686 ^ _3551;
  wire _46688 = _46685 ^ _46687;
  wire _46689 = _5012 ^ _30232;
  wire _46690 = _4298 ^ _360;
  wire _46691 = _46689 ^ _46690;
  wire _46692 = _5020 ^ _12113;
  wire _46693 = _12114 ^ _3562;
  wire _46694 = _46692 ^ _46693;
  wire _46695 = _46691 ^ _46694;
  wire _46696 = _46688 ^ _46695;
  wire _46697 = _46683 ^ _46696;
  wire _46698 = _46670 ^ _46697;
  wire _46699 = _8790 ^ _3574;
  wire _46700 = _40454 ^ _46699;
  wire _46701 = _2021 ^ _2801;
  wire _46702 = _46701 ^ _33228;
  wire _46703 = _46700 ^ _46702;
  wire _46704 = _4324 ^ _27843;
  wire _46705 = _3587 ^ _12135;
  wire _46706 = _46704 ^ _46705;
  wire _46707 = _10490 ^ _16801;
  wire _46708 = _46707 ^ _19722;
  wire _46709 = _46706 ^ _46708;
  wire _46710 = _46703 ^ _46709;
  wire _46711 = uncoded_block[847] ^ uncoded_block[855];
  wire _46712 = _8808 ^ _46711;
  wire _46713 = uncoded_block[859] ^ uncoded_block[864];
  wire _46714 = _8812 ^ _46713;
  wire _46715 = _46712 ^ _46714;
  wire _46716 = _27452 ^ _12150;
  wire _46717 = _46716 ^ _26612;
  wire _46718 = _46715 ^ _46717;
  wire _46719 = _5078 ^ _2838;
  wire _46720 = _2058 ^ _12704;
  wire _46721 = _46719 ^ _46720;
  wire _46722 = _14829 ^ _11062;
  wire _46723 = uncoded_block[909] ^ uncoded_block[914];
  wire _46724 = _1284 ^ _46723;
  wire _46725 = _46722 ^ _46724;
  wire _46726 = _46721 ^ _46725;
  wire _46727 = _46718 ^ _46726;
  wire _46728 = _46710 ^ _46727;
  wire _46729 = _3631 ^ _31995;
  wire _46730 = _3630 ^ _46729;
  wire _46731 = _2857 ^ _5773;
  wire _46732 = _452 ^ _22105;
  wire _46733 = _46731 ^ _46732;
  wire _46734 = _46730 ^ _46733;
  wire _46735 = _1303 ^ _1307;
  wire _46736 = _43070 ^ _46735;
  wire _46737 = _7680 ^ _11646;
  wire _46738 = _2093 ^ _468;
  wire _46739 = _46737 ^ _46738;
  wire _46740 = _46736 ^ _46739;
  wire _46741 = _46734 ^ _46740;
  wire _46742 = uncoded_block[977] ^ uncoded_block[983];
  wire _46743 = _46742 ^ _2102;
  wire _46744 = _16338 ^ _3663;
  wire _46745 = _46743 ^ _46744;
  wire _46746 = _25292 ^ _488;
  wire _46747 = _46745 ^ _46746;
  wire _46748 = uncoded_block[1012] ^ uncoded_block[1016];
  wire _46749 = _46748 ^ _494;
  wire _46750 = _12752 ^ _4417;
  wire _46751 = _46749 ^ _46750;
  wire _46752 = _34925 ^ _2129;
  wire _46753 = _6475 ^ _38937;
  wire _46754 = _46752 ^ _46753;
  wire _46755 = _46751 ^ _46754;
  wire _46756 = _46747 ^ _46755;
  wire _46757 = _46741 ^ _46756;
  wire _46758 = _46728 ^ _46757;
  wire _46759 = _46698 ^ _46758;
  wire _46760 = _46642 ^ _46759;
  wire _46761 = _15870 ^ _32856;
  wire _46762 = _519 ^ _2916;
  wire _46763 = _522 ^ _15395;
  wire _46764 = _46762 ^ _46763;
  wire _46765 = _46761 ^ _46764;
  wire _46766 = _11122 ^ _2146;
  wire _46767 = _8895 ^ _8904;
  wire _46768 = _46766 ^ _46767;
  wire _46769 = _22149 ^ _11137;
  wire _46770 = uncoded_block[1096] ^ uncoded_block[1100];
  wire _46771 = _46770 ^ _14372;
  wire _46772 = _46769 ^ _46771;
  wire _46773 = _46768 ^ _46772;
  wire _46774 = _46765 ^ _46773;
  wire _46775 = _2941 ^ _14376;
  wire _46776 = _36958 ^ _46775;
  wire _46777 = _14380 ^ _41288;
  wire _46778 = _25789 ^ _46777;
  wire _46779 = _46776 ^ _46778;
  wire _46780 = uncoded_block[1144] ^ uncoded_block[1151];
  wire _46781 = _46780 ^ _3727;
  wire _46782 = _29878 ^ _3734;
  wire _46783 = _46781 ^ _46782;
  wire _46784 = _3739 ^ _5872;
  wire _46785 = _40540 ^ _46784;
  wire _46786 = _46783 ^ _46785;
  wire _46787 = _46779 ^ _46786;
  wire _46788 = _46774 ^ _46787;
  wire _46789 = _27539 ^ _35354;
  wire _46790 = _2200 ^ _6525;
  wire _46791 = _46789 ^ _46790;
  wire _46792 = _597 ^ _2206;
  wire _46793 = _7163 ^ _2210;
  wire _46794 = _46792 ^ _46793;
  wire _46795 = _46791 ^ _46794;
  wire _46796 = _2216 ^ _7765;
  wire _46797 = _46796 ^ _24914;
  wire _46798 = _5891 ^ _1439;
  wire _46799 = _21722 ^ _46798;
  wire _46800 = _46797 ^ _46799;
  wire _46801 = _46795 ^ _46800;
  wire _46802 = uncoded_block[1237] ^ uncoded_block[1245];
  wire _46803 = uncoded_block[1251] ^ uncoded_block[1257];
  wire _46804 = _46802 ^ _46803;
  wire _46805 = _32492 ^ _46804;
  wire _46806 = _3786 ^ _12832;
  wire _46807 = _21734 ^ _46806;
  wire _46808 = _46805 ^ _46807;
  wire _46809 = _35377 ^ _13379;
  wire _46810 = _13380 ^ _30797;
  wire _46811 = _3015 ^ _17927;
  wire _46812 = _46810 ^ _46811;
  wire _46813 = _46809 ^ _46812;
  wire _46814 = _46808 ^ _46813;
  wire _46815 = _46801 ^ _46814;
  wire _46816 = _46788 ^ _46815;
  wire _46817 = _3808 ^ _2261;
  wire _46818 = _4538 ^ _46817;
  wire _46819 = uncoded_block[1319] ^ uncoded_block[1324];
  wire _46820 = _21293 ^ _46819;
  wire _46821 = _656 ^ _1494;
  wire _46822 = _46820 ^ _46821;
  wire _46823 = _46818 ^ _46822;
  wire _46824 = _26736 ^ _45065;
  wire _46825 = _32515 ^ _46824;
  wire _46826 = uncoded_block[1363] ^ uncoded_block[1374];
  wire _46827 = _46826 ^ _12305;
  wire _46828 = _7219 ^ _12307;
  wire _46829 = _46827 ^ _46828;
  wire _46830 = _46825 ^ _46829;
  wire _46831 = _46823 ^ _46830;
  wire _46832 = uncoded_block[1391] ^ uncoded_block[1399];
  wire _46833 = _5950 ^ _46832;
  wire _46834 = _4578 ^ _9585;
  wire _46835 = _46833 ^ _46834;
  wire _46836 = _13947 ^ _17461;
  wire _46837 = _704 ^ _11792;
  wire _46838 = _46836 ^ _46837;
  wire _46839 = _46835 ^ _46838;
  wire _46840 = uncoded_block[1436] ^ uncoded_block[1441];
  wire _46841 = _23604 ^ _46840;
  wire _46842 = _25861 ^ _46841;
  wire _46843 = _1541 ^ _9033;
  wire _46844 = _46843 ^ _35806;
  wire _46845 = _46842 ^ _46844;
  wire _46846 = _46839 ^ _46845;
  wire _46847 = _46831 ^ _46846;
  wire _46848 = _37044 ^ _38225;
  wire _46849 = uncoded_block[1473] ^ uncoded_block[1479];
  wire _46850 = _5983 ^ _46849;
  wire _46851 = _23181 ^ _11809;
  wire _46852 = _46850 ^ _46851;
  wire _46853 = _46848 ^ _46852;
  wire _46854 = _12896 ^ _19890;
  wire _46855 = _46854 ^ _28370;
  wire _46856 = _5337 ^ _754;
  wire _46857 = _29971 ^ _46856;
  wire _46858 = _46855 ^ _46857;
  wire _46859 = _46853 ^ _46858;
  wire _46860 = uncoded_block[1521] ^ uncoded_block[1525];
  wire _46861 = _46860 ^ _1582;
  wire _46862 = uncoded_block[1531] ^ uncoded_block[1535];
  wire _46863 = _46862 ^ _15009;
  wire _46864 = _46861 ^ _46863;
  wire _46865 = _6008 ^ _13471;
  wire _46866 = _14496 ^ _9070;
  wire _46867 = _46865 ^ _46866;
  wire _46868 = _46864 ^ _46867;
  wire _46869 = _1596 ^ _4640;
  wire _46870 = _46869 ^ _20393;
  wire _46871 = _7285 ^ _4647;
  wire _46872 = _6663 ^ _21821;
  wire _46873 = _46871 ^ _46872;
  wire _46874 = _46870 ^ _46873;
  wire _46875 = _46868 ^ _46874;
  wire _46876 = _46859 ^ _46875;
  wire _46877 = _46847 ^ _46876;
  wire _46878 = _46816 ^ _46877;
  wire _46879 = uncoded_block[1586] ^ uncoded_block[1594];
  wire _46880 = _46879 ^ _3934;
  wire _46881 = _3151 ^ _26343;
  wire _46882 = _46880 ^ _46881;
  wire _46883 = _31740 ^ _7908;
  wire _46884 = _29997 ^ _25906;
  wire _46885 = _46883 ^ _46884;
  wire _46886 = _46882 ^ _46885;
  wire _46887 = _35064 ^ _23658;
  wire _46888 = _10754 ^ _20901;
  wire _46889 = _46887 ^ _46888;
  wire _46890 = _42179 ^ _41405;
  wire _46891 = _46889 ^ _46890;
  wire _46892 = _46886 ^ _46891;
  wire _46893 = _14011 ^ _822;
  wire _46894 = _2419 ^ _3180;
  wire _46895 = _46893 ^ _46894;
  wire _46896 = _19471 ^ _830;
  wire _46897 = _7325 ^ _17040;
  wire _46898 = _46896 ^ _46897;
  wire _46899 = _46895 ^ _46898;
  wire _46900 = _34660 ^ _41420;
  wire _46901 = _1669 ^ _9120;
  wire _46902 = _22314 ^ _848;
  wire _46903 = _46901 ^ _46902;
  wire _46904 = _46900 ^ _46903;
  wire _46905 = _46899 ^ _46904;
  wire _46906 = _46892 ^ _46905;
  wire _46907 = _10778 ^ _3200;
  wire _46908 = _20923 ^ uncoded_block[1722];
  wire _46909 = _46907 ^ _46908;
  wire _46910 = _46906 ^ _46909;
  wire _46911 = _46878 ^ _46910;
  wire _46912 = _46760 ^ _46911;
  wire _46913 = uncoded_block[6] ^ uncoded_block[9];
  wire _46914 = _4710 ^ _46913;
  wire _46915 = _17058 ^ _3998;
  wire _46916 = _46914 ^ _46915;
  wire _46917 = _1693 ^ _6732;
  wire _46918 = _42206 ^ _46917;
  wire _46919 = _46916 ^ _46918;
  wire _46920 = _15594 ^ _3232;
  wire _46921 = _37915 ^ _46920;
  wire _46922 = _25 ^ _7364;
  wire _46923 = _46922 ^ _14581;
  wire _46924 = _46921 ^ _46923;
  wire _46925 = _46919 ^ _46924;
  wire _46926 = _26393 ^ _1712;
  wire _46927 = _2481 ^ _6750;
  wire _46928 = _46926 ^ _46927;
  wire _46929 = _15603 ^ _4026;
  wire _46930 = _43273 ^ _46929;
  wire _46931 = _46928 ^ _46930;
  wire _46932 = _14068 ^ _4028;
  wire _46933 = _46932 ^ _20477;
  wire _46934 = _15103 ^ _18090;
  wire _46935 = _12451 ^ _2502;
  wire _46936 = _46934 ^ _46935;
  wire _46937 = _46933 ^ _46936;
  wire _46938 = _46931 ^ _46937;
  wire _46939 = _46925 ^ _46938;
  wire _46940 = _3262 ^ _4042;
  wire _46941 = _22819 ^ _11918;
  wire _46942 = _46940 ^ _46941;
  wire _46943 = uncoded_block[144] ^ uncoded_block[150];
  wire _46944 = _15114 ^ _46943;
  wire _46945 = uncoded_block[154] ^ uncoded_block[157];
  wire _46946 = _46945 ^ _21906;
  wire _46947 = _46944 ^ _46946;
  wire _46948 = _46942 ^ _46947;
  wire _46949 = _4053 ^ _937;
  wire _46950 = _46949 ^ _31400;
  wire _46951 = _17604 ^ _8012;
  wire _46952 = _46950 ^ _46951;
  wire _46953 = _46948 ^ _46952;
  wire _46954 = _18111 ^ _10277;
  wire _46955 = _4068 ^ _3291;
  wire _46956 = _46954 ^ _46955;
  wire _46957 = _30963 ^ _27295;
  wire _46958 = _14105 ^ _2545;
  wire _46959 = _46957 ^ _46958;
  wire _46960 = _46956 ^ _46959;
  wire _46961 = _15144 ^ _39154;
  wire _46962 = _31411 ^ _46961;
  wire _46963 = uncoded_block[261] ^ uncoded_block[267];
  wire _46964 = _46963 ^ _985;
  wire _46965 = _34736 ^ _46964;
  wire _46966 = _46962 ^ _46965;
  wire _46967 = _46960 ^ _46966;
  wire _46968 = _46953 ^ _46967;
  wire _46969 = _46939 ^ _46968;
  wire _46970 = _14124 ^ _10303;
  wire _46971 = _1796 ^ _11428;
  wire _46972 = _46970 ^ _46971;
  wire _46973 = _14133 ^ _12515;
  wire _46974 = _4109 ^ _46973;
  wire _46975 = _46972 ^ _46974;
  wire _46976 = _22866 ^ _15671;
  wire _46977 = _4830 ^ _4832;
  wire _46978 = _46976 ^ _46977;
  wire _46979 = _21947 ^ _9240;
  wire _46980 = uncoded_block[335] ^ uncoded_block[342];
  wire _46981 = _46980 ^ _3359;
  wire _46982 = _46979 ^ _46981;
  wire _46983 = _46978 ^ _46982;
  wire _46984 = _46975 ^ _46983;
  wire _46985 = _3362 ^ _6228;
  wire _46986 = _14666 ^ _46985;
  wire _46987 = _5548 ^ _1835;
  wire _46988 = _46987 ^ _9796;
  wire _46989 = _46986 ^ _46988;
  wire _46990 = _40363 ^ _26474;
  wire _46991 = _11468 ^ _28478;
  wire _46992 = _46990 ^ _46991;
  wire _46993 = _46989 ^ _46992;
  wire _46994 = _46984 ^ _46993;
  wire _46995 = _2629 ^ _38785;
  wire _46996 = _18175 ^ _4874;
  wire _46997 = _46995 ^ _46996;
  wire _46998 = _9816 ^ _1063;
  wire _46999 = _46998 ^ _4880;
  wire _47000 = _46997 ^ _46999;
  wire _47001 = _21052 ^ _11486;
  wire _47002 = _19621 ^ _5584;
  wire _47003 = _47001 ^ _47002;
  wire _47004 = _1871 ^ _4181;
  wire _47005 = _1874 ^ _4186;
  wire _47006 = _47004 ^ _47005;
  wire _47007 = _47003 ^ _47006;
  wire _47008 = _47000 ^ _47007;
  wire _47009 = _1082 ^ _12025;
  wire _47010 = _12028 ^ _20588;
  wire _47011 = _47009 ^ _47010;
  wire _47012 = _5600 ^ _30167;
  wire _47013 = _6279 ^ _6921;
  wire _47014 = _47012 ^ _47013;
  wire _47015 = _47011 ^ _47014;
  wire _47016 = _12034 ^ _5611;
  wire _47017 = _4908 ^ _10945;
  wire _47018 = _47016 ^ _47017;
  wire _47019 = _4910 ^ _18206;
  wire _47020 = _6289 ^ _4922;
  wire _47021 = _47019 ^ _47020;
  wire _47022 = _47018 ^ _47021;
  wire _47023 = _47015 ^ _47022;
  wire _47024 = _47008 ^ _47023;
  wire _47025 = _46994 ^ _47024;
  wire _47026 = _46969 ^ _47025;
  wire _47027 = _14719 ^ _6298;
  wire _47028 = _36820 ^ _47027;
  wire _47029 = uncoded_block[554] ^ uncoded_block[558];
  wire _47030 = _14725 ^ _47029;
  wire _47031 = uncoded_block[559] ^ uncoded_block[566];
  wire _47032 = _47031 ^ _4223;
  wire _47033 = _47030 ^ _47032;
  wire _47034 = _47028 ^ _47033;
  wire _47035 = _4224 ^ _4941;
  wire _47036 = _47035 ^ _1134;
  wire _47037 = _3478 ^ _15247;
  wire _47038 = _1140 ^ _47037;
  wire _47039 = _47036 ^ _47038;
  wire _47040 = _47034 ^ _47039;
  wire _47041 = _2709 ^ _14218;
  wire _47042 = _13174 ^ _47041;
  wire _47043 = _20121 ^ _7565;
  wire _47044 = _47042 ^ _47043;
  wire _47045 = _1948 ^ _6966;
  wire _47046 = _14744 ^ _47045;
  wire _47047 = _12071 ^ _6330;
  wire _47048 = _47047 ^ _22953;
  wire _47049 = _47046 ^ _47048;
  wire _47050 = _47044 ^ _47049;
  wire _47051 = _47040 ^ _47050;
  wire _47052 = _15766 ^ _28908;
  wire _47053 = _23848 ^ _47052;
  wire _47054 = _304 ^ _2739;
  wire _47055 = _4262 ^ _1173;
  wire _47056 = _47054 ^ _47055;
  wire _47057 = _47053 ^ _47056;
  wire _47058 = uncoded_block[667] ^ uncoded_block[674];
  wire _47059 = _47058 ^ _10434;
  wire _47060 = _1968 ^ _32764;
  wire _47061 = _47059 ^ _47060;
  wire _47062 = _2754 ^ _29756;
  wire _47063 = uncoded_block[701] ^ uncoded_block[707];
  wire _47064 = _11562 ^ _47063;
  wire _47065 = _47062 ^ _47064;
  wire _47066 = _47061 ^ _47065;
  wire _47067 = _47057 ^ _47066;
  wire _47068 = uncoded_block[727] ^ uncoded_block[731];
  wire _47069 = _38450 ^ _47068;
  wire _47070 = _25672 ^ _47069;
  wire _47071 = _41193 ^ _34048;
  wire _47072 = _21600 ^ _5013;
  wire _47073 = _47071 ^ _47072;
  wire _47074 = _47070 ^ _47073;
  wire _47075 = _21139 ^ _2003;
  wire _47076 = _47075 ^ _20162;
  wire _47077 = _3561 ^ _8787;
  wire _47078 = _7021 ^ _5715;
  wire _47079 = _47077 ^ _47078;
  wire _47080 = _47076 ^ _47079;
  wire _47081 = _47074 ^ _47080;
  wire _47082 = _47067 ^ _47081;
  wire _47083 = _47051 ^ _47082;
  wire _47084 = _19218 ^ _1225;
  wire _47085 = _47084 ^ _3575;
  wire _47086 = _382 ^ _4316;
  wire _47087 = _47086 ^ _9395;
  wire _47088 = _47085 ^ _47087;
  wire _47089 = _15814 ^ _5042;
  wire _47090 = _9397 ^ _3584;
  wire _47091 = _47089 ^ _47090;
  wire _47092 = _30673 ^ _45721;
  wire _47093 = _47091 ^ _47092;
  wire _47094 = _47088 ^ _47093;
  wire _47095 = _7043 ^ _5058;
  wire _47096 = _405 ^ _1262;
  wire _47097 = _47095 ^ _47096;
  wire _47098 = _41224 ^ _7653;
  wire _47099 = _47097 ^ _47098;
  wire _47100 = _2831 ^ _7060;
  wire _47101 = _8820 ^ _13797;
  wire _47102 = _47100 ^ _47101;
  wire _47103 = _14827 ^ _4355;
  wire _47104 = _47103 ^ _430;
  wire _47105 = _47102 ^ _47104;
  wire _47106 = _47099 ^ _47105;
  wire _47107 = _47094 ^ _47106;
  wire _47108 = _3622 ^ _19251;
  wire _47109 = _3625 ^ _12712;
  wire _47110 = _47108 ^ _47109;
  wire _47111 = uncoded_block[923] ^ uncoded_block[932];
  wire _47112 = _3631 ^ _47111;
  wire _47113 = _1299 ^ _2084;
  wire _47114 = _47112 ^ _47113;
  wire _47115 = _47110 ^ _47114;
  wire _47116 = _17828 ^ _12175;
  wire _47117 = _47116 ^ _36089;
  wire _47118 = uncoded_block[969] ^ uncoded_block[971];
  wire _47119 = _2093 ^ _47118;
  wire _47120 = _2877 ^ _32425;
  wire _47121 = _47119 ^ _47120;
  wire _47122 = _47117 ^ _47121;
  wire _47123 = _47115 ^ _47122;
  wire _47124 = _5789 ^ _476;
  wire _47125 = _47124 ^ _3660;
  wire _47126 = _1318 ^ _4401;
  wire _47127 = _479 ^ _11101;
  wire _47128 = _47126 ^ _47127;
  wire _47129 = _47125 ^ _47128;
  wire _47130 = _2112 ^ _4405;
  wire _47131 = _18335 ^ _47130;
  wire _47132 = _4409 ^ _8296;
  wire _47133 = uncoded_block[1020] ^ uncoded_block[1024];
  wire _47134 = _9996 ^ _47133;
  wire _47135 = _47132 ^ _47134;
  wire _47136 = _47131 ^ _47135;
  wire _47137 = _47129 ^ _47136;
  wire _47138 = _47123 ^ _47137;
  wire _47139 = _47107 ^ _47138;
  wire _47140 = _47083 ^ _47139;
  wire _47141 = _47026 ^ _47140;
  wire _47142 = _18801 ^ _501;
  wire _47143 = _5810 ^ _38937;
  wire _47144 = _47142 ^ _47143;
  wire _47145 = _29410 ^ _23966;
  wire _47146 = uncoded_block[1065] ^ uncoded_block[1069];
  wire _47147 = _2916 ^ _47146;
  wire _47148 = _47145 ^ _47147;
  wire _47149 = _47144 ^ _47148;
  wire _47150 = _12770 ^ _6486;
  wire _47151 = _47150 ^ _25777;
  wire _47152 = _13858 ^ _36552;
  wire _47153 = _47151 ^ _47152;
  wire _47154 = _47149 ^ _47153;
  wire _47155 = _9484 ^ _2938;
  wire _47156 = _3714 ^ _4455;
  wire _47157 = _47155 ^ _47156;
  wire _47158 = _33312 ^ _8343;
  wire _47159 = _30329 ^ _25332;
  wire _47160 = _47158 ^ _47159;
  wire _47161 = _47157 ^ _47160;
  wire _47162 = _2180 ^ _2185;
  wire _47163 = _47162 ^ _5191;
  wire _47164 = _16897 ^ _22630;
  wire _47165 = _47163 ^ _47164;
  wire _47166 = _47161 ^ _47165;
  wire _47167 = _47154 ^ _47166;
  wire _47168 = _4481 ^ _17397;
  wire _47169 = _2196 ^ _3747;
  wire _47170 = _47168 ^ _47169;
  wire _47171 = _47170 ^ _7165;
  wire _47172 = _7765 ^ _1428;
  wire _47173 = _28297 ^ _47172;
  wire _47174 = _31219 ^ _6532;
  wire _47175 = _47174 ^ _13358;
  wire _47176 = _47173 ^ _47175;
  wire _47177 = _47171 ^ _47176;
  wire _47178 = _615 ^ _3772;
  wire _47179 = _47178 ^ _41312;
  wire _47180 = _1451 ^ _5901;
  wire _47181 = _5902 ^ _3004;
  wire _47182 = _47180 ^ _47181;
  wire _47183 = _47179 ^ _47182;
  wire _47184 = _3786 ^ _32500;
  wire _47185 = _47184 ^ _19364;
  wire _47186 = _3797 ^ _24482;
  wire _47187 = uncoded_block[1289] ^ uncoded_block[1299];
  wire _47188 = _47187 ^ _646;
  wire _47189 = _47186 ^ _47188;
  wire _47190 = _47185 ^ _47189;
  wire _47191 = _47183 ^ _47190;
  wire _47192 = _47177 ^ _47191;
  wire _47193 = _47167 ^ _47192;
  wire _47194 = _23134 ^ _14436;
  wire _47195 = _47194 ^ _22218;
  wire _47196 = _18436 ^ _40941;
  wire _47197 = _13402 ^ _47196;
  wire _47198 = _47195 ^ _47197;
  wire _47199 = _3045 ^ _1504;
  wire _47200 = _47199 ^ _37433;
  wire _47201 = _680 ^ _2289;
  wire _47202 = _47201 ^ _14964;
  wire _47203 = _47200 ^ _47202;
  wire _47204 = _47198 ^ _47203;
  wire _47205 = uncoded_block[1389] ^ uncoded_block[1396];
  wire _47206 = _47205 ^ _5293;
  wire _47207 = _32112 ^ _47206;
  wire _47208 = _14968 ^ _15489;
  wire _47209 = _40956 ^ _7844;
  wire _47210 = _47208 ^ _47209;
  wire _47211 = _47207 ^ _47210;
  wire _47212 = _22242 ^ _17470;
  wire _47213 = _19402 ^ _47212;
  wire _47214 = uncoded_block[1439] ^ uncoded_block[1444];
  wire _47215 = _47214 ^ _3084;
  wire _47216 = _47215 ^ _3866;
  wire _47217 = _47213 ^ _47216;
  wire _47218 = _47211 ^ _47217;
  wire _47219 = _47204 ^ _47218;
  wire _47220 = _4596 ^ _8455;
  wire _47221 = _19882 ^ _733;
  wire _47222 = _47220 ^ _47221;
  wire _47223 = _44354 ^ _42143;
  wire _47224 = _47222 ^ _47223;
  wire _47225 = _1565 ^ _3890;
  wire _47226 = _3109 ^ _41762;
  wire _47227 = _47225 ^ _47226;
  wire _47228 = uncoded_block[1509] ^ uncoded_block[1514];
  wire _47229 = _3894 ^ _47228;
  wire _47230 = uncoded_block[1517] ^ uncoded_block[1522];
  wire _47231 = _9621 ^ _47230;
  wire _47232 = _47229 ^ _47231;
  wire _47233 = _47227 ^ _47232;
  wire _47234 = _47224 ^ _47233;
  wire _47235 = uncoded_block[1529] ^ uncoded_block[1535];
  wire _47236 = _9626 ^ _47235;
  wire _47237 = _3906 ^ _6651;
  wire _47238 = _47236 ^ _47237;
  wire _47239 = _1589 ^ _30858;
  wire _47240 = _7277 ^ _24094;
  wire _47241 = _47239 ^ _47240;
  wire _47242 = _47238 ^ _47241;
  wire _47243 = uncoded_block[1566] ^ uncoded_block[1573];
  wire _47244 = _47243 ^ _6663;
  wire _47245 = _32158 ^ _47244;
  wire _47246 = _2383 ^ _32567;
  wire _47247 = _47246 ^ _22743;
  wire _47248 = _47245 ^ _47247;
  wire _47249 = _47242 ^ _47248;
  wire _47250 = _47234 ^ _47249;
  wire _47251 = _47219 ^ _47250;
  wire _47252 = _47193 ^ _47251;
  wire _47253 = uncoded_block[1608] ^ uncoded_block[1612];
  wire _47254 = _12373 ^ _47253;
  wire _47255 = _18014 ^ _47254;
  wire _47256 = _6042 ^ _6680;
  wire _47257 = _47256 ^ _41399;
  wire _47258 = _47255 ^ _47257;
  wire _47259 = _3942 ^ _19929;
  wire _47260 = _47259 ^ _40642;
  wire _47261 = _4674 ^ _13506;
  wire _47262 = _14529 ^ _47261;
  wire _47263 = _47260 ^ _47262;
  wire _47264 = _47258 ^ _47263;
  wire _47265 = _7319 ^ _19470;
  wire _47266 = _41411 ^ _47265;
  wire _47267 = _42187 ^ _3183;
  wire _47268 = _7325 ^ _10766;
  wire _47269 = _47267 ^ _47268;
  wire _47270 = _47266 ^ _47269;
  wire _47271 = _16058 ^ _35471;
  wire _47272 = _47271 ^ _30022;
  wire _47273 = uncoded_block[1700] ^ uncoded_block[1707];
  wire _47274 = _47273 ^ _11879;
  wire _47275 = _6072 ^ _2444;
  wire _47276 = _47274 ^ _47275;
  wire _47277 = _47272 ^ _47276;
  wire _47278 = _47270 ^ _47277;
  wire _47279 = _47264 ^ _47278;
  wire _47280 = _47279 ^ uncoded_block[1722];
  wire _47281 = _47252 ^ _47280;
  wire _47282 = _47141 ^ _47281;
  wire _47283 = _2453 ^ _4;
  wire _47284 = _46150 ^ _3217;
  wire _47285 = _47283 ^ _47284;
  wire _47286 = _25940 ^ _22330;
  wire _47287 = _47285 ^ _47286;
  wire _47288 = _3227 ^ _7965;
  wire _47289 = uncoded_block[45] ^ uncoded_block[51];
  wire _47290 = _47289 ^ _1700;
  wire _47291 = _47288 ^ _47290;
  wire _47292 = _7364 ^ _1705;
  wire _47293 = _2475 ^ _7367;
  wire _47294 = _47292 ^ _47293;
  wire _47295 = _47291 ^ _47294;
  wire _47296 = _47287 ^ _47295;
  wire _47297 = _14060 ^ _22805;
  wire _47298 = _17578 ^ _42;
  wire _47299 = _47297 ^ _47298;
  wire _47300 = _4026 ^ _15097;
  wire _47301 = _7986 ^ _17584;
  wire _47302 = _47300 ^ _47301;
  wire _47303 = _47299 ^ _47302;
  wire _47304 = _1722 ^ _5453;
  wire _47305 = _47304 ^ _18565;
  wire _47306 = _3256 ^ _4042;
  wire _47307 = uncoded_block[135] ^ uncoded_block[139];
  wire _47308 = _47307 ^ _11918;
  wire _47309 = _47306 ^ _47308;
  wire _47310 = _47305 ^ _47309;
  wire _47311 = _47303 ^ _47310;
  wire _47312 = _47296 ^ _47311;
  wire _47313 = _15114 ^ _17097;
  wire _47314 = _1744 ^ _8003;
  wire _47315 = _47313 ^ _47314;
  wire _47316 = _16604 ^ _81;
  wire _47317 = _42884 ^ _47316;
  wire _47318 = _47315 ^ _47317;
  wire _47319 = _19539 ^ _2524;
  wire _47320 = uncoded_block[181] ^ uncoded_block[185];
  wire _47321 = _47320 ^ _4773;
  wire _47322 = _47319 ^ _47321;
  wire _47323 = _15135 ^ _5486;
  wire _47324 = _33496 ^ _47323;
  wire _47325 = _47322 ^ _47324;
  wire _47326 = _47318 ^ _47325;
  wire _47327 = _959 ^ _101;
  wire _47328 = _47327 ^ _46958;
  wire _47329 = _15143 ^ _45193;
  wire _47330 = _47328 ^ _47329;
  wire _47331 = _8612 ^ _6179;
  wire _47332 = _47331 ^ _20998;
  wire _47333 = _4095 ^ _4098;
  wire _47334 = _30542 ^ _47333;
  wire _47335 = _47332 ^ _47334;
  wire _47336 = _47330 ^ _47335;
  wire _47337 = _47326 ^ _47336;
  wire _47338 = _47312 ^ _47337;
  wire _47339 = _7440 ^ _14642;
  wire _47340 = _10872 ^ _2568;
  wire _47341 = _47339 ^ _47340;
  wire _47342 = _20527 ^ _40716;
  wire _47343 = _15159 ^ _4819;
  wire _47344 = _47342 ^ _47343;
  wire _47345 = _47341 ^ _47344;
  wire _47346 = _4820 ^ _1807;
  wire _47347 = _1810 ^ _4111;
  wire _47348 = _47346 ^ _47347;
  wire _47349 = _1000 ^ _8056;
  wire _47350 = _3340 ^ _1818;
  wire _47351 = _47349 ^ _47350;
  wire _47352 = _47348 ^ _47351;
  wire _47353 = _47345 ^ _47352;
  wire _47354 = _18147 ^ _1821;
  wire _47355 = _3353 ^ _161;
  wire _47356 = _47354 ^ _47355;
  wire _47357 = _11990 ^ _6221;
  wire _47358 = _6227 ^ _21030;
  wire _47359 = _47357 ^ _47358;
  wire _47360 = _47356 ^ _47359;
  wire _47361 = _8079 ^ _20056;
  wire _47362 = _3370 ^ _47361;
  wire _47363 = _19599 ^ _7483;
  wire _47364 = _20058 ^ _47363;
  wire _47365 = _47362 ^ _47364;
  wire _47366 = _47360 ^ _47365;
  wire _47367 = _47353 ^ _47366;
  wire _47368 = _19604 ^ _2623;
  wire _47369 = _5559 ^ _41525;
  wire _47370 = _47368 ^ _47369;
  wire _47371 = uncoded_block[409] ^ uncoded_block[414];
  wire _47372 = _47371 ^ _5565;
  wire _47373 = _13112 ^ _4872;
  wire _47374 = _47372 ^ _47373;
  wire _47375 = _47370 ^ _47374;
  wire _47376 = _32702 ^ _6254;
  wire _47377 = _47376 ^ _30589;
  wire _47378 = _4176 ^ _1070;
  wire _47379 = _1075 ^ _30591;
  wire _47380 = _47378 ^ _47379;
  wire _47381 = _47377 ^ _47380;
  wire _47382 = _47375 ^ _47381;
  wire _47383 = _29702 ^ _12028;
  wire _47384 = _16691 ^ _47383;
  wire _47385 = _17197 ^ _26950;
  wire _47386 = _47384 ^ _47385;
  wire _47387 = _229 ^ _9295;
  wire _47388 = _26952 ^ _47387;
  wire _47389 = _32722 ^ _10947;
  wire _47390 = _10948 ^ _16711;
  wire _47391 = _47389 ^ _47390;
  wire _47392 = _47388 ^ _47391;
  wire _47393 = _47386 ^ _47392;
  wire _47394 = _47382 ^ _47393;
  wire _47395 = _47367 ^ _47394;
  wire _47396 = _47338 ^ _47395;
  wire _47397 = _31482 ^ _4928;
  wire _47398 = _2684 ^ _5628;
  wire _47399 = _4933 ^ _6304;
  wire _47400 = _47398 ^ _47399;
  wire _47401 = _47397 ^ _47400;
  wire _47402 = _31907 ^ _3465;
  wire _47403 = _1927 ^ _23387;
  wire _47404 = _47402 ^ _47403;
  wire _47405 = _11526 ^ _9325;
  wire _47406 = _47405 ^ _44911;
  wire _47407 = _47404 ^ _47406;
  wire _47408 = _47401 ^ _47407;
  wire _47409 = _8148 ^ _4952;
  wire _47410 = _47409 ^ _1147;
  wire _47411 = _41570 ^ _5652;
  wire _47412 = _13178 ^ _20125;
  wire _47413 = _47411 ^ _47412;
  wire _47414 = _47410 ^ _47413;
  wire _47415 = _12618 ^ _5658;
  wire _47416 = _14745 ^ _290;
  wire _47417 = _47415 ^ _47416;
  wire _47418 = _44551 ^ _39633;
  wire _47419 = _47417 ^ _47418;
  wire _47420 = _47414 ^ _47419;
  wire _47421 = _47408 ^ _47420;
  wire _47422 = _19181 ^ _18705;
  wire _47423 = _1173 ^ _17742;
  wire _47424 = _47422 ^ _47423;
  wire _47425 = _1181 ^ _5678;
  wire _47426 = _11553 ^ _47425;
  wire _47427 = _47424 ^ _47426;
  wire _47428 = _22491 ^ _12093;
  wire _47429 = _13740 ^ _10447;
  wire _47430 = _3535 ^ _1194;
  wire _47431 = _47429 ^ _47430;
  wire _47432 = _47428 ^ _47431;
  wire _47433 = _47427 ^ _47432;
  wire _47434 = _6367 ^ _5691;
  wire _47435 = _47434 ^ _45699;
  wire _47436 = _7605 ^ _2770;
  wire _47437 = uncoded_block[741] ^ uncoded_block[749];
  wire _47438 = _47437 ^ _1214;
  wire _47439 = _47436 ^ _47438;
  wire _47440 = _47435 ^ _47439;
  wire _47441 = _11012 ^ _9914;
  wire _47442 = _2784 ^ _14278;
  wire _47443 = _47441 ^ _47442;
  wire _47444 = _13219 ^ _18277;
  wire _47445 = _372 ^ _374;
  wire _47446 = _47444 ^ _47445;
  wire _47447 = _47443 ^ _47446;
  wire _47448 = _47440 ^ _47447;
  wire _47449 = _47433 ^ _47448;
  wire _47450 = _47421 ^ _47449;
  wire _47451 = _12125 ^ _11595;
  wire _47452 = uncoded_block[811] ^ uncoded_block[816];
  wire _47453 = _47452 ^ _7634;
  wire _47454 = _3587 ^ _34067;
  wire _47455 = _47453 ^ _47454;
  wire _47456 = _47451 ^ _47455;
  wire _47457 = _16801 ^ _12138;
  wire _47458 = _4337 ^ _5057;
  wire _47459 = _47457 ^ _47458;
  wire _47460 = _8808 ^ _4340;
  wire _47461 = _47460 ^ _46329;
  wire _47462 = _47459 ^ _47461;
  wire _47463 = _47456 ^ _47462;
  wire _47464 = uncoded_block[856] ^ uncoded_block[860];
  wire _47465 = _47464 ^ _9948;
  wire _47466 = _47465 ^ _22087;
  wire _47467 = _6416 ^ _11620;
  wire _47468 = _47467 ^ _22090;
  wire _47469 = _47466 ^ _47468;
  wire _47470 = _11059 ^ _15342;
  wire _47471 = _1277 ^ _5758;
  wire _47472 = _47470 ^ _47471;
  wire _47473 = _5759 ^ _2065;
  wire _47474 = uncoded_block[911] ^ uncoded_block[917];
  wire _47475 = _47474 ^ _18775;
  wire _47476 = _47473 ^ _47475;
  wire _47477 = _47472 ^ _47476;
  wire _47478 = _47469 ^ _47477;
  wire _47479 = _47463 ^ _47478;
  wire _47480 = _4368 ^ _4370;
  wire _47481 = uncoded_block[928] ^ uncoded_block[933];
  wire _47482 = _47481 ^ _2079;
  wire _47483 = _47480 ^ _47482;
  wire _47484 = uncoded_block[953] ^ uncoded_block[960];
  wire _47485 = _4381 ^ _47484;
  wire _47486 = _38111 ^ _47485;
  wire _47487 = _47483 ^ _47486;
  wire _47488 = _16330 ^ _2094;
  wire _47489 = _3656 ^ _4390;
  wire _47490 = uncoded_block[978] ^ uncoded_block[983];
  wire _47491 = _5114 ^ _47490;
  wire _47492 = _47489 ^ _47491;
  wire _47493 = _47488 ^ _47492;
  wire _47494 = _47487 ^ _47493;
  wire _47495 = _7093 ^ _14850;
  wire _47496 = _47495 ^ _28238;
  wire _47497 = _484 ^ _13835;
  wire _47498 = _12739 ^ _47497;
  wire _47499 = _47496 ^ _47498;
  wire _47500 = _494 ^ _8874;
  wire _47501 = _31602 ^ _47500;
  wire _47502 = _8875 ^ _5806;
  wire _47503 = _47502 ^ _32023;
  wire _47504 = _47501 ^ _47503;
  wire _47505 = _47499 ^ _47504;
  wire _47506 = _47494 ^ _47505;
  wire _47507 = _47479 ^ _47506;
  wire _47508 = _47450 ^ _47507;
  wire _47509 = _47396 ^ _47508;
  wire _47510 = _38940 ^ _9466;
  wire _47511 = _1363 ^ _5825;
  wire _47512 = _2142 ^ _25773;
  wire _47513 = _47511 ^ _47512;
  wire _47514 = _47510 ^ _47513;
  wire _47515 = _527 ^ _5832;
  wire _47516 = uncoded_block[1080] ^ uncoded_block[1087];
  wire _47517 = _47516 ^ _12774;
  wire _47518 = _47515 ^ _47517;
  wire _47519 = _5840 ^ _5842;
  wire _47520 = _40884 ^ _2161;
  wire _47521 = _47519 ^ _47520;
  wire _47522 = _47518 ^ _47521;
  wire _47523 = _47514 ^ _47522;
  wire _47524 = uncoded_block[1118] ^ uncoded_block[1123];
  wire _47525 = _15890 ^ _47524;
  wire _47526 = _2944 ^ _23523;
  wire _47527 = _47525 ^ _47526;
  wire _47528 = _15896 ^ _14380;
  wire _47529 = _20269 ^ _32468;
  wire _47530 = _47528 ^ _47529;
  wire _47531 = _47527 ^ _47530;
  wire _47532 = _11711 ^ _2958;
  wire _47533 = _13876 ^ _47532;
  wire _47534 = _24444 ^ _29882;
  wire _47535 = _47533 ^ _47534;
  wire _47536 = _47531 ^ _47535;
  wire _47537 = _47523 ^ _47536;
  wire _47538 = _17396 ^ _1417;
  wire _47539 = _47538 ^ _16395;
  wire _47540 = _24910 ^ _21259;
  wire _47541 = _2206 ^ _3755;
  wire _47542 = _47540 ^ _47541;
  wire _47543 = _47539 ^ _47542;
  wire _47544 = _2217 ^ _1428;
  wire _47545 = _3763 ^ _10059;
  wire _47546 = _47544 ^ _47545;
  wire _47547 = _5218 ^ _31228;
  wire _47548 = _47547 ^ _9524;
  wire _47549 = _47546 ^ _47548;
  wire _47550 = _47543 ^ _47549;
  wire _47551 = uncoded_block[1245] ^ uncoded_block[1250];
  wire _47552 = _10627 ^ _47551;
  wire _47553 = _47552 ^ _45816;
  wire _47554 = _13369 ^ _3004;
  wire _47555 = _7788 ^ _5905;
  wire _47556 = _47554 ^ _47555;
  wire _47557 = _47553 ^ _47556;
  wire _47558 = _3794 ^ _6557;
  wire _47559 = _44694 ^ _47558;
  wire _47560 = _28317 ^ _11195;
  wire _47561 = _7193 ^ _17927;
  wire _47562 = _47560 ^ _47561;
  wire _47563 = _47559 ^ _47562;
  wire _47564 = _47557 ^ _47563;
  wire _47565 = _47550 ^ _47564;
  wire _47566 = _47537 ^ _47565;
  wire _47567 = _2254 ^ _3807;
  wire _47568 = _17435 ^ _26726;
  wire _47569 = _47567 ^ _47568;
  wire _47570 = _20319 ^ _5929;
  wire _47571 = _47569 ^ _47570;
  wire _47572 = _6578 ^ _2276;
  wire _47573 = _47572 ^ _33783;
  wire _47574 = uncoded_block[1347] ^ uncoded_block[1354];
  wire _47575 = _47574 ^ _12857;
  wire _47576 = _7821 ^ _1504;
  wire _47577 = _47575 ^ _47576;
  wire _47578 = _47573 ^ _47577;
  wire _47579 = _47571 ^ _47578;
  wire _47580 = _10103 ^ _5285;
  wire _47581 = _3048 ^ _47580;
  wire _47582 = _3059 ^ _688;
  wire _47583 = _47582 ^ _24512;
  wire _47584 = _47581 ^ _47583;
  wire _47585 = _25856 ^ _8435;
  wire _47586 = _47585 ^ _16958;
  wire _47587 = _16463 ^ _9588;
  wire _47588 = _2308 ^ _23604;
  wire _47589 = _47587 ^ _47588;
  wire _47590 = _47586 ^ _47589;
  wire _47591 = _47584 ^ _47590;
  wire _47592 = _47579 ^ _47591;
  wire _47593 = _3081 ^ _14978;
  wire _47594 = _3861 ^ _5305;
  wire _47595 = _47593 ^ _47594;
  wire _47596 = _3088 ^ _4596;
  wire _47597 = _36636 ^ _47596;
  wire _47598 = _47595 ^ _47597;
  wire _47599 = _8455 ^ _10136;
  wire _47600 = uncoded_block[1480] ^ uncoded_block[1487];
  wire _47601 = _735 ^ _47600;
  wire _47602 = _47599 ^ _47601;
  wire _47603 = uncoded_block[1498] ^ uncoded_block[1504];
  wire _47604 = _12898 ^ _47603;
  wire _47605 = _24536 ^ _47604;
  wire _47606 = _47602 ^ _47605;
  wire _47607 = _47598 ^ _47606;
  wire _47608 = _1574 ^ _6642;
  wire _47609 = _47608 ^ _46472;
  wire _47610 = uncoded_block[1522] ^ uncoded_block[1527];
  wire _47611 = _47610 ^ _8474;
  wire _47612 = _12914 ^ _1587;
  wire _47613 = _47611 ^ _47612;
  wire _47614 = _47609 ^ _47613;
  wire _47615 = _3909 ^ _2367;
  wire _47616 = _47615 ^ _19438;
  wire _47617 = _28378 ^ _31732;
  wire _47618 = _47617 ^ _25447;
  wire _47619 = _47616 ^ _47618;
  wire _47620 = _47614 ^ _47619;
  wire _47621 = _47607 ^ _47620;
  wire _47622 = _47592 ^ _47621;
  wire _47623 = _47566 ^ _47622;
  wire _47624 = _16510 ^ _15026;
  wire _47625 = uncoded_block[1576] ^ uncoded_block[1579];
  wire _47626 = _4647 ^ _47625;
  wire _47627 = _47624 ^ _47626;
  wire _47628 = _18952 ^ _788;
  wire _47629 = _47628 ^ _3147;
  wire _47630 = _47627 ^ _47629;
  wire _47631 = _11294 ^ _8502;
  wire _47632 = _1625 ^ _1627;
  wire _47633 = _47631 ^ _47632;
  wire _47634 = uncoded_block[1615] ^ uncoded_block[1621];
  wire _47635 = uncoded_block[1622] ^ uncoded_block[1626];
  wire _47636 = _47634 ^ _47635;
  wire _47637 = _33843 ^ _47636;
  wire _47638 = _47633 ^ _47637;
  wire _47639 = _47630 ^ _47638;
  wire _47640 = _2404 ^ _20900;
  wire _47641 = _13500 ^ _1647;
  wire _47642 = _47640 ^ _47641;
  wire _47643 = _11313 ^ _21385;
  wire _47644 = _47642 ^ _47643;
  wire _47645 = _16052 ^ _6059;
  wire _47646 = _20911 ^ _47645;
  wire _47647 = _12398 ^ _5406;
  wire _47648 = _3190 ^ _6066;
  wire _47649 = _47647 ^ _47648;
  wire _47650 = _47646 ^ _47649;
  wire _47651 = _47644 ^ _47650;
  wire _47652 = _47639 ^ _47651;
  wire _47653 = _3972 ^ _845;
  wire _47654 = _16551 ^ _854;
  wire _47655 = _47653 ^ _47654;
  wire _47656 = _47655 ^ _10217;
  wire _47657 = _47652 ^ _47656;
  wire _47658 = _47623 ^ _47657;
  wire _47659 = _47509 ^ _47658;
  wire _47660 = _3210 ^ _32201;
  wire _47661 = _6724 ^ _6083;
  wire _47662 = _47660 ^ _47661;
  wire _47663 = _8 ^ _10226;
  wire _47664 = _872 ^ _23249;
  wire _47665 = _47663 ^ _47664;
  wire _47666 = _47662 ^ _47665;
  wire _47667 = _11 ^ _14569;
  wire _47668 = _18 ^ _14571;
  wire _47669 = _47667 ^ _47668;
  wire _47670 = _32212 ^ _38299;
  wire _47671 = _19503 ^ _47670;
  wire _47672 = _47669 ^ _47671;
  wire _47673 = _47666 ^ _47672;
  wire _47674 = _2472 ^ _10806;
  wire _47675 = uncoded_block[65] ^ uncoded_block[79];
  wire _47676 = _47675 ^ _11364;
  wire _47677 = _47674 ^ _47676;
  wire _47678 = _17578 ^ _9713;
  wire _47679 = _903 ^ _6758;
  wire _47680 = _47678 ^ _47679;
  wire _47681 = _47677 ^ _47680;
  wire _47682 = _9718 ^ _7377;
  wire _47683 = _9166 ^ _6126;
  wire _47684 = _47682 ^ _47683;
  wire _47685 = _6769 ^ _29611;
  wire _47686 = _2502 ^ _917;
  wire _47687 = _47685 ^ _47686;
  wire _47688 = _47684 ^ _47687;
  wire _47689 = _47681 ^ _47688;
  wire _47690 = _47673 ^ _47689;
  wire _47691 = _1736 ^ _64;
  wire _47692 = _20964 ^ _47691;
  wire _47693 = _16600 ^ _6780;
  wire _47694 = _5469 ^ _2514;
  wire _47695 = _47693 ^ _47694;
  wire _47696 = _47692 ^ _47695;
  wire _47697 = _74 ^ _11928;
  wire _47698 = _5473 ^ _19539;
  wire _47699 = _47697 ^ _47698;
  wire _47700 = _10272 ^ _34716;
  wire _47701 = _47699 ^ _47700;
  wire _47702 = _47696 ^ _47701;
  wire _47703 = _20010 ^ _22839;
  wire _47704 = _21919 ^ _4787;
  wire _47705 = _104 ^ _6814;
  wire _47706 = _47704 ^ _47705;
  wire _47707 = _47703 ^ _47706;
  wire _47708 = _1774 ^ _6824;
  wire _47709 = _47708 ^ _37956;
  wire _47710 = uncoded_block[269] ^ uncoded_block[274];
  wire _47711 = _8620 ^ _47710;
  wire _47712 = _34730 ^ _47711;
  wire _47713 = _47709 ^ _47712;
  wire _47714 = _47707 ^ _47713;
  wire _47715 = _47702 ^ _47714;
  wire _47716 = _47690 ^ _47715;
  wire _47717 = _43314 ^ _11425;
  wire _47718 = _29238 ^ _28817;
  wire _47719 = _17635 ^ _4111;
  wire _47720 = _47718 ^ _47719;
  wire _47721 = _47717 ^ _47720;
  wire _47722 = _17639 ^ _5528;
  wire _47723 = _47722 ^ _12518;
  wire _47724 = _8058 ^ _11983;
  wire _47725 = _47724 ^ _35556;
  wire _47726 = _47723 ^ _47725;
  wire _47727 = _47721 ^ _47726;
  wire _47728 = _1825 ^ _6217;
  wire _47729 = _3355 ^ _7465;
  wire _47730 = _47728 ^ _47729;
  wire _47731 = _2601 ^ _39567;
  wire _47732 = _16657 ^ _47731;
  wire _47733 = _47730 ^ _47732;
  wire _47734 = uncoded_block[372] ^ uncoded_block[376];
  wire _47735 = _1838 ^ _47734;
  wire _47736 = _4854 ^ _1841;
  wire _47737 = _47735 ^ _47736;
  wire _47738 = _1842 ^ _4149;
  wire _47739 = _3381 ^ _12541;
  wire _47740 = _47738 ^ _47739;
  wire _47741 = _47737 ^ _47740;
  wire _47742 = _47733 ^ _47741;
  wire _47743 = _47727 ^ _47742;
  wire _47744 = _177 ^ _2622;
  wire _47745 = _16177 ^ _190;
  wire _47746 = _47744 ^ _47745;
  wire _47747 = _3394 ^ _4871;
  wire _47748 = _24248 ^ _34771;
  wire _47749 = _47747 ^ _47748;
  wire _47750 = _47746 ^ _47749;
  wire _47751 = uncoded_block[433] ^ uncoded_block[441];
  wire _47752 = _47751 ^ _206;
  wire _47753 = _3409 ^ _1867;
  wire _47754 = _47752 ^ _47753;
  wire _47755 = _1870 ^ _3415;
  wire _47756 = _2653 ^ _10927;
  wire _47757 = _47755 ^ _47756;
  wire _47758 = _47754 ^ _47757;
  wire _47759 = _47750 ^ _47758;
  wire _47760 = _5590 ^ _5598;
  wire _47761 = _3419 ^ _47760;
  wire _47762 = _5603 ^ _6279;
  wire _47763 = _17691 ^ _47762;
  wire _47764 = _47761 ^ _47763;
  wire _47765 = _1887 ^ _3437;
  wire _47766 = _9840 ^ _3444;
  wire _47767 = _47765 ^ _47766;
  wire _47768 = _22924 ^ _1111;
  wire _47769 = uncoded_block[534] ^ uncoded_block[539];
  wire _47770 = _9309 ^ _47769;
  wire _47771 = _47768 ^ _47770;
  wire _47772 = _47767 ^ _47771;
  wire _47773 = _47764 ^ _47772;
  wire _47774 = _47759 ^ _47773;
  wire _47775 = _47743 ^ _47774;
  wire _47776 = _47716 ^ _47775;
  wire _47777 = _14721 ^ _246;
  wire _47778 = _47777 ^ _16719;
  wire _47779 = _40776 ^ _38416;
  wire _47780 = _47778 ^ _47779;
  wire _47781 = uncoded_block[574] ^ uncoded_block[579];
  wire _47782 = _13698 ^ _47781;
  wire _47783 = _11527 ^ _1141;
  wire _47784 = _47782 ^ _47783;
  wire _47785 = _2709 ^ _16233;
  wire _47786 = _41566 ^ _47785;
  wire _47787 = _47784 ^ _47786;
  wire _47788 = _47780 ^ _47787;
  wire _47789 = _7564 ^ _14743;
  wire _47790 = _2720 ^ _8749;
  wire _47791 = _47789 ^ _47790;
  wire _47792 = _1161 ^ _12624;
  wire _47793 = _47792 ^ _12626;
  wire _47794 = _47791 ^ _47793;
  wire _47795 = _20638 ^ _5671;
  wire _47796 = _40796 ^ _47795;
  wire _47797 = _9886 ^ _2748;
  wire _47798 = _8177 ^ _1971;
  wire _47799 = _47797 ^ _47798;
  wire _47800 = _47796 ^ _47799;
  wire _47801 = _47794 ^ _47800;
  wire _47802 = _47788 ^ _47801;
  wire _47803 = _2750 ^ _4271;
  wire _47804 = _47803 ^ _34436;
  wire _47805 = _4989 ^ _14255;
  wire _47806 = _10448 ^ _33205;
  wire _47807 = _47805 ^ _47806;
  wire _47808 = _47804 ^ _47807;
  wire _47809 = uncoded_block[715] ^ uncoded_block[722];
  wire _47810 = _47809 ^ _9904;
  wire _47811 = _5693 ^ _5005;
  wire _47812 = _47810 ^ _47811;
  wire _47813 = _1206 ^ _2770;
  wire _47814 = _5699 ^ _5013;
  wire _47815 = _47813 ^ _47814;
  wire _47816 = _47812 ^ _47815;
  wire _47817 = _47808 ^ _47816;
  wire _47818 = _2777 ^ _11012;
  wire _47819 = _17774 ^ _8781;
  wire _47820 = _47818 ^ _47819;
  wire _47821 = _17776 ^ _2791;
  wire _47822 = _2792 ^ _368;
  wire _47823 = _47821 ^ _47822;
  wire _47824 = _47820 ^ _47823;
  wire _47825 = _25691 ^ _3570;
  wire _47826 = _1225 ^ _2799;
  wire _47827 = _47825 ^ _47826;
  wire _47828 = _6392 ^ _9395;
  wire _47829 = _47827 ^ _47828;
  wire _47830 = _47824 ^ _47829;
  wire _47831 = _47817 ^ _47830;
  wire _47832 = _47802 ^ _47831;
  wire _47833 = _16793 ^ _31971;
  wire _47834 = _2029 ^ _37698;
  wire _47835 = _47833 ^ _47834;
  wire _47836 = uncoded_block[838] ^ uncoded_block[841];
  wire _47837 = _23003 ^ _47836;
  wire _47838 = _34470 ^ _12141;
  wire _47839 = _47837 ^ _47838;
  wire _47840 = _47835 ^ _47839;
  wire _47841 = _15330 ^ _7649;
  wire _47842 = _7650 ^ _35281;
  wire _47843 = _47841 ^ _47842;
  wire _47844 = _33671 ^ _41628;
  wire _47845 = _11056 ^ _2059;
  wire _47846 = _47844 ^ _47845;
  wire _47847 = _47843 ^ _47846;
  wire _47848 = _47840 ^ _47847;
  wire _47849 = _11060 ^ _8826;
  wire _47850 = _28965 ^ _2065;
  wire _47851 = _47849 ^ _47850;
  wire _47852 = _46723 ^ _21644;
  wire _47853 = _16310 ^ _47852;
  wire _47854 = _47851 ^ _47853;
  wire _47855 = _39692 ^ _2076;
  wire _47856 = _9968 ^ _5096;
  wire _47857 = _47855 ^ _47856;
  wire _47858 = _5102 ^ _16834;
  wire _47859 = _47857 ^ _47858;
  wire _47860 = _47854 ^ _47859;
  wire _47861 = _47848 ^ _47860;
  wire _47862 = _29387 ^ _8275;
  wire _47863 = uncoded_block[960] ^ uncoded_block[964];
  wire _47864 = _7680 ^ _47863;
  wire _47865 = _47862 ^ _47864;
  wire _47866 = _6447 ^ _468;
  wire _47867 = _4390 ^ _5114;
  wire _47868 = _47866 ^ _47867;
  wire _47869 = _47865 ^ _47868;
  wire _47870 = _3660 ^ _43083;
  wire _47871 = uncoded_block[995] ^ uncoded_block[999];
  wire _47872 = _47871 ^ _24858;
  wire _47873 = _484 ^ _4409;
  wire _47874 = _47872 ^ _47873;
  wire _47875 = _47870 ^ _47874;
  wire _47876 = _47869 ^ _47875;
  wire _47877 = _37743 ^ _9996;
  wire _47878 = _47877 ^ _26649;
  wire _47879 = _13288 ^ _34925;
  wire _47880 = _35319 ^ _47879;
  wire _47881 = _47878 ^ _47880;
  wire _47882 = _21219 ^ _36542;
  wire _47883 = _12762 ^ _7117;
  wire _47884 = _4433 ^ _3685;
  wire _47885 = _47883 ^ _47884;
  wire _47886 = _47882 ^ _47885;
  wire _47887 = _47881 ^ _47886;
  wire _47888 = _47876 ^ _47887;
  wire _47889 = _47861 ^ _47888;
  wire _47890 = _47832 ^ _47889;
  wire _47891 = _47776 ^ _47890;
  wire _47892 = _12213 ^ _527;
  wire _47893 = _47892 ^ _15882;
  wire _47894 = _3696 ^ _12774;
  wire _47895 = _37371 ^ _47894;
  wire _47896 = _47893 ^ _47895;
  wire _47897 = _5840 ^ _8330;
  wire _47898 = uncoded_block[1106] ^ uncoded_block[1113];
  wire _47899 = _3707 ^ _47898;
  wire _47900 = _47897 ^ _47899;
  wire _47901 = _13323 ^ _8921;
  wire _47902 = _47900 ^ _47901;
  wire _47903 = _47896 ^ _47902;
  wire _47904 = _2942 ^ _18832;
  wire _47905 = _19322 ^ _4462;
  wire _47906 = _47904 ^ _47905;
  wire _47907 = _14383 ^ _24900;
  wire _47908 = _47906 ^ _47907;
  wire _47909 = _32056 ^ _3728;
  wire _47910 = _47909 ^ _16892;
  wire _47911 = _26244 ^ _11160;
  wire _47912 = _47911 ^ _22630;
  wire _47913 = _47910 ^ _47912;
  wire _47914 = _47908 ^ _47913;
  wire _47915 = _47903 ^ _47914;
  wire _47916 = _24450 ^ _30764;
  wire _47917 = _5201 ^ _5203;
  wire _47918 = _16397 ^ _2206;
  wire _47919 = _47917 ^ _47918;
  wire _47920 = _47916 ^ _47919;
  wire _47921 = _14910 ^ _7767;
  wire _47922 = _5215 ^ _6532;
  wire _47923 = _47922 ^ _13358;
  wire _47924 = _47921 ^ _47923;
  wire _47925 = _47920 ^ _47924;
  wire _47926 = _43145 ^ _8385;
  wire _47927 = _7175 ^ _47926;
  wire _47928 = _44300 ^ _5234;
  wire _47929 = _47928 ^ _38581;
  wire _47930 = _47927 ^ _47929;
  wire _47931 = _1459 ^ _10075;
  wire _47932 = _30786 ^ _47931;
  wire _47933 = _5908 ^ _3794;
  wire _47934 = _12837 ^ _2251;
  wire _47935 = _47933 ^ _47934;
  wire _47936 = _47932 ^ _47935;
  wire _47937 = _47930 ^ _47936;
  wire _47938 = _47925 ^ _47937;
  wire _47939 = _47915 ^ _47938;
  wire _47940 = _5246 ^ _2254;
  wire _47941 = _47940 ^ _24485;
  wire _47942 = _14430 ^ _5926;
  wire _47943 = _24938 ^ _47942;
  wire _47944 = _47941 ^ _47943;
  wire _47945 = uncoded_block[1322] ^ uncoded_block[1324];
  wire _47946 = _9555 ^ _47945;
  wire _47947 = _47946 ^ _658;
  wire _47948 = _5931 ^ _9563;
  wire _47949 = _47948 ^ _43546;
  wire _47950 = _47947 ^ _47949;
  wire _47951 = _47944 ^ _47950;
  wire _47952 = _1501 ^ _3041;
  wire _47953 = _33363 ^ _15477;
  wire _47954 = _47952 ^ _47953;
  wire _47955 = _3047 ^ _4563;
  wire _47956 = _46438 ^ _47955;
  wire _47957 = _47954 ^ _47956;
  wire _47958 = _22229 ^ _3834;
  wire _47959 = _47958 ^ _25851;
  wire _47960 = uncoded_block[1389] ^ uncoded_block[1393];
  wire _47961 = _47960 ^ _4571;
  wire _47962 = _47961 ^ _29943;
  wire _47963 = _47959 ^ _47962;
  wire _47964 = _47957 ^ _47963;
  wire _47965 = _47951 ^ _47964;
  wire _47966 = _4578 ^ _4580;
  wire _47967 = uncoded_block[1414] ^ uncoded_block[1417];
  wire _47968 = _47967 ^ _10120;
  wire _47969 = _47966 ^ _47968;
  wire _47970 = uncoded_block[1429] ^ uncoded_block[1435];
  wire _47971 = _11239 ^ _47970;
  wire _47972 = _36206 ^ _47971;
  wire _47973 = _47969 ^ _47972;
  wire _47974 = _1540 ^ _2321;
  wire _47975 = _16473 ^ _6620;
  wire _47976 = _47974 ^ _47975;
  wire _47977 = _16474 ^ _3088;
  wire _47978 = _726 ^ _20855;
  wire _47979 = _47977 ^ _47978;
  wire _47980 = _47976 ^ _47979;
  wire _47981 = _47973 ^ _47980;
  wire _47982 = _2338 ^ _733;
  wire _47983 = uncoded_block[1478] ^ uncoded_block[1484];
  wire _47984 = _735 ^ _47983;
  wire _47985 = _47982 ^ _47984;
  wire _47986 = _2349 ^ _5329;
  wire _47987 = _3890 ^ _3109;
  wire _47988 = _47986 ^ _47987;
  wire _47989 = _47985 ^ _47988;
  wire _47990 = _748 ^ _4616;
  wire _47991 = _15002 ^ _6642;
  wire _47992 = _47990 ^ _47991;
  wire _47993 = _27622 ^ _39436;
  wire _47994 = _47992 ^ _47993;
  wire _47995 = _47989 ^ _47994;
  wire _47996 = _47981 ^ _47995;
  wire _47997 = _47965 ^ _47996;
  wire _47998 = _47939 ^ _47997;
  wire _47999 = _15007 ^ _9064;
  wire _48000 = _19903 ^ _1590;
  wire _48001 = _47999 ^ _48000;
  wire _48002 = _9070 ^ _7888;
  wire _48003 = _23637 ^ _48002;
  wire _48004 = _48001 ^ _48003;
  wire _48005 = _2372 ^ _6019;
  wire _48006 = uncoded_block[1571] ^ uncoded_block[1577];
  wire _48007 = _16510 ^ _48006;
  wire _48008 = _48005 ^ _48007;
  wire _48009 = _25008 ^ _5371;
  wire _48010 = _24105 ^ _48009;
  wire _48011 = _48008 ^ _48010;
  wire _48012 = _48004 ^ _48011;
  wire _48013 = _3151 ^ _1625;
  wire _48014 = _18012 ^ _48013;
  wire _48015 = _25905 ^ _805;
  wire _48016 = _22290 ^ _48015;
  wire _48017 = _48014 ^ _48016;
  wire _48018 = _3941 ^ _12947;
  wire _48019 = _48018 ^ _1640;
  wire _48020 = _3949 ^ _42179;
  wire _48021 = _48019 ^ _48020;
  wire _48022 = _48017 ^ _48021;
  wire _48023 = _48012 ^ _48022;
  wire _48024 = _17529 ^ _820;
  wire _48025 = _822 ^ _17032;
  wire _48026 = _48024 ^ _48025;
  wire _48027 = _1662 ^ _9113;
  wire _48028 = _31761 ^ _48027;
  wire _48029 = _48026 ^ _48028;
  wire _48030 = _4693 ^ _14543;
  wire _48031 = _48030 ^ _3191;
  wire _48032 = _18041 ^ _1669;
  wire _48033 = _8533 ^ _2435;
  wire _48034 = _48032 ^ _48033;
  wire _48035 = _48031 ^ _48034;
  wire _48036 = _48029 ^ _48035;
  wire _48037 = _20439 ^ uncoded_block[1716];
  wire _48038 = _48036 ^ _48037;
  wire _48039 = _48023 ^ _48038;
  wire _48040 = _47998 ^ _48039;
  wire _48041 = _47891 ^ _48040;
  wire _48042 = _3995 ^ _42204;
  wire _48043 = _39487 ^ _48042;
  wire _48044 = _13537 ^ _35096;
  wire _48045 = _9143 ^ _6095;
  wire _48046 = _48044 ^ _48045;
  wire _48047 = _48043 ^ _48046;
  wire _48048 = _4009 ^ _886;
  wire _48049 = _4722 ^ _48048;
  wire _48050 = _12996 ^ _9705;
  wire _48051 = _28765 ^ _6750;
  wire _48052 = _48050 ^ _48051;
  wire _48053 = _48049 ^ _48052;
  wire _48054 = _48047 ^ _48053;
  wire _48055 = _19980 ^ _15603;
  wire _48056 = _4026 ^ _14068;
  wire _48057 = _48055 ^ _48056;
  wire _48058 = _9718 ^ _15101;
  wire _48059 = uncoded_block[109] ^ uncoded_block[115];
  wire _48060 = _50 ^ _48059;
  wire _48061 = _48058 ^ _48060;
  wire _48062 = _48057 ^ _48061;
  wire _48063 = _33056 ^ _6771;
  wire _48064 = _48063 ^ _28448;
  wire _48065 = _6136 ^ _10830;
  wire _48066 = _5459 ^ _48065;
  wire _48067 = _48064 ^ _48066;
  wire _48068 = _48062 ^ _48067;
  wire _48069 = _48054 ^ _48068;
  wire _48070 = _67 ^ _932;
  wire _48071 = _1749 ^ _46182;
  wire _48072 = _48070 ^ _48071;
  wire _48073 = _2521 ^ _82;
  wire _48074 = _85 ^ _4062;
  wire _48075 = _48073 ^ _48074;
  wire _48076 = _48072 ^ _48075;
  wire _48077 = _947 ^ _3284;
  wire _48078 = _16116 ^ _10849;
  wire _48079 = _48077 ^ _48078;
  wire _48080 = _953 ^ _3296;
  wire _48081 = _14105 ^ _17617;
  wire _48082 = _48080 ^ _48081;
  wire _48083 = _48079 ^ _48082;
  wire _48084 = _48076 ^ _48083;
  wire _48085 = uncoded_block[237] ^ uncoded_block[242];
  wire _48086 = _10289 ^ _48085;
  wire _48087 = _38744 ^ _48086;
  wire _48088 = _4797 ^ _39154;
  wire _48089 = _48088 ^ _33934;
  wire _48090 = _48087 ^ _48089;
  wire _48091 = _23749 ^ _10871;
  wire _48092 = _4105 ^ _135;
  wire _48093 = _24211 ^ _48092;
  wire _48094 = _48091 ^ _48093;
  wire _48095 = _48090 ^ _48094;
  wire _48096 = _48084 ^ _48095;
  wire _48097 = _48069 ^ _48096;
  wire _48098 = _17142 ^ _1810;
  wire _48099 = _4111 ^ _31847;
  wire _48100 = _48098 ^ _48099;
  wire _48101 = _3340 ^ _149;
  wire _48102 = _41502 ^ _1014;
  wire _48103 = _48101 ^ _48102;
  wire _48104 = _48100 ^ _48103;
  wire _48105 = _2584 ^ _9240;
  wire _48106 = _48105 ^ _12525;
  wire _48107 = _4840 ^ _8652;
  wire _48108 = _4132 ^ _6863;
  wire _48109 = _48107 ^ _48108;
  wire _48110 = _48106 ^ _48109;
  wire _48111 = _48104 ^ _48110;
  wire _48112 = uncoded_block[362] ^ uncoded_block[367];
  wire _48113 = _48112 ^ _1838;
  wire _48114 = uncoded_block[373] ^ uncoded_block[380];
  wire _48115 = _48114 ^ _3377;
  wire _48116 = _48113 ^ _48115;
  wire _48117 = uncoded_block[387] ^ uncoded_block[393];
  wire _48118 = _3380 ^ _48117;
  wire _48119 = _6881 ^ _15696;
  wire _48120 = _48118 ^ _48119;
  wire _48121 = _48116 ^ _48120;
  wire _48122 = _183 ^ _4867;
  wire _48123 = _4868 ^ _9812;
  wire _48124 = _48122 ^ _48123;
  wire _48125 = _11479 ^ _14163;
  wire _48126 = _6254 ^ _28103;
  wire _48127 = _48125 ^ _48126;
  wire _48128 = _48124 ^ _48127;
  wire _48129 = _48121 ^ _48128;
  wire _48130 = _48111 ^ _48129;
  wire _48131 = _5578 ^ _1864;
  wire _48132 = _48131 ^ _26496;
  wire _48133 = _10926 ^ _9281;
  wire _48134 = _1079 ^ _1878;
  wire _48135 = _48133 ^ _48134;
  wire _48136 = _48132 ^ _48135;
  wire _48137 = _222 ^ _8694;
  wire _48138 = _19127 ^ _48137;
  wire _48139 = _24727 ^ _6919;
  wire _48140 = _7521 ^ _13674;
  wire _48141 = _48139 ^ _48140;
  wire _48142 = _48138 ^ _48141;
  wire _48143 = _48136 ^ _48142;
  wire _48144 = _8705 ^ _23370;
  wire _48145 = _48144 ^ _41142;
  wire _48146 = _4922 ^ _240;
  wire _48147 = _46254 ^ _48146;
  wire _48148 = _48145 ^ _48147;
  wire _48149 = _1905 ^ _14197;
  wire _48150 = _48149 ^ _24740;
  wire _48151 = uncoded_block[547] ^ uncoded_block[552];
  wire _48152 = uncoded_block[553] ^ uncoded_block[558];
  wire _48153 = _48151 ^ _48152;
  wire _48154 = uncoded_block[566] ^ uncoded_block[572];
  wire _48155 = _8725 ^ _48154;
  wire _48156 = _48153 ^ _48155;
  wire _48157 = _48150 ^ _48156;
  wire _48158 = _48148 ^ _48157;
  wire _48159 = _48143 ^ _48158;
  wire _48160 = _48130 ^ _48159;
  wire _48161 = _48097 ^ _48160;
  wire _48162 = _1931 ^ _15747;
  wire _48163 = _4946 ^ _31915;
  wire _48164 = _48162 ^ _48163;
  wire _48165 = _9330 ^ _1939;
  wire _48166 = _14737 ^ _277;
  wire _48167 = _48165 ^ _48166;
  wire _48168 = _48164 ^ _48167;
  wire _48169 = _278 ^ _4242;
  wire _48170 = _7564 ^ _3495;
  wire _48171 = _48169 ^ _48170;
  wire _48172 = _15261 ^ _7576;
  wire _48173 = _48172 ^ _46666;
  wire _48174 = _48171 ^ _48173;
  wire _48175 = _48168 ^ _48174;
  wire _48176 = _28908 ^ _304;
  wire _48177 = _21109 ^ _48176;
  wire _48178 = _3513 ^ _4262;
  wire _48179 = _28915 ^ _16752;
  wire _48180 = _48178 ^ _48179;
  wire _48181 = _48177 ^ _48180;
  wire _48182 = _2750 ^ _2754;
  wire _48183 = _47798 ^ _48182;
  wire _48184 = _4272 ^ _2757;
  wire _48185 = uncoded_block[704] ^ uncoded_block[711];
  wire _48186 = _14250 ^ _48185;
  wire _48187 = _48184 ^ _48186;
  wire _48188 = _48183 ^ _48187;
  wire _48189 = _48181 ^ _48188;
  wire _48190 = _48175 ^ _48189;
  wire _48191 = _28171 ^ _342;
  wire _48192 = _5691 ^ _7603;
  wire _48193 = _15788 ^ _350;
  wire _48194 = _48192 ^ _48193;
  wire _48195 = _48191 ^ _48194;
  wire _48196 = _5010 ^ _1999;
  wire _48197 = _1210 ^ _2778;
  wire _48198 = _48196 ^ _48197;
  wire _48199 = _2784 ^ _1221;
  wire _48200 = _25230 ^ _48199;
  wire _48201 = _48198 ^ _48200;
  wire _48202 = _48195 ^ _48201;
  wire _48203 = _25694 ^ _4311;
  wire _48204 = _14279 ^ _48203;
  wire _48205 = _19222 ^ _1233;
  wire _48206 = _383 ^ _5039;
  wire _48207 = _48205 ^ _48206;
  wire _48208 = _48204 ^ _48207;
  wire _48209 = _10485 ^ _5046;
  wire _48210 = _34063 ^ _48209;
  wire _48211 = _45332 ^ _3587;
  wire _48212 = uncoded_block[825] ^ uncoded_block[836];
  wire _48213 = _48212 ^ _14809;
  wire _48214 = _48211 ^ _48213;
  wire _48215 = _48210 ^ _48214;
  wire _48216 = _48208 ^ _48215;
  wire _48217 = _48202 ^ _48216;
  wire _48218 = _48190 ^ _48217;
  wire _48219 = _2820 ^ _8809;
  wire _48220 = _32395 ^ _48219;
  wire _48221 = _2046 ^ _408;
  wire _48222 = _13244 ^ _1266;
  wire _48223 = _48221 ^ _48222;
  wire _48224 = _48220 ^ _48223;
  wire _48225 = _12150 ^ _4347;
  wire _48226 = _5753 ^ _17811;
  wire _48227 = _48225 ^ _48226;
  wire _48228 = _25262 ^ _1280;
  wire _48229 = _2070 ^ _5092;
  wire _48230 = _48228 ^ _48229;
  wire _48231 = _48227 ^ _48230;
  wire _48232 = _48224 ^ _48231;
  wire _48233 = _12714 ^ _2857;
  wire _48234 = _48233 ^ _44220;
  wire _48235 = _4377 ^ _1302;
  wire _48236 = _14326 ^ _4382;
  wire _48237 = _48235 ^ _48236;
  wire _48238 = _48234 ^ _48237;
  wire _48239 = _35692 ^ _12179;
  wire _48240 = _7682 ^ _8847;
  wire _48241 = _48239 ^ _48240;
  wire _48242 = _5112 ^ _471;
  wire _48243 = _10537 ^ _2102;
  wire _48244 = _48242 ^ _48243;
  wire _48245 = _48241 ^ _48244;
  wire _48246 = _48238 ^ _48245;
  wire _48247 = _48232 ^ _48246;
  wire _48248 = _1318 ^ _2883;
  wire _48249 = _7691 ^ _38929;
  wire _48250 = _48248 ^ _48249;
  wire _48251 = _1327 ^ _2890;
  wire _48252 = _2118 ^ _2894;
  wire _48253 = _48251 ^ _48252;
  wire _48254 = _48250 ^ _48253;
  wire _48255 = uncoded_block[1028] ^ uncoded_block[1036];
  wire _48256 = _8872 ^ _48255;
  wire _48257 = uncoded_block[1037] ^ uncoded_block[1043];
  wire _48258 = _48257 ^ _46364;
  wire _48259 = _48256 ^ _48258;
  wire _48260 = _17858 ^ _23502;
  wire _48261 = _48259 ^ _48260;
  wire _48262 = _48254 ^ _48261;
  wire _48263 = _3689 ^ _2924;
  wire _48264 = _20251 ^ _42054;
  wire _48265 = _48263 ^ _48264;
  wire _48266 = _20253 ^ _5840;
  wire _48267 = uncoded_block[1101] ^ uncoded_block[1109];
  wire _48268 = _33305 ^ _48267;
  wire _48269 = _48266 ^ _48268;
  wire _48270 = _48265 ^ _48269;
  wire _48271 = _552 ^ _1388;
  wire _48272 = _10587 ^ _33312;
  wire _48273 = _48271 ^ _48272;
  wire _48274 = _35343 ^ _2953;
  wire _48275 = _26234 ^ _48274;
  wire _48276 = _48273 ^ _48275;
  wire _48277 = _48270 ^ _48276;
  wire _48278 = _48262 ^ _48277;
  wire _48279 = _48247 ^ _48278;
  wire _48280 = _48218 ^ _48279;
  wire _48281 = _48161 ^ _48280;
  wire _48282 = _10597 ^ _27532;
  wire _48283 = _48282 ^ _5189;
  wire _48284 = _3733 ^ _22627;
  wire _48285 = uncoded_block[1166] ^ uncoded_block[1171];
  wire _48286 = _6511 ^ _48285;
  wire _48287 = _48284 ^ _48286;
  wire _48288 = _48283 ^ _48287;
  wire _48289 = _32064 ^ _2193;
  wire _48290 = _6520 ^ _13883;
  wire _48291 = _48289 ^ _48290;
  wire _48292 = _12810 ^ _18389;
  wire _48293 = _36576 ^ _48292;
  wire _48294 = _48291 ^ _48293;
  wire _48295 = _48288 ^ _48294;
  wire _48296 = uncoded_block[1204] ^ uncoded_block[1210];
  wire _48297 = _48296 ^ _26694;
  wire _48298 = _12813 ^ _2220;
  wire _48299 = _48297 ^ _48298;
  wire _48300 = _610 ^ _16407;
  wire _48301 = _48299 ^ _48300;
  wire _48302 = _43141 ^ _31231;
  wire _48303 = _17911 ^ _6543;
  wire _48304 = _48302 ^ _48303;
  wire _48305 = _20801 ^ _34563;
  wire _48306 = _7779 ^ _48305;
  wire _48307 = _48304 ^ _48306;
  wire _48308 = _48301 ^ _48307;
  wire _48309 = _48295 ^ _48308;
  wire _48310 = _4523 ^ _1463;
  wire _48311 = _28656 ^ _48310;
  wire _48312 = _3794 ^ _26271;
  wire _48313 = _29913 ^ _4531;
  wire _48314 = _48312 ^ _48313;
  wire _48315 = _48311 ^ _48314;
  wire _48316 = _8984 ^ _23131;
  wire _48317 = _26276 ^ _2262;
  wire _48318 = _48316 ^ _48317;
  wire _48319 = uncoded_block[1318] ^ uncoded_block[1325];
  wire _48320 = _48319 ^ _657;
  wire _48321 = _48320 ^ _3035;
  wire _48322 = _48318 ^ _48321;
  wire _48323 = _48315 ^ _48322;
  wire _48324 = _13399 ^ _10092;
  wire _48325 = _17938 ^ _5268;
  wire _48326 = _48324 ^ _48325;
  wire _48327 = _21303 ^ _6587;
  wire _48328 = _48327 ^ _35396;
  wire _48329 = _48326 ^ _48328;
  wire _48330 = _6594 ^ _7824;
  wire _48331 = _21763 ^ _48330;
  wire _48332 = _22687 ^ _11782;
  wire _48333 = _2293 ^ _4569;
  wire _48334 = _48332 ^ _48333;
  wire _48335 = _48331 ^ _48334;
  wire _48336 = _48329 ^ _48335;
  wire _48337 = _48323 ^ _48336;
  wire _48338 = _48309 ^ _48337;
  wire _48339 = _4571 ^ _29090;
  wire _48340 = _4578 ^ _701;
  wire _48341 = _48339 ^ _48340;
  wire _48342 = _3853 ^ _32948;
  wire _48343 = _21783 ^ _2318;
  wire _48344 = _48342 ^ _48343;
  wire _48345 = _48341 ^ _48344;
  wire _48346 = uncoded_block[1444] ^ uncoded_block[1447];
  wire _48347 = _4590 ^ _48346;
  wire _48348 = _3865 ^ _726;
  wire _48349 = _48347 ^ _48348;
  wire _48350 = _16977 ^ _41757;
  wire _48351 = _47599 ^ _48350;
  wire _48352 = _48349 ^ _48351;
  wire _48353 = _48345 ^ _48352;
  wire _48354 = _12342 ^ _10706;
  wire _48355 = _48354 ^ _46464;
  wire _48356 = _3890 ^ _11260;
  wire _48357 = _1571 ^ _7262;
  wire _48358 = _48356 ^ _48357;
  wire _48359 = _48355 ^ _48358;
  wire _48360 = _15002 ^ _9055;
  wire _48361 = _27621 ^ _2357;
  wire _48362 = _48360 ^ _48361;
  wire _48363 = _27193 ^ _21349;
  wire _48364 = _48362 ^ _48363;
  wire _48365 = _48359 ^ _48364;
  wire _48366 = _48353 ^ _48365;
  wire _48367 = _15009 ^ _1589;
  wire _48368 = _1590 ^ _18492;
  wire _48369 = _48367 ^ _48368;
  wire _48370 = _43217 ^ _3914;
  wire _48371 = _48370 ^ _30440;
  wire _48372 = _48369 ^ _48371;
  wire _48373 = _24102 ^ _15026;
  wire _48374 = _10163 ^ _1609;
  wire _48375 = _48373 ^ _48374;
  wire _48376 = _46487 ^ _5368;
  wire _48377 = _48376 ^ _23646;
  wire _48378 = _48375 ^ _48377;
  wire _48379 = _48372 ^ _48378;
  wire _48380 = _8499 ^ _5373;
  wire _48381 = _48380 ^ _35452;
  wire _48382 = _16031 ^ _18020;
  wire _48383 = _7912 ^ _807;
  wire _48384 = _48382 ^ _48383;
  wire _48385 = _48381 ^ _48384;
  wire _48386 = _1639 ^ _18965;
  wire _48387 = _7309 ^ _2411;
  wire _48388 = _48386 ^ _48387;
  wire _48389 = _6054 ^ _25024;
  wire _48390 = _48388 ^ _48389;
  wire _48391 = _48385 ^ _48390;
  wire _48392 = _48379 ^ _48391;
  wire _48393 = _48366 ^ _48392;
  wire _48394 = _48338 ^ _48393;
  wire _48395 = _10196 ^ _22303;
  wire _48396 = _19939 ^ _17538;
  wire _48397 = _48395 ^ _48396;
  wire _48398 = _6061 ^ _14543;
  wire _48399 = _48398 ^ _3191;
  wire _48400 = _48397 ^ _48399;
  wire _48401 = _6066 ^ _9677;
  wire _48402 = _48401 ^ _20919;
  wire _48403 = uncoded_block[1702] ^ uncoded_block[1707];
  wire _48404 = _48403 ^ _12407;
  wire _48405 = _48404 ^ _856;
  wire _48406 = _48402 ^ _48405;
  wire _48407 = _48400 ^ _48406;
  wire _48408 = _48407 ^ uncoded_block[1719];
  wire _48409 = _48394 ^ _48408;
  wire _48410 = _48281 ^ _48409;
  wire _48411 = _19959 ^ _42204;
  wire _48412 = _37908 ^ _48411;
  wire _48413 = _7351 ^ _4001;
  wire _48414 = uncoded_block[35] ^ uncoded_block[40];
  wire _48415 = _48414 ^ _20457;
  wire _48416 = _48413 ^ _48415;
  wire _48417 = _48412 ^ _48416;
  wire _48418 = uncoded_block[48] ^ uncoded_block[54];
  wire _48419 = _12425 ^ _48418;
  wire _48420 = _16572 ^ _20465;
  wire _48421 = _48419 ^ _48420;
  wire _48422 = _2474 ^ _34289;
  wire _48423 = _11357 ^ _897;
  wire _48424 = _48422 ^ _48423;
  wire _48425 = _48421 ^ _48424;
  wire _48426 = _48417 ^ _48425;
  wire _48427 = _46927 ^ _45162;
  wire _48428 = _4739 ^ _16584;
  wire _48429 = _48428 ^ _15608;
  wire _48430 = _48427 ^ _48429;
  wire _48431 = _9166 ^ _20957;
  wire _48432 = uncoded_block[116] ^ uncoded_block[120];
  wire _48433 = _48432 ^ _10821;
  wire _48434 = _48431 ^ _48433;
  wire _48435 = _13017 ^ _1735;
  wire _48436 = _15112 ^ _1736;
  wire _48437 = _48435 ^ _48436;
  wire _48438 = _48434 ^ _48437;
  wire _48439 = _48430 ^ _48438;
  wire _48440 = _48426 ^ _48439;
  wire _48441 = _6136 ^ _1742;
  wire _48442 = _8000 ^ _71;
  wire _48443 = _48441 ^ _48442;
  wire _48444 = _73 ^ _6144;
  wire _48445 = _1749 ^ _81;
  wire _48446 = _48444 ^ _48445;
  wire _48447 = _48443 ^ _48446;
  wire _48448 = _5477 ^ _2525;
  wire _48449 = _15631 ^ _3284;
  wire _48450 = _48448 ^ _48449;
  wire _48451 = uncoded_block[198] ^ uncoded_block[203];
  wire _48452 = _48451 ^ _97;
  wire _48453 = _3292 ^ _17116;
  wire _48454 = _48452 ^ _48453;
  wire _48455 = _48450 ^ _48454;
  wire _48456 = _48447 ^ _48455;
  wire _48457 = _1774 ^ _23300;
  wire _48458 = _37159 ^ _48457;
  wire _48459 = uncoded_block[239] ^ uncoded_block[244];
  wire _48460 = _970 ^ _48459;
  wire _48461 = _16626 ^ _13053;
  wire _48462 = _48460 ^ _48461;
  wire _48463 = _48458 ^ _48462;
  wire _48464 = uncoded_block[265] ^ uncoded_block[270];
  wire _48465 = _10297 ^ _48464;
  wire _48466 = _38753 ^ _48465;
  wire _48467 = _12506 ^ _8632;
  wire _48468 = _18607 ^ _48467;
  wire _48469 = _48466 ^ _48468;
  wire _48470 = _48463 ^ _48469;
  wire _48471 = _48456 ^ _48470;
  wire _48472 = _48440 ^ _48471;
  wire _48473 = _19574 ^ _3332;
  wire _48474 = _48473 ^ _20537;
  wire _48475 = _15168 ^ _6208;
  wire _48476 = uncoded_block[321] ^ uncoded_block[326];
  wire _48477 = _48476 ^ _8063;
  wire _48478 = _48475 ^ _48477;
  wire _48479 = _48474 ^ _48478;
  wire _48480 = _15173 ^ _6217;
  wire _48481 = _48480 ^ _11452;
  wire _48482 = _2599 ^ _11455;
  wire _48483 = _20554 ^ _12530;
  wire _48484 = _48482 ^ _48483;
  wire _48485 = _48481 ^ _48484;
  wire _48486 = _48479 ^ _48485;
  wire _48487 = _26032 ^ _16662;
  wire _48488 = uncoded_block[373] ^ uncoded_block[378];
  wire _48489 = _1838 ^ _48488;
  wire _48490 = _48487 ^ _48489;
  wire _48491 = _28090 ^ _13102;
  wire _48492 = _3383 ^ _10910;
  wire _48493 = _48491 ^ _48492;
  wire _48494 = _48490 ^ _48493;
  wire _48495 = _1048 ^ _41525;
  wire _48496 = _11473 ^ _21508;
  wire _48497 = _48495 ^ _48496;
  wire _48498 = _19613 ^ _14160;
  wire _48499 = uncoded_block[425] ^ uncoded_block[428];
  wire _48500 = _48499 ^ _32297;
  wire _48501 = _48498 ^ _48500;
  wire _48502 = _48497 ^ _48501;
  wire _48503 = _48494 ^ _48502;
  wire _48504 = _48486 ^ _48503;
  wire _48505 = _17181 ^ _9275;
  wire _48506 = _42297 ^ _48505;
  wire _48507 = uncoded_block[447] ^ uncoded_block[452];
  wire _48508 = _48507 ^ _1075;
  wire _48509 = _48508 ^ _5585;
  wire _48510 = _48506 ^ _48509;
  wire _48511 = _21058 ^ _48134;
  wire _48512 = uncoded_block[472] ^ uncoded_block[478];
  wire _48513 = _3418 ^ _48512;
  wire _48514 = _5598 ^ _7516;
  wire _48515 = _48513 ^ _48514;
  wire _48516 = _48511 ^ _48515;
  wire _48517 = _48510 ^ _48516;
  wire _48518 = _43357 ^ _228;
  wire _48519 = _48518 ^ _37227;
  wire _48520 = _9294 ^ _3439;
  wire _48521 = uncoded_block[514] ^ uncoded_block[524];
  wire _48522 = _48521 ^ _1900;
  wire _48523 = _48520 ^ _48522;
  wire _48524 = _48519 ^ _48523;
  wire _48525 = _6929 ^ _21550;
  wire _48526 = _48525 ^ _38410;
  wire _48527 = _4937 ^ _5633;
  wire _48528 = _22005 ^ _48527;
  wire _48529 = _48526 ^ _48528;
  wire _48530 = _48524 ^ _48529;
  wire _48531 = _48517 ^ _48530;
  wire _48532 = _48504 ^ _48531;
  wire _48533 = _48472 ^ _48532;
  wire _48534 = _6942 ^ _4224;
  wire _48535 = _40404 ^ _48534;
  wire _48536 = _4941 ^ _19652;
  wire _48537 = _31915 ^ _3478;
  wire _48538 = _48536 ^ _48537;
  wire _48539 = _48535 ^ _48538;
  wire _48540 = _2700 ^ _4236;
  wire _48541 = _8149 ^ _1142;
  wire _48542 = _48540 ^ _48541;
  wire _48543 = _5646 ^ _1146;
  wire _48544 = _48543 ^ _14222;
  wire _48545 = _48542 ^ _48544;
  wire _48546 = _48539 ^ _48545;
  wire _48547 = _13713 ^ _31060;
  wire _48548 = _28901 ^ _11543;
  wire _48549 = _48547 ^ _48548;
  wire _48550 = _4255 ^ _12624;
  wire _48551 = _48550 ^ _21579;
  wire _48552 = _48549 ^ _48551;
  wire _48553 = uncoded_block[661] ^ uncoded_block[664];
  wire _48554 = _40030 ^ _48553;
  wire _48555 = _4264 ^ _311;
  wire _48556 = _48554 ^ _48555;
  wire _48557 = _8176 ^ _6349;
  wire _48558 = _48557 ^ _14245;
  wire _48559 = _48556 ^ _48558;
  wire _48560 = _48552 ^ _48559;
  wire _48561 = _48546 ^ _48560;
  wire _48562 = _3527 ^ _326;
  wire _48563 = _6358 ^ _3529;
  wire _48564 = _48562 ^ _48563;
  wire _48565 = _4989 ^ _14250;
  wire _48566 = _48565 ^ _18256;
  wire _48567 = _48564 ^ _48566;
  wire _48568 = _31946 ^ _1196;
  wire _48569 = _4286 ^ _18730;
  wire _48570 = _31527 ^ _48569;
  wire _48571 = _48568 ^ _48570;
  wire _48572 = _48567 ^ _48571;
  wire _48573 = uncoded_block[737] ^ uncoded_block[742];
  wire _48574 = _48573 ^ _5012;
  wire _48575 = _8778 ^ _1214;
  wire _48576 = _48574 ^ _48575;
  wire _48577 = _5017 ^ _3559;
  wire _48578 = _48577 ^ _13763;
  wire _48579 = _48576 ^ _48578;
  wire _48580 = _17776 ^ _11019;
  wire _48581 = _48580 ^ _25690;
  wire _48582 = _17284 ^ _2015;
  wire _48583 = _1224 ^ _10475;
  wire _48584 = _48582 ^ _48583;
  wire _48585 = _48581 ^ _48584;
  wire _48586 = _48579 ^ _48585;
  wire _48587 = _48572 ^ _48586;
  wire _48588 = _48561 ^ _48587;
  wire _48589 = _375 ^ _382;
  wire _48590 = _48589 ^ _30669;
  wire _48591 = _389 ^ _1238;
  wire _48592 = _48591 ^ _8229;
  wire _48593 = _48590 ^ _48592;
  wire _48594 = _11597 ^ _5051;
  wire _48595 = _17793 ^ _2033;
  wire _48596 = _48594 ^ _48595;
  wire _48597 = _401 ^ _5058;
  wire _48598 = _11609 ^ _7643;
  wire _48599 = _48597 ^ _48598;
  wire _48600 = _48596 ^ _48599;
  wire _48601 = _48593 ^ _48600;
  wire _48602 = _8237 ^ _2047;
  wire _48603 = _9948 ^ _27452;
  wire _48604 = _48602 ^ _48603;
  wire _48605 = _12150 ^ _16815;
  wire _48606 = _8820 ^ _2058;
  wire _48607 = _48605 ^ _48606;
  wire _48608 = _48604 ^ _48607;
  wire _48609 = uncoded_block[898] ^ uncoded_block[902];
  wire _48610 = _48609 ^ _2065;
  wire _48611 = _4356 ^ _48610;
  wire _48612 = _431 ^ _2070;
  wire _48613 = _3628 ^ _18775;
  wire _48614 = _48612 ^ _48613;
  wire _48615 = _48611 ^ _48614;
  wire _48616 = _48608 ^ _48615;
  wire _48617 = _48601 ^ _48616;
  wire _48618 = uncoded_block[927] ^ uncoded_block[935];
  wire _48619 = _48618 ^ _2083;
  wire _48620 = _2856 ^ _48619;
  wire _48621 = uncoded_block[943] ^ uncoded_block[947];
  wire _48622 = _6439 ^ _48621;
  wire _48623 = _48622 ^ _4383;
  wire _48624 = _48620 ^ _48623;
  wire _48625 = _1307 ^ _7680;
  wire _48626 = _48625 ^ _23033;
  wire _48627 = _3657 ^ _3659;
  wire _48628 = _29828 ^ _48627;
  wire _48629 = _48626 ^ _48628;
  wire _48630 = _48624 ^ _48629;
  wire _48631 = _5118 ^ _19275;
  wire _48632 = _5798 ^ _24858;
  wire _48633 = _48631 ^ _48632;
  wire _48634 = _4409 ^ _4412;
  wire _48635 = uncoded_block[1020] ^ uncoded_block[1026];
  wire _48636 = _8871 ^ _48635;
  wire _48637 = _48634 ^ _48636;
  wire _48638 = _48633 ^ _48637;
  wire _48639 = _11668 ^ _1342;
  wire _48640 = _34924 ^ _48639;
  wire _48641 = uncoded_block[1038] ^ uncoded_block[1042];
  wire _48642 = _48641 ^ _514;
  wire _48643 = _3681 ^ _2136;
  wire _48644 = _48642 ^ _48643;
  wire _48645 = _48640 ^ _48644;
  wire _48646 = _48638 ^ _48645;
  wire _48647 = _48630 ^ _48646;
  wire _48648 = _48617 ^ _48647;
  wire _48649 = _48588 ^ _48648;
  wire _48650 = _48533 ^ _48649;
  wire _48651 = _1359 ^ _11120;
  wire _48652 = uncoded_block[1061] ^ uncoded_block[1067];
  wire _48653 = _48652 ^ _5158;
  wire _48654 = _48651 ^ _48653;
  wire _48655 = _25774 ^ _7724;
  wire _48656 = _7725 ^ _536;
  wire _48657 = _48655 ^ _48656;
  wire _48658 = _48654 ^ _48657;
  wire _48659 = _537 ^ _42741;
  wire _48660 = _48659 ^ _40138;
  wire _48661 = _14882 ^ _12782;
  wire _48662 = _48661 ^ _8921;
  wire _48663 = _48660 ^ _48662;
  wire _48664 = _48658 ^ _48663;
  wire _48665 = _2942 ^ _20265;
  wire _48666 = _15896 ^ _20266;
  wire _48667 = _48665 ^ _48666;
  wire _48668 = _5859 ^ _7141;
  wire _48669 = _48668 ^ _2187;
  wire _48670 = _48667 ^ _48669;
  wire _48671 = _19330 ^ _23532;
  wire _48672 = _43884 ^ _6519;
  wire _48673 = _48671 ^ _48672;
  wire _48674 = uncoded_block[1181] ^ uncoded_block[1185];
  wire _48675 = _48674 ^ _2971;
  wire _48676 = _38970 ^ _7160;
  wire _48677 = _48675 ^ _48676;
  wire _48678 = _48673 ^ _48677;
  wire _48679 = _48670 ^ _48678;
  wire _48680 = _48664 ^ _48679;
  wire _48681 = _8370 ^ _1425;
  wire _48682 = _23544 ^ _2982;
  wire _48683 = _48681 ^ _48682;
  wire _48684 = _10620 ^ _10059;
  wire _48685 = _7168 ^ _612;
  wire _48686 = _48684 ^ _48685;
  wire _48687 = _48683 ^ _48686;
  wire _48688 = _18400 ^ _5219;
  wire _48689 = uncoded_block[1238] ^ uncoded_block[1247];
  wire _48690 = _48689 ^ _6543;
  wire _48691 = _48688 ^ _48690;
  wire _48692 = _19358 ^ _1455;
  wire _48693 = _3003 ^ _6550;
  wire _48694 = _48692 ^ _48693;
  wire _48695 = _48691 ^ _48694;
  wire _48696 = _48687 ^ _48695;
  wire _48697 = _3008 ^ _6554;
  wire _48698 = _16419 ^ _10638;
  wire _48699 = _48697 ^ _48698;
  wire _48700 = _10077 ^ _13380;
  wire _48701 = _48700 ^ _1470;
  wire _48702 = _48699 ^ _48701;
  wire _48703 = _6563 ^ _20812;
  wire _48704 = _48703 ^ _26727;
  wire _48705 = _1490 ^ _22672;
  wire _48706 = _3030 ^ _48705;
  wire _48707 = _48704 ^ _48706;
  wire _48708 = _48702 ^ _48707;
  wire _48709 = _48696 ^ _48708;
  wire _48710 = _48680 ^ _48709;
  wire _48711 = uncoded_block[1357] ^ uncoded_block[1361];
  wire _48712 = _5272 ^ _48711;
  wire _48713 = _13407 ^ _24954;
  wire _48714 = _48712 ^ _48713;
  wire _48715 = _45452 ^ _48714;
  wire _48716 = _12866 ^ _19861;
  wire _48717 = _48716 ^ _15968;
  wire _48718 = _21774 ^ _26747;
  wire _48719 = _5293 ^ _9585;
  wire _48720 = _48718 ^ _48719;
  wire _48721 = _48717 ^ _48720;
  wire _48722 = _48715 ^ _48721;
  wire _48723 = _17461 ^ _14466;
  wire _48724 = _15980 ^ _8443;
  wire _48725 = _48723 ^ _48724;
  wire _48726 = _17470 ^ _5304;
  wire _48727 = _716 ^ _1543;
  wire _48728 = _48726 ^ _48727;
  wire _48729 = _48725 ^ _48728;
  wire _48730 = _18470 ^ _3881;
  wire _48731 = _6626 ^ _48730;
  wire _48732 = _736 ^ _3101;
  wire _48733 = _739 ^ _16981;
  wire _48734 = _48732 ^ _48733;
  wire _48735 = _48731 ^ _48734;
  wire _48736 = _48729 ^ _48735;
  wire _48737 = _48722 ^ _48736;
  wire _48738 = _16483 ^ _7257;
  wire _48739 = _1573 ^ _43960;
  wire _48740 = _48738 ^ _48739;
  wire _48741 = _19897 ^ _8473;
  wire _48742 = _34222 ^ _48741;
  wire _48743 = _11272 ^ _13979;
  wire _48744 = _3908 ^ _1589;
  wire _48745 = _48743 ^ _48744;
  wire _48746 = _48742 ^ _48745;
  wire _48747 = _48740 ^ _48746;
  wire _48748 = uncoded_block[1556] ^ uncoded_block[1560];
  wire _48749 = _43217 ^ _48748;
  wire _48750 = _31729 ^ _48749;
  wire _48751 = _2372 ^ _37871;
  wire _48752 = _7285 ^ _47625;
  wire _48753 = _48751 ^ _48752;
  wire _48754 = _48750 ^ _48753;
  wire _48755 = _22284 ^ _24566;
  wire _48756 = _8500 ^ _2396;
  wire _48757 = _3157 ^ _804;
  wire _48758 = _48756 ^ _48757;
  wire _48759 = _48755 ^ _48758;
  wire _48760 = _48754 ^ _48759;
  wire _48761 = _48747 ^ _48760;
  wire _48762 = _48737 ^ _48761;
  wire _48763 = _48710 ^ _48762;
  wire _48764 = _7298 ^ _7300;
  wire _48765 = uncoded_block[1627] ^ uncoded_block[1634];
  wire _48766 = _6046 ^ _48765;
  wire _48767 = _48764 ^ _48766;
  wire _48768 = _3949 ^ _23223;
  wire _48769 = _48767 ^ _48768;
  wire _48770 = _18030 ^ _14011;
  wire _48771 = uncoded_block[1662] ^ uncoded_block[1666];
  wire _48772 = _48771 ^ _3182;
  wire _48773 = _48770 ^ _48772;
  wire _48774 = uncoded_block[1674] ^ uncoded_block[1678];
  wire _48775 = _6700 ^ _48774;
  wire _48776 = _48775 ^ _26829;
  wire _48777 = _48773 ^ _48776;
  wire _48778 = _48769 ^ _48777;
  wire _48779 = _6066 ^ _3972;
  wire _48780 = _5409 ^ _9120;
  wire _48781 = _48779 ^ _48780;
  wire _48782 = _3976 ^ _3979;
  wire _48783 = _2438 ^ _26369;
  wire _48784 = _48782 ^ _48783;
  wire _48785 = _48781 ^ _48784;
  wire _48786 = _48785 ^ _17554;
  wire _48787 = _48778 ^ _48786;
  wire _48788 = _48763 ^ _48787;
  wire _48789 = _48650 ^ _48788;
  wire _48790 = _7347 ^ _3995;
  wire _48791 = _7 ^ _46150;
  wire _48792 = _48790 ^ _48791;
  wire _48793 = _11344 ^ _3227;
  wire _48794 = _36711 ^ _48793;
  wire _48795 = _48792 ^ _48794;
  wire _48796 = _18 ^ _20457;
  wire _48797 = _3232 ^ _8556;
  wire _48798 = _48796 ^ _48797;
  wire _48799 = _12996 ^ _13553;
  wire _48800 = uncoded_block[70] ^ uncoded_block[75];
  wire _48801 = _34 ^ _48800;
  wire _48802 = _48799 ^ _48801;
  wire _48803 = _48798 ^ _48802;
  wire _48804 = _48795 ^ _48803;
  wire _48805 = _20472 ^ _7981;
  wire _48806 = _23704 ^ _48805;
  wire _48807 = _4026 ^ _3249;
  wire _48808 = _48807 ^ _31798;
  wire _48809 = _48806 ^ _48808;
  wire _48810 = uncoded_block[105] ^ uncoded_block[109];
  wire _48811 = _48810 ^ _7990;
  wire _48812 = _48432 ^ _13016;
  wire _48813 = _48811 ^ _48812;
  wire _48814 = uncoded_block[132] ^ uncoded_block[138];
  wire _48815 = _48814 ^ _4043;
  wire _48816 = _1734 ^ _48815;
  wire _48817 = _48813 ^ _48816;
  wire _48818 = _48809 ^ _48817;
  wire _48819 = _48804 ^ _48818;
  wire _48820 = _17097 ^ _7397;
  wire _48821 = _48820 ^ _19535;
  wire _48822 = _30519 ^ _8591;
  wire _48823 = uncoded_block[172] ^ uncoded_block[178];
  wire _48824 = _48823 ^ _8009;
  wire _48825 = _48822 ^ _48824;
  wire _48826 = _48821 ^ _48825;
  wire _48827 = _4772 ^ _3283;
  wire _48828 = _4777 ^ _14099;
  wire _48829 = _48827 ^ _48828;
  wire _48830 = uncoded_block[215] ^ uncoded_block[224];
  wire _48831 = _33082 ^ _48830;
  wire _48832 = uncoded_block[225] ^ uncoded_block[232];
  wire _48833 = _48832 ^ _2550;
  wire _48834 = _48831 ^ _48833;
  wire _48835 = _48829 ^ _48834;
  wire _48836 = _48826 ^ _48835;
  wire _48837 = _7423 ^ _16622;
  wire _48838 = _48837 ^ _26433;
  wire _48839 = _116 ^ _31834;
  wire _48840 = _8041 ^ _22855;
  wire _48841 = _48839 ^ _48840;
  wire _48842 = _48838 ^ _48841;
  wire _48843 = _4102 ^ _26895;
  wire _48844 = _20524 ^ _48843;
  wire _48845 = uncoded_block[285] ^ uncoded_block[290];
  wire _48846 = _4105 ^ _48845;
  wire _48847 = _11968 ^ _48846;
  wire _48848 = _48844 ^ _48847;
  wire _48849 = _48842 ^ _48848;
  wire _48850 = _48836 ^ _48849;
  wire _48851 = _48819 ^ _48850;
  wire _48852 = _19076 ^ _33529;
  wire _48853 = _3338 ^ _3340;
  wire _48854 = _1008 ^ _2583;
  wire _48855 = _48853 ^ _48854;
  wire _48856 = _48852 ^ _48855;
  wire _48857 = _16153 ^ _24225;
  wire _48858 = _30994 ^ _34356;
  wire _48859 = _48857 ^ _48858;
  wire _48860 = _48856 ^ _48859;
  wire _48861 = _2602 ^ _21030;
  wire _48862 = _48861 ^ _37596;
  wire _48863 = _13101 ^ _10907;
  wire _48864 = _10896 ^ _48863;
  wire _48865 = _48862 ^ _48864;
  wire _48866 = _5554 ^ _8661;
  wire _48867 = _48866 ^ _6885;
  wire _48868 = uncoded_block[409] ^ uncoded_block[417];
  wire _48869 = _3391 ^ _48868;
  wire _48870 = uncoded_block[418] ^ uncoded_block[424];
  wire _48871 = _48870 ^ _1062;
  wire _48872 = _48869 ^ _48871;
  wire _48873 = _48867 ^ _48872;
  wire _48874 = _48865 ^ _48873;
  wire _48875 = _48860 ^ _48874;
  wire _48876 = _4169 ^ _5577;
  wire _48877 = _19616 ^ _48876;
  wire _48878 = _1864 ^ _33565;
  wire _48879 = _48878 ^ _13663;
  wire _48880 = _48877 ^ _48879;
  wire _48881 = _16691 ^ _43727;
  wire _48882 = _16693 ^ _5598;
  wire _48883 = _48882 ^ _36813;
  wire _48884 = _48881 ^ _48883;
  wire _48885 = _48880 ^ _48884;
  wire _48886 = _8117 ^ _4905;
  wire _48887 = _48886 ^ _48140;
  wire _48888 = _9295 ^ _4910;
  wire _48889 = _19638 ^ _1108;
  wire _48890 = _48888 ^ _48889;
  wire _48891 = _48887 ^ _48890;
  wire _48892 = _13684 ^ _1900;
  wire _48893 = _48892 ^ _24278;
  wire _48894 = _41554 ^ _1913;
  wire _48895 = _32727 ^ _48894;
  wire _48896 = _48893 ^ _48895;
  wire _48897 = _48891 ^ _48896;
  wire _48898 = _48885 ^ _48897;
  wire _48899 = _48875 ^ _48898;
  wire _48900 = _48851 ^ _48899;
  wire _48901 = _8138 ^ _43374;
  wire _48902 = _3468 ^ _10399;
  wire _48903 = _1133 ^ _1138;
  wire _48904 = _48902 ^ _48903;
  wire _48905 = _48901 ^ _48904;
  wire _48906 = _1938 ^ _37253;
  wire _48907 = _20117 ^ _48906;
  wire _48908 = _46272 ^ _22470;
  wire _48909 = _48907 ^ _48908;
  wire _48910 = _48905 ^ _48909;
  wire _48911 = _28147 ^ _7570;
  wire _48912 = _7565 ^ _48911;
  wire _48913 = _12075 ^ _1161;
  wire _48914 = _14746 ^ _48913;
  wire _48915 = _48912 ^ _48914;
  wire _48916 = _16241 ^ _2729;
  wire _48917 = _6338 ^ _25206;
  wire _48918 = _48916 ^ _48917;
  wire _48919 = _3514 ^ _3516;
  wire _48920 = _36021 ^ _48919;
  wire _48921 = _48918 ^ _48920;
  wire _48922 = _48915 ^ _48921;
  wire _48923 = _48910 ^ _48922;
  wire _48924 = _1971 ^ _6983;
  wire _48925 = _34032 ^ _48924;
  wire _48926 = _1974 ^ _22493;
  wire _48927 = _48926 ^ _15286;
  wire _48928 = _48925 ^ _48927;
  wire _48929 = uncoded_block[704] ^ uncoded_block[709];
  wire _48930 = _48929 ^ _2762;
  wire _48931 = _19201 ^ _2765;
  wire _48932 = _48930 ^ _48931;
  wire _48933 = uncoded_block[725] ^ uncoded_block[731];
  wire _48934 = _48933 ^ _1206;
  wire _48935 = _4289 ^ _353;
  wire _48936 = _48934 ^ _48935;
  wire _48937 = _48932 ^ _48936;
  wire _48938 = _48928 ^ _48937;
  wire _48939 = _14266 ^ _5017;
  wire _48940 = _3559 ^ _8781;
  wire _48941 = _48939 ^ _48940;
  wire _48942 = _4301 ^ _17776;
  wire _48943 = _48942 ^ _12668;
  wire _48944 = _48941 ^ _48943;
  wire _48945 = _41600 ^ _28189;
  wire _48946 = _3575 ^ _47086;
  wire _48947 = _48945 ^ _48946;
  wire _48948 = _48944 ^ _48947;
  wire _48949 = _48938 ^ _48948;
  wire _48950 = _48923 ^ _48949;
  wire _48951 = _20175 ^ _22523;
  wire _48952 = _5046 ^ _14290;
  wire _48953 = uncoded_block[824] ^ uncoded_block[827];
  wire _48954 = _48953 ^ _7039;
  wire _48955 = _48952 ^ _48954;
  wire _48956 = _48951 ^ _48955;
  wire _48957 = _47457 ^ _47095;
  wire _48958 = _3597 ^ _2820;
  wire _48959 = _11048 ^ _8812;
  wire _48960 = _48958 ^ _48959;
  wire _48961 = _48957 ^ _48960;
  wire _48962 = _48956 ^ _48961;
  wire _48963 = _5067 ^ _46331;
  wire _48964 = _20696 ^ _11056;
  wire _48965 = _22542 ^ _48964;
  wire _48966 = _48963 ^ _48965;
  wire _48967 = _11059 ^ _1273;
  wire _48968 = _48967 ^ _31573;
  wire _48969 = _5758 ^ _1278;
  wire _48970 = _48969 ^ _25728;
  wire _48971 = _48968 ^ _48970;
  wire _48972 = _48966 ^ _48971;
  wire _48973 = _48962 ^ _48972;
  wire _48974 = _44973 ^ _24833;
  wire _48975 = _2076 ^ _16827;
  wire _48976 = _4371 ^ _448;
  wire _48977 = _48975 ^ _48976;
  wire _48978 = _48974 ^ _48977;
  wire _48979 = _2078 ^ _15355;
  wire _48980 = _48979 ^ _9976;
  wire _48981 = _7680 ^ _12179;
  wire _48982 = _28592 ^ _48981;
  wire _48983 = _48980 ^ _48982;
  wire _48984 = _48978 ^ _48983;
  wire _48985 = _2093 ^ _19268;
  wire _48986 = _48985 ^ _8854;
  wire _48987 = uncoded_block[990] ^ uncoded_block[996];
  wire _48988 = _48987 ^ _5798;
  wire _48989 = _44228 ^ _48988;
  wire _48990 = _48986 ^ _48989;
  wire _48991 = uncoded_block[1007] ^ uncoded_block[1015];
  wire _48992 = _2114 ^ _48991;
  wire _48993 = _48992 ^ _31169;
  wire _48994 = _44635 ^ _3676;
  wire _48995 = _12758 ^ _38937;
  wire _48996 = _48994 ^ _48995;
  wire _48997 = _48993 ^ _48996;
  wire _48998 = _48990 ^ _48997;
  wire _48999 = _48984 ^ _48998;
  wire _49000 = _48973 ^ _48999;
  wire _49001 = _48950 ^ _49000;
  wire _49002 = _48900 ^ _49001;
  wire _49003 = uncoded_block[1050] ^ uncoded_block[1056];
  wire _49004 = _514 ^ _49003;
  wire _49005 = _7117 ^ _6483;
  wire _49006 = _49004 ^ _49005;
  wire _49007 = _23502 ^ _36546;
  wire _49008 = _49006 ^ _49007;
  wire _49009 = _3692 ^ _20251;
  wire _49010 = _10575 ^ _1373;
  wire _49011 = _49009 ^ _49010;
  wire _49012 = _23070 ^ _42057;
  wire _49013 = _49011 ^ _49012;
  wire _49014 = _49008 ^ _49013;
  wire _49015 = _545 ^ _10585;
  wire _49016 = _49015 ^ _15411;
  wire _49017 = _15894 ^ _12795;
  wire _49018 = _17377 ^ _49017;
  wire _49019 = _49016 ^ _49018;
  wire _49020 = _2953 ^ _5184;
  wire _49021 = _49020 ^ _38162;
  wire _49022 = _3733 ^ _32884;
  wire _49023 = _2189 ^ _10602;
  wire _49024 = _49022 ^ _49023;
  wire _49025 = _49021 ^ _49024;
  wire _49026 = _49019 ^ _49025;
  wire _49027 = _49014 ^ _49026;
  wire _49028 = uncoded_block[1186] ^ uncoded_block[1191];
  wire _49029 = _592 ^ _49028;
  wire _49030 = _29034 ^ _49029;
  wire _49031 = _1420 ^ _11719;
  wire _49032 = _17400 ^ _1425;
  wire _49033 = _49031 ^ _49032;
  wire _49034 = _49030 ^ _49033;
  wire _49035 = _11171 ^ _10617;
  wire _49036 = _12813 ^ _23105;
  wire _49037 = _49035 ^ _49036;
  wire _49038 = _6532 ^ _4504;
  wire _49039 = _14919 ^ _43141;
  wire _49040 = _49038 ^ _49039;
  wire _49041 = _49037 ^ _49040;
  wire _49042 = _49034 ^ _49041;
  wire _49043 = uncoded_block[1238] ^ uncoded_block[1245];
  wire _49044 = _49043 ^ _5229;
  wire _49045 = _8385 ^ _32082;
  wire _49046 = _49044 ^ _49045;
  wire _49047 = _1456 ^ _22197;
  wire _49048 = _9533 ^ _23123;
  wire _49049 = _49047 ^ _49048;
  wire _49050 = _49046 ^ _49049;
  wire _49051 = _639 ^ _641;
  wire _49052 = _642 ^ _4532;
  wire _49053 = _49051 ^ _49052;
  wire _49054 = _4536 ^ _8991;
  wire _49055 = _49054 ^ _41329;
  wire _49056 = _49053 ^ _49055;
  wire _49057 = _49050 ^ _49056;
  wire _49058 = _49042 ^ _49057;
  wire _49059 = _49027 ^ _49058;
  wire _49060 = _1486 ^ _19375;
  wire _49061 = _16435 ^ _4551;
  wire _49062 = _49060 ^ _49061;
  wire _49063 = _5259 ^ _7815;
  wire _49064 = _9003 ^ _11771;
  wire _49065 = _49063 ^ _49064;
  wire _49066 = _49062 ^ _49065;
  wire _49067 = uncoded_block[1351] ^ uncoded_block[1359];
  wire _49068 = _49067 ^ _27157;
  wire _49069 = _2283 ^ _5281;
  wire _49070 = _49068 ^ _49069;
  wire _49071 = uncoded_block[1378] ^ uncoded_block[1384];
  wire _49072 = _49071 ^ _11782;
  wire _49073 = _17947 ^ _49072;
  wire _49074 = _49070 ^ _49073;
  wire _49075 = _49066 ^ _49074;
  wire _49076 = _692 ^ _13416;
  wire _49077 = _49076 ^ _46449;
  wire _49078 = _3847 ^ _15492;
  wire _49079 = _5964 ^ _24058;
  wire _49080 = _49078 ^ _49079;
  wire _49081 = _49077 ^ _49080;
  wire _49082 = _2314 ^ _3083;
  wire _49083 = _20352 ^ _49082;
  wire _49084 = _9034 ^ _46458;
  wire _49085 = _49083 ^ _49084;
  wire _49086 = _49081 ^ _49085;
  wire _49087 = _49075 ^ _49086;
  wire _49088 = uncoded_block[1456] ^ uncoded_block[1461];
  wire _49089 = _49088 ^ _2336;
  wire _49090 = _49089 ^ _42519;
  wire _49091 = uncoded_block[1470] ^ uncoded_block[1474];
  wire _49092 = _49091 ^ _2342;
  wire _49093 = _49092 ^ _48354;
  wire _49094 = _49090 ^ _49093;
  wire _49095 = _13967 ^ _2352;
  wire _49096 = _13451 ^ _49095;
  wire _49097 = uncoded_block[1500] ^ uncoded_block[1505];
  wire _49098 = _49097 ^ _3112;
  wire _49099 = _49098 ^ _13456;
  wire _49100 = _49096 ^ _49099;
  wire _49101 = _49094 ^ _49100;
  wire _49102 = _9055 ^ _5341;
  wire _49103 = _49102 ^ _10720;
  wire _49104 = _3906 ^ _1589;
  wire _49105 = _32972 ^ _49104;
  wire _49106 = _49103 ^ _49105;
  wire _49107 = _13472 ^ _767;
  wire _49108 = _31729 ^ _49107;
  wire _49109 = _22731 ^ _11283;
  wire _49110 = _7891 ^ _15026;
  wire _49111 = _49109 ^ _49110;
  wire _49112 = _49108 ^ _49111;
  wire _49113 = _49106 ^ _49112;
  wire _49114 = _49101 ^ _49113;
  wire _49115 = _49087 ^ _49114;
  wire _49116 = _49059 ^ _49115;
  wire _49117 = _13478 ^ _15535;
  wire _49118 = _49117 ^ _16022;
  wire _49119 = _15031 ^ _20401;
  wire _49120 = _49119 ^ _14516;
  wire _49121 = _49118 ^ _49120;
  wire _49122 = uncoded_block[1599] ^ uncoded_block[1604];
  wire _49123 = _49122 ^ _1625;
  wire _49124 = _4662 ^ _17020;
  wire _49125 = _49123 ^ _49124;
  wire _49126 = _29145 ^ _36260;
  wire _49127 = _49125 ^ _49126;
  wire _49128 = _49121 ^ _49127;
  wire _49129 = _48386 ^ _18027;
  wire _49130 = _3172 ^ _9106;
  wire _49131 = _10760 ^ _7927;
  wire _49132 = _49130 ^ _49131;
  wire _49133 = _49129 ^ _49132;
  wire _49134 = _3182 ^ _3186;
  wire _49135 = _9110 ^ _49134;
  wire _49136 = _836 ^ _30900;
  wire _49137 = _49136 ^ _32190;
  wire _49138 = _49135 ^ _49137;
  wire _49139 = _49133 ^ _49138;
  wire _49140 = _49128 ^ _49139;
  wire _49141 = _6068 ^ _3976;
  wire _49142 = _7335 ^ _3988;
  wire _49143 = _49141 ^ _49142;
  wire _49144 = _49143 ^ uncoded_block[1721];
  wire _49145 = _49140 ^ _49144;
  wire _49146 = _49116 ^ _49145;
  wire _49147 = _49002 ^ _49146;
  wire _49148 = _4710 ^ _6080;
  wire _49149 = _2454 ^ _3998;
  wire _49150 = _49148 ^ _49149;
  wire _49151 = _13537 ^ _11343;
  wire _49152 = uncoded_block[28] ^ uncoded_block[34];
  wire _49153 = _7959 ^ _49152;
  wire _49154 = _49151 ^ _49153;
  wire _49155 = _49150 ^ _49154;
  wire _49156 = _879 ^ _10796;
  wire _49157 = _20457 ^ _6099;
  wire _49158 = _49156 ^ _49157;
  wire _49159 = _1700 ^ _12996;
  wire _49160 = _49159 ^ _14581;
  wire _49161 = _49158 ^ _49160;
  wire _49162 = _49155 ^ _49161;
  wire _49163 = uncoded_block[68] ^ uncoded_block[73];
  wire _49164 = _49163 ^ _5443;
  wire _49165 = _49164 ^ _6751;
  wire _49166 = _9713 ^ _46;
  wire _49167 = _42592 ^ _49166;
  wire _49168 = _49165 ^ _49167;
  wire _49169 = uncoded_block[97] ^ uncoded_block[103];
  wire _49170 = _49169 ^ _50;
  wire _49171 = uncoded_block[112] ^ uncoded_block[121];
  wire _49172 = _49171 ^ _20961;
  wire _49173 = _49170 ^ _49172;
  wire _49174 = _13017 ^ _4042;
  wire _49175 = _23720 ^ _11918;
  wire _49176 = _49174 ^ _49175;
  wire _49177 = _49173 ^ _49176;
  wire _49178 = _49168 ^ _49177;
  wire _49179 = _49162 ^ _49178;
  wire _49180 = uncoded_block[143] ^ uncoded_block[150];
  wire _49181 = _49180 ^ _24182;
  wire _49182 = _6785 ^ _8589;
  wire _49183 = _49181 ^ _49182;
  wire _49184 = uncoded_block[172] ^ uncoded_block[177];
  wire _49185 = _8591 ^ _49184;
  wire _49186 = _5477 ^ _4062;
  wire _49187 = _49185 ^ _49186;
  wire _49188 = _49183 ^ _49187;
  wire _49189 = _6156 ^ _32247;
  wire _49190 = _1764 ^ _21459;
  wire _49191 = _46188 ^ _49190;
  wire _49192 = _49189 ^ _49191;
  wire _49193 = _49188 ^ _49192;
  wire _49194 = _3296 ^ _14105;
  wire _49195 = _4076 ^ _20990;
  wire _49196 = _49194 ^ _49195;
  wire _49197 = _3308 ^ _31834;
  wire _49198 = _46196 ^ _49197;
  wire _49199 = _49196 ^ _49198;
  wire _49200 = _1786 ^ _13609;
  wire _49201 = _26000 ^ _985;
  wire _49202 = _49200 ^ _49201;
  wire _49203 = uncoded_block[273] ^ uncoded_block[278];
  wire _49204 = _49203 ^ _12506;
  wire _49205 = _11424 ^ _1804;
  wire _49206 = _49204 ^ _49205;
  wire _49207 = _49202 ^ _49206;
  wire _49208 = _49199 ^ _49207;
  wire _49209 = _49193 ^ _49208;
  wire _49210 = _49179 ^ _49209;
  wire _49211 = _2573 ^ _10312;
  wire _49212 = _49211 ^ _20535;
  wire _49213 = _22866 ^ _9233;
  wire _49214 = _13618 ^ _49213;
  wire _49215 = _49212 ^ _49214;
  wire _49216 = _150 ^ _152;
  wire _49217 = _49216 ^ _16153;
  wire _49218 = _6857 ^ _10323;
  wire _49219 = _49218 ^ _46219;
  wire _49220 = _49217 ^ _49219;
  wire _49221 = _49215 ^ _49220;
  wire _49222 = _30123 ^ _2602;
  wire _49223 = _33119 ^ _5548;
  wire _49224 = _49222 ^ _49223;
  wire _49225 = _1835 ^ _169;
  wire _49226 = _6876 ^ _19599;
  wire _49227 = _49225 ^ _49226;
  wire _49228 = _49224 ^ _49227;
  wire _49229 = uncoded_block[396] ^ uncoded_block[401];
  wire _49230 = _3383 ^ _49229;
  wire _49231 = uncoded_block[404] ^ uncoded_block[409];
  wire _49232 = _2625 ^ _49231;
  wire _49233 = _49230 ^ _49232;
  wire _49234 = uncoded_block[410] ^ uncoded_block[417];
  wire _49235 = _49234 ^ _24707;
  wire _49236 = _49235 ^ _35963;
  wire _49237 = _49233 ^ _49236;
  wire _49238 = _49228 ^ _49237;
  wire _49239 = _49221 ^ _49238;
  wire _49240 = _13117 ^ _5577;
  wire _49241 = _21974 ^ _1069;
  wire _49242 = _49240 ^ _49241;
  wire _49243 = _38796 ^ _9282;
  wire _49244 = _49242 ^ _49243;
  wire _49245 = _9284 ^ _1084;
  wire _49246 = uncoded_block[475] ^ uncoded_block[481];
  wire _49247 = _49246 ^ _8694;
  wire _49248 = _17198 ^ _1093;
  wire _49249 = _49247 ^ _49248;
  wire _49250 = _49245 ^ _49249;
  wire _49251 = _49244 ^ _49250;
  wire _49252 = _13140 ^ _43733;
  wire _49253 = uncoded_block[511] ^ uncoded_block[516];
  wire _49254 = _49253 ^ _19638;
  wire _49255 = _29288 ^ _49254;
  wire _49256 = _49252 ^ _49255;
  wire _49257 = _1899 ^ _30173;
  wire _49258 = _1905 ^ _24279;
  wire _49259 = _14198 ^ _3453;
  wire _49260 = _49258 ^ _49259;
  wire _49261 = _49257 ^ _49260;
  wire _49262 = _49256 ^ _49261;
  wire _49263 = _49251 ^ _49262;
  wire _49264 = _49239 ^ _49263;
  wire _49265 = _49210 ^ _49264;
  wire _49266 = _6300 ^ _1913;
  wire _49267 = _49266 ^ _26086;
  wire _49268 = uncoded_block[564] ^ uncoded_block[569];
  wire _49269 = _4937 ^ _49268;
  wire _49270 = _49269 ^ _48536;
  wire _49271 = _49267 ^ _49270;
  wire _49272 = _270 ^ _18222;
  wire _49273 = _41939 ^ _49272;
  wire _49274 = _25640 ^ _7558;
  wire _49275 = _28516 ^ _49274;
  wire _49276 = _49273 ^ _49275;
  wire _49277 = _49271 ^ _49276;
  wire _49278 = _8738 ^ _1942;
  wire _49279 = _49278 ^ _14222;
  wire _49280 = uncoded_block[615] ^ uncoded_block[623];
  wire _49281 = _49280 ^ _5658;
  wire _49282 = _8161 ^ _12621;
  wire _49283 = _49281 ^ _49282;
  wire _49284 = _49279 ^ _49283;
  wire _49285 = _297 ^ _304;
  wire _49286 = _14749 ^ _49285;
  wire _49287 = _46283 ^ _37271;
  wire _49288 = _49286 ^ _49287;
  wire _49289 = _49284 ^ _49288;
  wire _49290 = _49277 ^ _49289;
  wire _49291 = _6352 ^ _23856;
  wire _49292 = _49291 ^ _15283;
  wire _49293 = _18719 ^ _18721;
  wire _49294 = _49293 ^ _46295;
  wire _49295 = _49292 ^ _49294;
  wire _49296 = _21126 ^ _6999;
  wire _49297 = _7603 ^ _32779;
  wire _49298 = _49296 ^ _49297;
  wire _49299 = _1996 ^ _33213;
  wire _49300 = uncoded_block[749] ^ uncoded_block[754];
  wire _49301 = _5013 ^ _49300;
  wire _49302 = _49299 ^ _49301;
  wire _49303 = _49298 ^ _49302;
  wire _49304 = _49295 ^ _49303;
  wire _49305 = uncoded_block[759] ^ uncoded_block[765];
  wire _49306 = _4298 ^ _49305;
  wire _49307 = _17776 ^ _6382;
  wire _49308 = _49306 ^ _49307;
  wire _49309 = uncoded_block[784] ^ uncoded_block[789];
  wire _49310 = _3568 ^ _49309;
  wire _49311 = _7621 ^ _49310;
  wire _49312 = _49308 ^ _49311;
  wire _49313 = _1232 ^ _3576;
  wire _49314 = _7629 ^ _1238;
  wire _49315 = _49313 ^ _49314;
  wire _49316 = _392 ^ _11030;
  wire _49317 = _1241 ^ _7037;
  wire _49318 = _49316 ^ _49317;
  wire _49319 = _49315 ^ _49318;
  wire _49320 = _49312 ^ _49319;
  wire _49321 = _49304 ^ _49320;
  wire _49322 = _49290 ^ _49321;
  wire _49323 = _1246 ^ _4330;
  wire _49324 = _49323 ^ _46322;
  wire _49325 = _8808 ^ _2820;
  wire _49326 = uncoded_block[850] ^ uncoded_block[855];
  wire _49327 = _49326 ^ _14300;
  wire _49328 = _49325 ^ _49327;
  wire _49329 = _49324 ^ _49328;
  wire _49330 = uncoded_block[864] ^ uncoded_block[867];
  wire _49331 = _2824 ^ _49330;
  wire _49332 = _49331 ^ _38488;
  wire _49333 = _11622 ^ _31572;
  wire _49334 = _49332 ^ _49333;
  wire _49335 = _49329 ^ _49334;
  wire _49336 = _47103 ^ _23913;
  wire _49337 = _3622 ^ _7070;
  wire _49338 = _49337 ^ _40091;
  wire _49339 = _49336 ^ _49338;
  wire _49340 = _17318 ^ _4370;
  wire _49341 = _7670 ^ _4377;
  wire _49342 = _49340 ^ _49341;
  wire _49343 = _19261 ^ _4381;
  wire _49344 = _4382 ^ _5105;
  wire _49345 = _49343 ^ _49344;
  wire _49346 = _49342 ^ _49345;
  wire _49347 = _49339 ^ _49346;
  wire _49348 = _49335 ^ _49347;
  wire _49349 = _10529 ^ _24388;
  wire _49350 = _49349 ^ _13271;
  wire _49351 = _37734 ^ _48243;
  wire _49352 = _49350 ^ _49351;
  wire _49353 = _1318 ^ _8293;
  wire _49354 = _28241 ^ _483;
  wire _49355 = _49353 ^ _49354;
  wire _49356 = _7703 ^ _2894;
  wire _49357 = _6460 ^ _49356;
  wire _49358 = _49355 ^ _49357;
  wire _49359 = _49352 ^ _49358;
  wire _49360 = _9454 ^ _9459;
  wire _49361 = _49360 ^ _7709;
  wire _49362 = _2910 ^ _24417;
  wire _49363 = _49362 ^ _49005;
  wire _49364 = _49361 ^ _49363;
  wire _49365 = uncoded_block[1067] ^ uncoded_block[1071];
  wire _49366 = _20247 ^ _49365;
  wire _49367 = _12770 ^ _5163;
  wire _49368 = _49366 ^ _49367;
  wire _49369 = _11687 ^ _20253;
  wire _49370 = _5840 ^ _1380;
  wire _49371 = _49369 ^ _49370;
  wire _49372 = _49368 ^ _49371;
  wire _49373 = _49364 ^ _49372;
  wire _49374 = _49359 ^ _49373;
  wire _49375 = _49348 ^ _49374;
  wire _49376 = _49322 ^ _49375;
  wire _49377 = _49265 ^ _49376;
  wire _49378 = _545 ^ _2164;
  wire _49379 = _49378 ^ _20764;
  wire _49380 = _8339 ^ _14376;
  wire _49381 = _49380 ^ _30330;
  wire _49382 = _49379 ^ _49381;
  wire _49383 = _38963 ^ _2185;
  wire _49384 = _49383 ^ _46392;
  wire _49385 = uncoded_block[1164] ^ uncoded_block[1170];
  wire _49386 = _49385 ^ _1410;
  wire _49387 = _585 ^ _590;
  wire _49388 = _49386 ^ _49387;
  wire _49389 = _49384 ^ _49388;
  wire _49390 = _49382 ^ _49389;
  wire _49391 = _592 ^ _2196;
  wire _49392 = _13346 ^ _24910;
  wire _49393 = _49391 ^ _49392;
  wire _49394 = _7160 ^ _8370;
  wire _49395 = _49394 ^ _26693;
  wire _49396 = _49393 ^ _49395;
  wire _49397 = uncoded_block[1215] ^ uncoded_block[1220];
  wire _49398 = _1427 ^ _49397;
  wire _49399 = _5891 ^ _13357;
  wire _49400 = _49398 ^ _49399;
  wire _49401 = uncoded_block[1235] ^ uncoded_block[1242];
  wire _49402 = _31228 ^ _49401;
  wire _49403 = _19829 ^ _2997;
  wire _49404 = _49402 ^ _49403;
  wire _49405 = _49400 ^ _49404;
  wire _49406 = _49396 ^ _49405;
  wire _49407 = _49390 ^ _49406;
  wire _49408 = _36165 ^ _37798;
  wire _49409 = _3784 ^ _3786;
  wire _49410 = _3010 ^ _29468;
  wire _49411 = _49409 ^ _49410;
  wire _49412 = _49408 ^ _49411;
  wire _49413 = _16924 ^ _45826;
  wire _49414 = uncoded_block[1301] ^ uncoded_block[1307];
  wire _49415 = _6564 ^ _49414;
  wire _49416 = _49413 ^ _49415;
  wire _49417 = _11759 ^ _3812;
  wire _49418 = _49417 ^ _43163;
  wire _49419 = _49416 ^ _49418;
  wire _49420 = _49412 ^ _49419;
  wire _49421 = _7815 ^ _18436;
  wire _49422 = _5260 ^ _49421;
  wire _49423 = _10097 ^ _7821;
  wire _49424 = _2283 ^ _9572;
  wire _49425 = _49423 ^ _49424;
  wire _49426 = _49422 ^ _49425;
  wire _49427 = _12305 ^ _32935;
  wire _49428 = _18444 ^ _1513;
  wire _49429 = _49427 ^ _49428;
  wire _49430 = _38613 ^ _13938;
  wire _49431 = uncoded_block[1404] ^ uncoded_block[1410];
  wire _49432 = _29090 ^ _49431;
  wire _49433 = _49430 ^ _49432;
  wire _49434 = _49429 ^ _49433;
  wire _49435 = _49426 ^ _49434;
  wire _49436 = _49420 ^ _49435;
  wire _49437 = _49407 ^ _49436;
  wire _49438 = uncoded_block[1411] ^ uncoded_block[1419];
  wire _49439 = _49438 ^ _3853;
  wire _49440 = _3075 ^ _2313;
  wire _49441 = _49439 ^ _49440;
  wire _49442 = _3861 ^ _45085;
  wire _49443 = _31702 ^ _49442;
  wire _49444 = _49441 ^ _49443;
  wire _49445 = _36635 ^ _3088;
  wire _49446 = _40962 ^ _49445;
  wire _49447 = _726 ^ _10136;
  wire _49448 = uncoded_block[1477] ^ uncoded_block[1483];
  wire _49449 = _4603 ^ _49448;
  wire _49450 = _49447 ^ _49449;
  wire _49451 = _49446 ^ _49450;
  wire _49452 = _49444 ^ _49451;
  wire _49453 = _7861 ^ _2349;
  wire _49454 = _49453 ^ _15512;
  wire _49455 = _24539 ^ _19429;
  wire _49456 = _43202 ^ _49455;
  wire _49457 = _49454 ^ _49456;
  wire _49458 = _11267 ^ _12352;
  wire _49459 = _3900 ^ _17499;
  wire _49460 = _49458 ^ _49459;
  wire _49461 = _46474 ^ _6008;
  wire _49462 = _33821 ^ _49461;
  wire _49463 = _49460 ^ _49462;
  wire _49464 = _49457 ^ _49463;
  wire _49465 = _49452 ^ _49464;
  wire _49466 = _17998 ^ _4638;
  wire _49467 = _44372 ^ _24102;
  wire _49468 = _49466 ^ _49467;
  wire _49469 = _14508 ^ _46488;
  wire _49470 = _49468 ^ _49469;
  wire _49471 = uncoded_block[1613] ^ uncoded_block[1617];
  wire _49472 = _49471 ^ _18020;
  wire _49473 = _46494 ^ _49472;
  wire _49474 = _46492 ^ _49473;
  wire _49475 = _49470 ^ _49474;
  wire _49476 = _6046 ^ _808;
  wire _49477 = _49476 ^ _24121;
  wire _49478 = _12949 ^ _1646;
  wire _49479 = _7312 ^ _10757;
  wire _49480 = _49478 ^ _49479;
  wire _49481 = _49477 ^ _49480;
  wire _49482 = _32178 ^ _14011;
  wire _49483 = _49482 ^ _21385;
  wire _49484 = _3182 ^ _11319;
  wire _49485 = _38272 ^ _49484;
  wire _49486 = _49483 ^ _49485;
  wire _49487 = _49481 ^ _49486;
  wire _49488 = _49475 ^ _49487;
  wire _49489 = _49465 ^ _49488;
  wire _49490 = _49437 ^ _49489;
  wire _49491 = _17538 ^ _23671;
  wire _49492 = _24130 ^ _2429;
  wire _49493 = _49491 ^ _49492;
  wire _49494 = _3968 ^ _3973;
  wire _49495 = _49494 ^ _15064;
  wire _49496 = _49493 ^ _49495;
  wire _49497 = _851 ^ _6072;
  wire _49498 = _49497 ^ _21402;
  wire _49499 = _49496 ^ _49498;
  wire _49500 = _49490 ^ _49499;
  wire _49501 = _49377 ^ _49500;
  wire _49502 = uncoded_block[4] ^ uncoded_block[19];
  wire _49503 = uncoded_block[25] ^ uncoded_block[63];
  wire _49504 = _49502 ^ _49503;
  wire _49505 = uncoded_block[86] ^ uncoded_block[107];
  wire _49506 = _14060 ^ _49505;
  wire _49507 = _49504 ^ _49506;
  wire _49508 = uncoded_block[126] ^ uncoded_block[145];
  wire _49509 = _49508 ^ _45938;
  wire _49510 = uncoded_block[164] ^ uncoded_block[187];
  wire _49511 = _49510 ^ _9200;
  wire _49512 = _49509 ^ _49511;
  wire _49513 = _49507 ^ _49512;
  wire _49514 = _32251 ^ _4081;
  wire _49515 = uncoded_block[235] ^ uncoded_block[246];
  wire _49516 = uncoded_block[261] ^ uncoded_block[285];
  wire _49517 = _49515 ^ _49516;
  wire _49518 = _49514 ^ _49517;
  wire _49519 = uncoded_block[290] ^ uncoded_block[302];
  wire _49520 = uncoded_block[311] ^ uncoded_block[331];
  wire _49521 = _49519 ^ _49520;
  wire _49522 = uncoded_block[340] ^ uncoded_block[349];
  wire _49523 = uncoded_block[355] ^ uncoded_block[366];
  wire _49524 = _49522 ^ _49523;
  wire _49525 = _49521 ^ _49524;
  wire _49526 = _49518 ^ _49525;
  wire _49527 = _49513 ^ _49526;
  wire _49528 = uncoded_block[376] ^ uncoded_block[395];
  wire _49529 = _49528 ^ _191;
  wire _49530 = uncoded_block[471] ^ uncoded_block[494];
  wire _49531 = _1874 ^ _49530;
  wire _49532 = _49529 ^ _49531;
  wire _49533 = uncoded_block[495] ^ uncoded_block[507];
  wire _49534 = uncoded_block[510] ^ uncoded_block[540];
  wire _49535 = _49533 ^ _49534;
  wire _49536 = uncoded_block[545] ^ uncoded_block[558];
  wire _49537 = uncoded_block[565] ^ uncoded_block[574];
  wire _49538 = _49536 ^ _49537;
  wire _49539 = _49535 ^ _49538;
  wire _49540 = _49532 ^ _49539;
  wire _49541 = uncoded_block[581] ^ uncoded_block[591];
  wire _49542 = uncoded_block[612] ^ uncoded_block[627];
  wire _49543 = _49541 ^ _49542;
  wire _49544 = _10984 ^ _15766;
  wire _49545 = _49543 ^ _49544;
  wire _49546 = uncoded_block[669] ^ uncoded_block[698];
  wire _49547 = _49546 ^ _4999;
  wire _49548 = uncoded_block[719] ^ uncoded_block[727];
  wire _49549 = _49548 ^ _14266;
  wire _49550 = _49547 ^ _49549;
  wire _49551 = _49545 ^ _49550;
  wire _49552 = _49540 ^ _49551;
  wire _49553 = _49527 ^ _49552;
  wire _49554 = uncoded_block[785] ^ uncoded_block[790];
  wire _49555 = _4301 ^ _49554;
  wire _49556 = uncoded_block[818] ^ uncoded_block[834];
  wire _49557 = _45716 ^ _49556;
  wire _49558 = _49555 ^ _49557;
  wire _49559 = uncoded_block[848] ^ uncoded_block[879];
  wire _49560 = uncoded_block[885] ^ uncoded_block[893];
  wire _49561 = _49559 ^ _49560;
  wire _49562 = uncoded_block[900] ^ uncoded_block[918];
  wire _49563 = uncoded_block[919] ^ uncoded_block[925];
  wire _49564 = _49562 ^ _49563;
  wire _49565 = _49561 ^ _49564;
  wire _49566 = _49558 ^ _49565;
  wire _49567 = uncoded_block[958] ^ uncoded_block[967];
  wire _49568 = uncoded_block[968] ^ uncoded_block[996];
  wire _49569 = _49567 ^ _49568;
  wire _49570 = uncoded_block[1000] ^ uncoded_block[1013];
  wire _49571 = uncoded_block[1016] ^ uncoded_block[1025];
  wire _49572 = _49570 ^ _49571;
  wire _49573 = _49569 ^ _49572;
  wire _49574 = uncoded_block[1026] ^ uncoded_block[1049];
  wire _49575 = uncoded_block[1064] ^ uncoded_block[1082];
  wire _49576 = _49574 ^ _49575;
  wire _49577 = uncoded_block[1102] ^ uncoded_block[1136];
  wire _49578 = _36955 ^ _49577;
  wire _49579 = _49576 ^ _49578;
  wire _49580 = _49573 ^ _49579;
  wire _49581 = _49566 ^ _49580;
  wire _49582 = _4462 ^ _8937;
  wire _49583 = uncoded_block[1188] ^ uncoded_block[1198];
  wire _49584 = uncoded_block[1209] ^ uncoded_block[1219];
  wire _49585 = _49583 ^ _49584;
  wire _49586 = _49582 ^ _49585;
  wire _49587 = uncoded_block[1222] ^ uncoded_block[1238];
  wire _49588 = uncoded_block[1248] ^ uncoded_block[1256];
  wire _49589 = _49587 ^ _49588;
  wire _49590 = uncoded_block[1266] ^ uncoded_block[1290];
  wire _49591 = uncoded_block[1295] ^ uncoded_block[1318];
  wire _49592 = _49590 ^ _49591;
  wire _49593 = _49589 ^ _49592;
  wire _49594 = _49586 ^ _49593;
  wire _49595 = uncoded_block[1327] ^ uncoded_block[1347];
  wire _49596 = uncoded_block[1355] ^ uncoded_block[1375];
  wire _49597 = _49595 ^ _49596;
  wire _49598 = _35016 ^ _3849;
  wire _49599 = _49597 ^ _49598;
  wire _49600 = uncoded_block[1430] ^ uncoded_block[1456];
  wire _49601 = uncoded_block[1470] ^ uncoded_block[1478];
  wire _49602 = _49600 ^ _49601;
  wire _49603 = uncoded_block[1488] ^ uncoded_block[1501];
  wire _49604 = uncoded_block[1521] ^ uncoded_block[1527];
  wire _49605 = _49603 ^ _49604;
  wire _49606 = _49602 ^ _49605;
  wire _49607 = _49599 ^ _49606;
  wire _49608 = _49594 ^ _49607;
  wire _49609 = _49581 ^ _49608;
  wire _49610 = _49553 ^ _49609;
  wire _49611 = uncoded_block[1537] ^ uncoded_block[1553];
  wire _49612 = _49611 ^ _38247;
  wire _49613 = uncoded_block[1592] ^ uncoded_block[1622];
  wire _49614 = _39838 ^ _49613;
  wire _49615 = _49612 ^ _49614;
  wire _49616 = uncoded_block[1626] ^ uncoded_block[1637];
  wire _49617 = _49616 ^ _20905;
  wire _49618 = _36687 ^ _7319;
  wire _49619 = _49617 ^ _49618;
  wire _49620 = _49615 ^ _49619;
  wire _49621 = uncoded_block[1691] ^ uncoded_block[1709];
  wire _49622 = _49621 ^ uncoded_block[1715];
  wire _49623 = _49620 ^ _49622;
  wire _49624 = _49610 ^ _49623;
  wire _49625 = uncoded_block[5] ^ uncoded_block[12];
  wire _49626 = _16560 ^ _49625;
  wire _49627 = uncoded_block[13] ^ uncoded_block[18];
  wire _49628 = _49627 ^ _3217;
  wire _49629 = _49626 ^ _49628;
  wire _49630 = _3220 ^ _11344;
  wire _49631 = _49630 ^ _46155;
  wire _49632 = _49629 ^ _49631;
  wire _49633 = _4008 ^ _8556;
  wire _49634 = _23697 ^ _2474;
  wire _49635 = _49633 ^ _49634;
  wire _49636 = _12435 ^ _34;
  wire _49637 = _35 ^ _34689;
  wire _49638 = _49636 ^ _49637;
  wire _49639 = _49635 ^ _49638;
  wire _49640 = _49632 ^ _49639;
  wire _49641 = _11363 ^ _14586;
  wire _49642 = _18077 ^ _6115;
  wire _49643 = _49641 ^ _49642;
  wire _49644 = _19025 ^ _50;
  wire _49645 = _45166 ^ _49644;
  wire _49646 = _49643 ^ _49645;
  wire _49647 = _5453 ^ _6769;
  wire _49648 = _2497 ^ _13016;
  wire _49649 = _49647 ^ _49648;
  wire _49650 = _3263 ^ _4760;
  wire _49651 = _49174 ^ _49650;
  wire _49652 = _49649 ^ _49651;
  wire _49653 = _49646 ^ _49652;
  wire _49654 = _49640 ^ _49653;
  wire _49655 = _6776 ^ _33909;
  wire _49656 = uncoded_block[151] ^ uncoded_block[157];
  wire _49657 = _1744 ^ _49656;
  wire _49658 = _49655 ^ _49657;
  wire _49659 = _15118 ^ _6785;
  wire _49660 = _4054 ^ _1752;
  wire _49661 = _49659 ^ _49660;
  wire _49662 = _49658 ^ _49661;
  wire _49663 = uncoded_block[172] ^ uncoded_block[179];
  wire _49664 = uncoded_block[182] ^ uncoded_block[185];
  wire _49665 = _49663 ^ _49664;
  wire _49666 = uncoded_block[186] ^ uncoded_block[191];
  wire _49667 = _49666 ^ _20500;
  wire _49668 = _49665 ^ _49667;
  wire _49669 = _32247 ^ _46188;
  wire _49670 = _49668 ^ _49669;
  wire _49671 = _49662 ^ _49670;
  wire _49672 = uncoded_block[205] ^ uncoded_block[212];
  wire _49673 = _49672 ^ _3296;
  wire _49674 = _20013 ^ _23739;
  wire _49675 = _49673 ^ _49674;
  wire _49676 = _6169 ^ _22380;
  wire _49677 = _49676 ^ _20510;
  wire _49678 = _49675 ^ _49677;
  wire _49679 = _2556 ^ _3309;
  wire _49680 = _37956 ^ _49679;
  wire _49681 = _120 ^ _21472;
  wire _49682 = _17132 ^ _49681;
  wire _49683 = _49680 ^ _49682;
  wire _49684 = _49678 ^ _49683;
  wire _49685 = _49671 ^ _49684;
  wire _49686 = _49654 ^ _49685;
  wire _49687 = uncoded_block[284] ^ uncoded_block[288];
  wire _49688 = _6834 ^ _49687;
  wire _49689 = _17635 ^ _1807;
  wire _49690 = _49688 ^ _49689;
  wire _49691 = _4824 ^ _4826;
  wire _49692 = _6845 ^ _3334;
  wire _49693 = _49691 ^ _49692;
  wire _49694 = _49690 ^ _49693;
  wire _49695 = _6846 ^ _1006;
  wire _49696 = _3347 ^ _11444;
  wire _49697 = _49695 ^ _49696;
  wire _49698 = _9235 ^ _4838;
  wire _49699 = _11984 ^ _4129;
  wire _49700 = _49698 ^ _49699;
  wire _49701 = _49697 ^ _49700;
  wire _49702 = _49694 ^ _49701;
  wire _49703 = _6218 ^ _8652;
  wire _49704 = _2599 ^ _9249;
  wire _49705 = _49703 ^ _49704;
  wire _49706 = _1838 ^ _13094;
  wire _49707 = _22413 ^ _49706;
  wire _49708 = _49705 ^ _49707;
  wire _49709 = _13101 ^ _31005;
  wire _49710 = _4151 ^ _8661;
  wire _49711 = _49709 ^ _49710;
  wire _49712 = _13646 ^ _3391;
  wire _49713 = _1054 ^ _12548;
  wire _49714 = _49712 ^ _49713;
  wire _49715 = _49711 ^ _49714;
  wire _49716 = _49708 ^ _49715;
  wire _49717 = _49702 ^ _49716;
  wire _49718 = _2638 ^ _8098;
  wire _49719 = _29270 ^ _49718;
  wire _49720 = _12559 ^ _6259;
  wire _49721 = _49720 ^ _2652;
  wire _49722 = _49719 ^ _49721;
  wire _49723 = _22907 ^ _23800;
  wire _49724 = uncoded_block[475] ^ uncoded_block[482];
  wire _49725 = _1082 ^ _49724;
  wire _49726 = _49723 ^ _49725;
  wire _49727 = _9832 ^ _27769;
  wire _49728 = _17197 ^ _49727;
  wire _49729 = _49726 ^ _49728;
  wire _49730 = _49722 ^ _49729;
  wire _49731 = _5604 ^ _21536;
  wire _49732 = _5607 ^ _5611;
  wire _49733 = _49731 ^ _49732;
  wire _49734 = _10943 ^ _4209;
  wire _49735 = _49733 ^ _49734;
  wire _49736 = _1108 ^ _1900;
  wire _49737 = _15230 ^ _3451;
  wire _49738 = _49736 ^ _49737;
  wire _49739 = _4217 ^ _25173;
  wire _49740 = _13689 ^ _4933;
  wire _49741 = _49739 ^ _49740;
  wire _49742 = _49738 ^ _49741;
  wire _49743 = _49735 ^ _49742;
  wire _49744 = _49730 ^ _49743;
  wire _49745 = _49717 ^ _49744;
  wire _49746 = _49686 ^ _49745;
  wire _49747 = _15236 ^ _8724;
  wire _49748 = uncoded_block[557] ^ uncoded_block[562];
  wire _49749 = _49748 ^ _24745;
  wire _49750 = _49747 ^ _49749;
  wire _49751 = _3472 ^ _28136;
  wire _49752 = _49751 ^ _28513;
  wire _49753 = _49750 ^ _49752;
  wire _49754 = uncoded_block[588] ^ uncoded_block[594];
  wire _49755 = _8143 ^ _49754;
  wire _49756 = _49755 ^ _24293;
  wire _49757 = _14219 ^ _13712;
  wire _49758 = _49756 ^ _49757;
  wire _49759 = _49753 ^ _49758;
  wire _49760 = _7567 ^ _1946;
  wire _49761 = _4963 ^ _287;
  wire _49762 = _49760 ^ _49761;
  wire _49763 = _293 ^ _9343;
  wire _49764 = _25652 ^ _49763;
  wire _49765 = _49762 ^ _49764;
  wire _49766 = _298 ^ _40796;
  wire _49767 = _7582 ^ _31072;
  wire _49768 = _3515 ^ _49767;
  wire _49769 = _49766 ^ _49768;
  wire _49770 = _49765 ^ _49769;
  wire _49771 = _49759 ^ _49770;
  wire _49772 = _3519 ^ _1971;
  wire _49773 = _49772 ^ _22491;
  wire _49774 = _4272 ^ _30641;
  wire _49775 = _49774 ^ _33200;
  wire _49776 = _49773 ^ _49775;
  wire _49777 = _6364 ^ _4996;
  wire _49778 = _33205 ^ _1194;
  wire _49779 = _49777 ^ _49778;
  wire _49780 = uncoded_block[719] ^ uncoded_block[724];
  wire _49781 = _49780 ^ _6999;
  wire _49782 = _1202 ^ _7005;
  wire _49783 = _49781 ^ _49782;
  wire _49784 = _49779 ^ _49783;
  wire _49785 = _49776 ^ _49784;
  wire _49786 = uncoded_block[739] ^ uncoded_block[747];
  wire _49787 = _49786 ^ _5704;
  wire _49788 = _5017 ^ _359;
  wire _49789 = _49787 ^ _49788;
  wire _49790 = uncoded_block[769] ^ uncoded_block[773];
  wire _49791 = _27427 ^ _49790;
  wire _49792 = _36469 ^ _5029;
  wire _49793 = _49791 ^ _49792;
  wire _49794 = _49789 ^ _49793;
  wire _49795 = _375 ^ _2022;
  wire _49796 = _38079 ^ _49795;
  wire _49797 = _11029 ^ _9397;
  wire _49798 = _46315 ^ _49797;
  wire _49799 = _49796 ^ _49798;
  wire _49800 = _49794 ^ _49799;
  wire _49801 = _49785 ^ _49800;
  wire _49802 = _49771 ^ _49801;
  wire _49803 = uncoded_block[823] ^ uncoded_block[831];
  wire _49804 = _12131 ^ _49803;
  wire _49805 = _49804 ^ _2816;
  wire _49806 = _11610 ^ _21165;
  wire _49807 = _49806 ^ _5067;
  wire _49808 = _49805 ^ _49807;
  wire _49809 = _17804 ^ _1266;
  wire _49810 = _12150 ^ _25719;
  wire _49811 = _49809 ^ _49810;
  wire _49812 = _11059 ^ _2061;
  wire _49813 = _22090 ^ _49812;
  wire _49814 = _49811 ^ _49813;
  wire _49815 = _49808 ^ _49814;
  wire _49816 = _3614 ^ _5085;
  wire _49817 = _2843 ^ _9960;
  wire _49818 = _49816 ^ _49817;
  wire _49819 = uncoded_block[906] ^ uncoded_block[910];
  wire _49820 = _8254 ^ _49819;
  wire _49821 = _49820 ^ _2853;
  wire _49822 = _49818 ^ _49821;
  wire _49823 = _15350 ^ _8835;
  wire _49824 = _12717 ^ _11076;
  wire _49825 = _49823 ^ _49824;
  wire _49826 = _13266 ^ _1303;
  wire _49827 = _11078 ^ _49826;
  wire _49828 = _49825 ^ _49827;
  wire _49829 = _49822 ^ _49828;
  wire _49830 = _49815 ^ _49829;
  wire _49831 = _14844 ^ _15363;
  wire _49832 = _25280 ^ _49831;
  wire _49833 = uncoded_block[975] ^ uncoded_block[981];
  wire _49834 = _19268 ^ _49833;
  wire _49835 = _49834 ^ _44228;
  wire _49836 = _49832 ^ _49835;
  wire _49837 = uncoded_block[992] ^ uncoded_block[998];
  wire _49838 = _15369 ^ _49837;
  wire _49839 = _49838 ^ _1328;
  wire _49840 = _14343 ^ _38127;
  wire _49841 = _49839 ^ _49840;
  wire _49842 = _49836 ^ _49841;
  wire _49843 = _495 ^ _36938;
  wire _49844 = _49843 ^ _44246;
  wire _49845 = _8309 ^ _519;
  wire _49846 = _47143 ^ _49845;
  wire _49847 = _49844 ^ _49846;
  wire _49848 = _10569 ^ _13851;
  wire _49849 = _3686 ^ _49848;
  wire _49850 = _13307 ^ _20251;
  wire _49851 = uncoded_block[1085] ^ uncoded_block[1090];
  wire _49852 = _10575 ^ _49851;
  wire _49853 = _49850 ^ _49852;
  wire _49854 = _49849 ^ _49853;
  wire _49855 = _49847 ^ _49854;
  wire _49856 = _49842 ^ _49855;
  wire _49857 = _49830 ^ _49856;
  wire _49858 = _49802 ^ _49857;
  wire _49859 = _49746 ^ _49858;
  wire _49860 = _1380 ^ _8336;
  wire _49861 = _37374 ^ _49860;
  wire _49862 = uncoded_block[1110] ^ uncoded_block[1118];
  wire _49863 = _49862 ^ _10587;
  wire _49864 = _2172 ^ _2945;
  wire _49865 = _49863 ^ _49864;
  wire _49866 = _49861 ^ _49865;
  wire _49867 = _4462 ^ _2953;
  wire _49868 = _22621 ^ _49867;
  wire _49869 = uncoded_block[1152] ^ uncoded_block[1157];
  wire _49870 = _49869 ^ _3733;
  wire _49871 = _24900 ^ _49870;
  wire _49872 = _49868 ^ _49871;
  wire _49873 = _49866 ^ _49872;
  wire _49874 = _15907 ^ _584;
  wire _49875 = _585 ^ _4482;
  wire _49876 = _49874 ^ _49875;
  wire _49877 = _35354 ^ _13346;
  wire _49878 = uncoded_block[1196] ^ uncoded_block[1202];
  wire _49879 = _1420 ^ _49878;
  wire _49880 = _49877 ^ _49879;
  wire _49881 = _49876 ^ _49880;
  wire _49882 = uncoded_block[1207] ^ uncoded_block[1210];
  wire _49883 = _2978 ^ _49882;
  wire _49884 = _27911 ^ _3763;
  wire _49885 = _49883 ^ _49884;
  wire _49886 = _3765 ^ _5891;
  wire _49887 = _13357 ^ _40166;
  wire _49888 = _49886 ^ _49887;
  wire _49889 = _49885 ^ _49888;
  wire _49890 = _49881 ^ _49889;
  wire _49891 = _49873 ^ _49890;
  wire _49892 = _31229 ^ _19829;
  wire _49893 = _49892 ^ _9528;
  wire _49894 = _26712 ^ _627;
  wire _49895 = _31657 ^ _49894;
  wire _49896 = _49893 ^ _49895;
  wire _49897 = uncoded_block[1272] ^ uncoded_block[1275];
  wire _49898 = _46419 ^ _49897;
  wire _49899 = _7792 ^ _631;
  wire _49900 = _49898 ^ _49899;
  wire _49901 = _6557 ^ _28317;
  wire _49902 = _18866 ^ _10646;
  wire _49903 = _49901 ^ _49902;
  wire _49904 = _49900 ^ _49903;
  wire _49905 = _49896 ^ _49904;
  wire _49906 = _4532 ^ _5917;
  wire _49907 = _32506 ^ _20816;
  wire _49908 = _49906 ^ _49907;
  wire _49909 = _21293 ^ _9555;
  wire _49910 = _47945 ^ _16435;
  wire _49911 = _49909 ^ _49910;
  wire _49912 = _49908 ^ _49911;
  wire _49913 = _5259 ^ _4553;
  wire _49914 = _4552 ^ _49913;
  wire _49915 = _13927 ^ _4556;
  wire _49916 = _15473 ^ _10097;
  wire _49917 = _49915 ^ _49916;
  wire _49918 = _49914 ^ _49917;
  wire _49919 = _49912 ^ _49918;
  wire _49920 = _49905 ^ _49919;
  wire _49921 = _49891 ^ _49920;
  wire _49922 = _15962 ^ _5281;
  wire _49923 = _35396 ^ _49922;
  wire _49924 = _3055 ^ _11781;
  wire _49925 = _17450 ^ _49924;
  wire _49926 = _49923 ^ _49925;
  wire _49927 = _11782 ^ _5952;
  wire _49928 = _3840 ^ _2296;
  wire _49929 = _49927 ^ _49928;
  wire _49930 = _701 ^ _3069;
  wire _49931 = _30395 ^ _49930;
  wire _49932 = _49929 ^ _49931;
  wire _49933 = _49926 ^ _49932;
  wire _49934 = _3850 ^ _24058;
  wire _49935 = _5968 ^ _2314;
  wire _49936 = _49934 ^ _49935;
  wire _49937 = _712 ^ _1541;
  wire _49938 = _49937 ^ _5977;
  wire _49939 = _49936 ^ _49938;
  wire _49940 = _3088 ^ _2336;
  wire _49941 = _10136 ^ _7247;
  wire _49942 = _49940 ^ _49941;
  wire _49943 = _13447 ^ _41366;
  wire _49944 = _49942 ^ _49943;
  wire _49945 = _49939 ^ _49944;
  wire _49946 = _49933 ^ _49945;
  wire _49947 = uncoded_block[1490] ^ uncoded_block[1494];
  wire _49948 = _740 ^ _49947;
  wire _49949 = _24084 ^ _6637;
  wire _49950 = _49948 ^ _49949;
  wire _49951 = _3898 ^ _15007;
  wire _49952 = _37856 ^ _49951;
  wire _49953 = _49950 ^ _49952;
  wire _49954 = uncoded_block[1535] ^ uncoded_block[1540];
  wire _49955 = _12914 ^ _49954;
  wire _49956 = _49955 ^ _1591;
  wire _49957 = _18492 ^ _5358;
  wire _49958 = _3914 ^ _15022;
  wire _49959 = _49957 ^ _49958;
  wire _49960 = _49956 ^ _49959;
  wire _49961 = _49953 ^ _49960;
  wire _49962 = _6019 ^ _16020;
  wire _49963 = _1608 ^ _3921;
  wire _49964 = _49962 ^ _49963;
  wire _49965 = _6031 ^ _15537;
  wire _49966 = _49965 ^ _15032;
  wire _49967 = _49964 ^ _49966;
  wire _49968 = _791 ^ _6674;
  wire _49969 = _8502 ^ _2396;
  wire _49970 = _49968 ^ _49969;
  wire _49971 = uncoded_block[1611] ^ uncoded_block[1617];
  wire _49972 = _5380 ^ _49971;
  wire _49973 = _40998 ^ _15551;
  wire _49974 = _49972 ^ _49973;
  wire _49975 = _49970 ^ _49974;
  wire _49976 = _49967 ^ _49975;
  wire _49977 = _49961 ^ _49976;
  wire _49978 = _49946 ^ _49977;
  wire _49979 = _49921 ^ _49978;
  wire _49980 = _18965 ^ _6689;
  wire _49981 = _49980 ^ _13501;
  wire _49982 = _9661 ^ _32178;
  wire _49983 = _49982 ^ _39076;
  wire _49984 = _49981 ^ _49983;
  wire _49985 = _2422 ^ _6059;
  wire _49986 = _37891 ^ _49985;
  wire _49987 = _2426 ^ _4693;
  wire _49988 = _837 ^ _6066;
  wire _49989 = _49987 ^ _49988;
  wire _49990 = _49986 ^ _49989;
  wire _49991 = _49984 ^ _49990;
  wire _49992 = _3973 ^ _26832;
  wire _49993 = _49992 ^ _40272;
  wire _49994 = _10780 ^ _861;
  wire _49995 = _49993 ^ _49994;
  wire _49996 = _49991 ^ _49995;
  wire _49997 = _49979 ^ _49996;
  wire _49998 = _49859 ^ _49997;
  wire _49999 = uncoded_block[9] ^ uncoded_block[14];
  wire _50000 = _49999 ^ _5423;
  wire _50001 = _45540 ^ _50000;
  wire _50002 = _12985 ^ _9694;
  wire _50003 = _50002 ^ _42209;
  wire _50004 = _50001 ^ _50003;
  wire _50005 = _15591 ^ _10234;
  wire _50006 = _12991 ^ _50005;
  wire _50007 = _12435 ^ _3241;
  wire _50008 = _43637 ^ _50007;
  wire _50009 = _50006 ^ _50008;
  wire _50010 = _50004 ^ _50009;
  wire _50011 = _11904 ^ _901;
  wire _50012 = _4735 ^ _11364;
  wire _50013 = _50011 ^ _50012;
  wire _50014 = uncoded_block[85] ^ uncoded_block[91];
  wire _50015 = _50014 ^ _6115;
  wire _50016 = _1719 ^ _6120;
  wire _50017 = _50015 ^ _50016;
  wire _50018 = _50013 ^ _50017;
  wire _50019 = _41454 ^ _914;
  wire _50020 = _48432 ^ _4754;
  wire _50021 = _50019 ^ _50020;
  wire _50022 = _3265 ^ _66;
  wire _50023 = _25076 ^ _50022;
  wire _50024 = _50021 ^ _50023;
  wire _50025 = _50018 ^ _50024;
  wire _50026 = _50010 ^ _50025;
  wire _50027 = _67 ^ _15623;
  wire _50028 = _4048 ^ _21905;
  wire _50029 = _50027 ^ _50028;
  wire _50030 = _29624 ^ _42888;
  wire _50031 = _16108 ^ _50030;
  wire _50032 = _50029 ^ _50031;
  wire _50033 = _85 ^ _5479;
  wire _50034 = _3279 ^ _50033;
  wire _50035 = _13588 ^ _6155;
  wire _50036 = _36332 ^ _50035;
  wire _50037 = _50034 ^ _50036;
  wire _50038 = _50032 ^ _50037;
  wire _50039 = _3291 ^ _8600;
  wire _50040 = _33500 ^ _50039;
  wire _50041 = _7415 ^ _102;
  wire _50042 = uncoded_block[221] ^ uncoded_block[226];
  wire _50043 = _50042 ^ _7422;
  wire _50044 = _50041 ^ _50043;
  wire _50045 = _50040 ^ _50044;
  wire _50046 = _10289 ^ _5503;
  wire _50047 = _4085 ^ _6180;
  wire _50048 = _50046 ^ _50047;
  wire _50049 = uncoded_block[248] ^ uncoded_block[253];
  wire _50050 = _50049 ^ _9761;
  wire _50051 = _50050 ^ _16630;
  wire _50052 = _50048 ^ _50051;
  wire _50053 = _50045 ^ _50052;
  wire _50054 = _50038 ^ _50053;
  wire _50055 = _50026 ^ _50054;
  wire _50056 = uncoded_block[267] ^ uncoded_block[275];
  wire _50057 = _12501 ^ _50056;
  wire _50058 = _5513 ^ _1796;
  wire _50059 = _50057 ^ _50058;
  wire _50060 = _1803 ^ _134;
  wire _50061 = _50060 ^ _31844;
  wire _50062 = _50059 ^ _50061;
  wire _50063 = _14133 ^ _41091;
  wire _50064 = _50063 ^ _28070;
  wire _50065 = _23764 ^ _4830;
  wire _50066 = _50065 ^ _3348;
  wire _50067 = _50064 ^ _50066;
  wire _50068 = _50062 ^ _50067;
  wire _50069 = _10887 ^ _1821;
  wire _50070 = _2592 ^ _9242;
  wire _50071 = _50069 ^ _50070;
  wire _50072 = _11450 ^ _5539;
  wire _50073 = _1024 ^ _11455;
  wire _50074 = _50072 ^ _50073;
  wire _50075 = _50071 ^ _50074;
  wire _50076 = uncoded_block[357] ^ uncoded_block[363];
  wire _50077 = _50076 ^ _168;
  wire _50078 = _17165 ^ _1036;
  wire _50079 = _50077 ^ _50078;
  wire _50080 = _7474 ^ _12538;
  wire _50081 = _10901 ^ _2613;
  wire _50082 = _50080 ^ _50081;
  wire _50083 = _50079 ^ _50082;
  wire _50084 = _50075 ^ _50083;
  wire _50085 = _50068 ^ _50084;
  wire _50086 = _3384 ^ _1849;
  wire _50087 = _37603 ^ _50086;
  wire _50088 = _4865 ^ _9810;
  wire _50089 = _50088 ^ _47372;
  wire _50090 = _50087 ^ _50089;
  wire _50091 = _8672 ^ _13115;
  wire _50092 = _14684 ^ _50091;
  wire _50093 = _1066 ^ _5574;
  wire _50094 = _205 ^ _1864;
  wire _50095 = _50093 ^ _50094;
  wire _50096 = _50092 ^ _50095;
  wire _50097 = _50090 ^ _50096;
  wire _50098 = _4176 ^ _12562;
  wire _50099 = _26495 ^ _1874;
  wire _50100 = _50098 ^ _50099;
  wire _50101 = _1083 ^ _5593;
  wire _50102 = _8687 ^ _50101;
  wire _50103 = _50100 ^ _50102;
  wire _50104 = _19627 ^ _9833;
  wire _50105 = _14183 ^ _4905;
  wire _50106 = _229 ^ _6283;
  wire _50107 = _50105 ^ _50106;
  wire _50108 = _50104 ^ _50107;
  wire _50109 = _50103 ^ _50108;
  wire _50110 = _50097 ^ _50109;
  wire _50111 = _50085 ^ _50110;
  wire _50112 = _50055 ^ _50111;
  wire _50113 = _3439 ^ _32722;
  wire _50114 = _37230 ^ _9301;
  wire _50115 = _50113 ^ _50114;
  wire _50116 = _34401 ^ _4928;
  wire _50117 = _50115 ^ _50116;
  wire _50118 = _1910 ^ _34404;
  wire _50119 = _1122 ^ _1916;
  wire _50120 = _5633 ^ _32327;
  wire _50121 = _50119 ^ _50120;
  wire _50122 = _50118 ^ _50121;
  wire _50123 = _50117 ^ _50122;
  wire _50124 = _13165 ^ _13698;
  wire _50125 = _50124 ^ _16723;
  wire _50126 = _10400 ^ _6948;
  wire _50127 = _9330 ^ _4236;
  wire _50128 = _50126 ^ _50127;
  wire _50129 = _50125 ^ _50128;
  wire _50130 = _2710 ^ _14739;
  wire _50131 = _38038 ^ _50130;
  wire _50132 = _17232 ^ _8744;
  wire _50133 = _50132 ^ _32339;
  wire _50134 = _50131 ^ _50133;
  wire _50135 = _50129 ^ _50134;
  wire _50136 = _50123 ^ _50135;
  wire _50137 = _5658 ^ _30199;
  wire _50138 = _21102 ^ _50137;
  wire _50139 = _17241 ^ _26990;
  wire _50140 = _50138 ^ _50139;
  wire _50141 = _8166 ^ _8755;
  wire _50142 = _5667 ^ _50141;
  wire _50143 = _2739 ^ _4262;
  wire _50144 = _50143 ^ _9888;
  wire _50145 = _50142 ^ _50144;
  wire _50146 = _50140 ^ _50145;
  wire _50147 = _6349 ^ _18247;
  wire _50148 = _31076 ^ _17754;
  wire _50149 = _50147 ^ _50148;
  wire _50150 = _45691 ^ _10447;
  wire _50151 = _4995 ^ _3535;
  wire _50152 = _50150 ^ _50151;
  wire _50153 = _50149 ^ _50152;
  wire _50154 = _24781 ^ _28925;
  wire _50155 = _7001 ^ _8201;
  wire _50156 = _50155 ^ _45313;
  wire _50157 = _50154 ^ _50156;
  wire _50158 = _50153 ^ _50157;
  wire _50159 = _50146 ^ _50158;
  wire _50160 = _50136 ^ _50159;
  wire _50161 = uncoded_block[750] ^ uncoded_block[758];
  wire _50162 = _50161 ^ _5019;
  wire _50163 = _32368 ^ _50162;
  wire _50164 = _1217 ^ _365;
  wire _50165 = _12113 ^ _15310;
  wire _50166 = _50164 ^ _50165;
  wire _50167 = _50163 ^ _50166;
  wire _50168 = _19217 ^ _5715;
  wire _50169 = _50168 ^ _27021;
  wire _50170 = _5033 ^ _3574;
  wire _50171 = _50170 ^ _48589;
  wire _50172 = _50169 ^ _50171;
  wire _50173 = _50167 ^ _50172;
  wire _50174 = uncoded_block[803] ^ uncoded_block[808];
  wire _50175 = _7029 ^ _50174;
  wire _50176 = _4324 ^ _22525;
  wire _50177 = _50175 ^ _50176;
  wire _50178 = _15320 ^ _33656;
  wire _50179 = _50178 ^ _18293;
  wire _50180 = _50177 ^ _50179;
  wire _50181 = _38481 ^ _3599;
  wire _50182 = _50181 ^ _36489;
  wire _50183 = _2046 ^ _5742;
  wire _50184 = _13244 ^ _2827;
  wire _50185 = _50183 ^ _50184;
  wire _50186 = _50182 ^ _50185;
  wire _50187 = _50180 ^ _50186;
  wire _50188 = _50173 ^ _50187;
  wire _50189 = _2831 ^ _5753;
  wire _50190 = _38488 ^ _50189;
  wire _50191 = _14821 ^ _1273;
  wire _50192 = _18307 ^ _5758;
  wire _50193 = _50191 ^ _50192;
  wire _50194 = _50190 ^ _50193;
  wire _50195 = _1278 ^ _2844;
  wire _50196 = _50195 ^ _34084;
  wire _50197 = _445 ^ _5772;
  wire _50198 = _29818 ^ _50197;
  wire _50199 = _50196 ^ _50198;
  wire _50200 = _50194 ^ _50199;
  wire _50201 = _6440 ^ _11078;
  wire _50202 = _4381 ^ _5105;
  wire _50203 = _464 ^ _11646;
  wire _50204 = _50202 ^ _50203;
  wire _50205 = _50201 ^ _50204;
  wire _50206 = _9981 ^ _11648;
  wire _50207 = _4390 ^ _8286;
  wire _50208 = _50206 ^ _50207;
  wire _50209 = _5790 ^ _7689;
  wire _50210 = _1317 ^ _24855;
  wire _50211 = _50209 ^ _50210;
  wire _50212 = _50208 ^ _50211;
  wire _50213 = _50205 ^ _50212;
  wire _50214 = _50200 ^ _50213;
  wire _50215 = _50188 ^ _50214;
  wire _50216 = _50160 ^ _50215;
  wire _50217 = _50112 ^ _50216;
  wire _50218 = _13277 ^ _28241;
  wire _50219 = _50218 ^ _2113;
  wire _50220 = _43469 ^ _9996;
  wire _50221 = _8871 ^ _1334;
  wire _50222 = _50220 ^ _50221;
  wire _50223 = _50219 ^ _50222;
  wire _50224 = _8301 ^ _2126;
  wire _50225 = _2127 ^ _2908;
  wire _50226 = _50224 ^ _50225;
  wire _50227 = _12199 ^ _22597;
  wire _50228 = _14867 ^ _1364;
  wire _50229 = _50227 ^ _50228;
  wire _50230 = _50226 ^ _50229;
  wire _50231 = _50223 ^ _50230;
  wire _50232 = _25773 ^ _8893;
  wire _50233 = _2147 ^ _12219;
  wire _50234 = _50232 ^ _50233;
  wire _50235 = _32865 ^ _542;
  wire _50236 = uncoded_block[1098] ^ uncoded_block[1106];
  wire _50237 = uncoded_block[1107] ^ uncoded_block[1111];
  wire _50238 = _50236 ^ _50237;
  wire _50239 = _50235 ^ _50238;
  wire _50240 = _50234 ^ _50239;
  wire _50241 = _552 ^ _13322;
  wire _50242 = uncoded_block[1122] ^ uncoded_block[1128];
  wire _50243 = _7736 ^ _50242;
  wire _50244 = _50241 ^ _50243;
  wire _50245 = _8343 ^ _565;
  wire _50246 = _50245 ^ _19326;
  wire _50247 = _50244 ^ _50246;
  wire _50248 = _50240 ^ _50247;
  wire _50249 = _50231 ^ _50248;
  wire _50250 = _17882 ^ _8354;
  wire _50251 = _24442 ^ _26244;
  wire _50252 = _50250 ^ _50251;
  wire _50253 = uncoded_block[1174] ^ uncoded_block[1178];
  wire _50254 = _18382 ^ _50253;
  wire _50255 = _50254 ^ _11716;
  wire _50256 = _50252 ^ _50255;
  wire _50257 = uncoded_block[1189] ^ uncoded_block[1194];
  wire _50258 = _50257 ^ _1421;
  wire _50259 = _11721 ^ _7162;
  wire _50260 = _50258 ^ _50259;
  wire _50261 = _6530 ^ _30351;
  wire _50262 = uncoded_block[1219] ^ uncoded_block[1225];
  wire _50263 = _50262 ^ _17411;
  wire _50264 = _50261 ^ _50263;
  wire _50265 = _50260 ^ _50264;
  wire _50266 = _50256 ^ _50265;
  wire _50267 = _8962 ^ _2995;
  wire _50268 = _50267 ^ _48303;
  wire _50269 = _20801 ^ _26712;
  wire _50270 = _11186 ^ _50269;
  wire _50271 = _50268 ^ _50270;
  wire _50272 = _6550 ^ _7179;
  wire _50273 = _628 ^ _5908;
  wire _50274 = _50272 ^ _50273;
  wire _50275 = _12837 ^ _8980;
  wire _50276 = _30797 ^ _3015;
  wire _50277 = _50275 ^ _50276;
  wire _50278 = _50274 ^ _50277;
  wire _50279 = _50271 ^ _50278;
  wire _50280 = _50266 ^ _50279;
  wire _50281 = _50249 ^ _50280;
  wire _50282 = uncoded_block[1306] ^ uncoded_block[1309];
  wire _50283 = _50282 ^ _1482;
  wire _50284 = _13389 ^ _50283;
  wire _50285 = _3811 ^ _23134;
  wire _50286 = _50285 ^ _4544;
  wire _50287 = _50284 ^ _50286;
  wire _50288 = _657 ^ _8998;
  wire _50289 = _50288 ^ _36183;
  wire _50290 = _9564 ^ _1498;
  wire _50291 = _1501 ^ _14442;
  wire _50292 = _50290 ^ _50291;
  wire _50293 = _50289 ^ _50292;
  wire _50294 = _50287 ^ _50293;
  wire _50295 = _5273 ^ _677;
  wire _50296 = _41730 ^ _50295;
  wire _50297 = _11776 ^ _10103;
  wire _50298 = _50297 ^ _24506;
  wire _50299 = _50296 ^ _50298;
  wire _50300 = _19861 ^ _5950;
  wire _50301 = _50300 ^ _48333;
  wire _50302 = _3065 ^ _14457;
  wire _50303 = uncoded_block[1407] ^ uncoded_block[1412];
  wire _50304 = _50303 ^ _20347;
  wire _50305 = _50302 ^ _50304;
  wire _50306 = _50301 ^ _50305;
  wire _50307 = _50299 ^ _50306;
  wire _50308 = _50294 ^ _50307;
  wire _50309 = uncoded_block[1424] ^ uncoded_block[1428];
  wire _50310 = _9588 ^ _50309;
  wire _50311 = _27598 ^ _50310;
  wire _50312 = _1531 ^ _2313;
  wire _50313 = _9595 ^ _14469;
  wire _50314 = _50312 ^ _50313;
  wire _50315 = _50311 ^ _50314;
  wire _50316 = _5305 ^ _8450;
  wire _50317 = _3865 ^ _3088;
  wire _50318 = _50316 ^ _50317;
  wire _50319 = _9602 ^ _29519;
  wire _50320 = _42517 ^ _50319;
  wire _50321 = _50318 ^ _50320;
  wire _50322 = _50315 ^ _50321;
  wire _50323 = _10701 ^ _31294;
  wire _50324 = uncoded_block[1485] ^ uncoded_block[1489];
  wire _50325 = _12342 ^ _50324;
  wire _50326 = _50323 ^ _50325;
  wire _50327 = _49947 ^ _747;
  wire _50328 = _15515 ^ _4616;
  wire _50329 = _50327 ^ _50328;
  wire _50330 = _50326 ^ _50329;
  wire _50331 = uncoded_block[1518] ^ uncoded_block[1524];
  wire _50332 = _50331 ^ _4623;
  wire _50333 = _4624 ^ _39050;
  wire _50334 = _50332 ^ _50333;
  wire _50335 = _6651 ^ _20387;
  wire _50336 = uncoded_block[1549] ^ uncoded_block[1552];
  wire _50337 = _16995 ^ _50336;
  wire _50338 = _50335 ^ _50337;
  wire _50339 = _50334 ^ _50338;
  wire _50340 = _50330 ^ _50339;
  wire _50341 = _50322 ^ _50340;
  wire _50342 = _50308 ^ _50341;
  wire _50343 = _50281 ^ _50342;
  wire _50344 = _769 ^ _10732;
  wire _50345 = _776 ^ _9072;
  wire _50346 = _50344 ^ _50345;
  wire _50347 = _6029 ^ _10171;
  wire _50348 = _17008 ^ _50347;
  wire _50349 = _50346 ^ _50348;
  wire _50350 = _9641 ^ _3935;
  wire _50351 = _3153 ^ _11303;
  wire _50352 = _12940 ^ _7297;
  wire _50353 = _50351 ^ _50352;
  wire _50354 = _50350 ^ _50353;
  wire _50355 = _50349 ^ _50354;
  wire _50356 = _7300 ^ _2400;
  wire _50357 = _31329 ^ _33852;
  wire _50358 = _50356 ^ _50357;
  wire _50359 = _3948 ^ _13500;
  wire _50360 = _24578 ^ _14011;
  wire _50361 = _50359 ^ _50360;
  wire _50362 = _50358 ^ _50361;
  wire _50363 = _3174 ^ _4687;
  wire _50364 = _24586 ^ _5406;
  wire _50365 = _50363 ^ _50364;
  wire _50366 = _17040 ^ _11324;
  wire _50367 = _7331 ^ _8527;
  wire _50368 = _50366 ^ _50367;
  wire _50369 = _50365 ^ _50368;
  wire _50370 = _50362 ^ _50369;
  wire _50371 = _50355 ^ _50370;
  wire _50372 = _11327 ^ _4700;
  wire _50373 = _847 ^ _11332;
  wire _50374 = _50372 ^ _50373;
  wire _50375 = _3201 ^ _7947;
  wire _50376 = _50374 ^ _50375;
  wire _50377 = _50371 ^ _50376;
  wire _50378 = _50343 ^ _50377;
  wire _50379 = _50217 ^ _50378;
  wire _50380 = _44790 ^ _27998;
  wire _50381 = _30035 ^ _50380;
  wire _50382 = _3224 ^ _6095;
  wire _50383 = _50382 ^ _7963;
  wire _50384 = _50381 ^ _50383;
  wire _50385 = _15591 ^ _6099;
  wire _50386 = _1705 ^ _34;
  wire _50387 = _50385 ^ _50386;
  wire _50388 = _897 ^ _2481;
  wire _50389 = _6755 ^ _15603;
  wire _50390 = _50388 ^ _50389;
  wire _50391 = _50387 ^ _50390;
  wire _50392 = _50384 ^ _50391;
  wire _50393 = _20952 ^ _4745;
  wire _50394 = _6762 ^ _2495;
  wire _50395 = _50393 ^ _50394;
  wire _50396 = _38721 ^ _4754;
  wire _50397 = _10820 ^ _50396;
  wire _50398 = _50395 ^ _50397;
  wire _50399 = _15112 ^ _64;
  wire _50400 = _10830 ^ _21901;
  wire _50401 = _50399 ^ _50400;
  wire _50402 = _71 ^ _3271;
  wire _50403 = uncoded_block[157] ^ uncoded_block[163];
  wire _50404 = uncoded_block[164] ^ uncoded_block[170];
  wire _50405 = _50403 ^ _50404;
  wire _50406 = _50402 ^ _50405;
  wire _50407 = _50401 ^ _50406;
  wire _50408 = _50398 ^ _50407;
  wire _50409 = _50392 ^ _50408;
  wire _50410 = _28037 ^ _4062;
  wire _50411 = _3283 ^ _2532;
  wire _50412 = _50410 ^ _50411;
  wire _50413 = _5486 ^ _97;
  wire _50414 = uncoded_block[211] ^ uncoded_block[219];
  wire _50415 = _50414 ^ _17617;
  wire _50416 = _50413 ^ _50415;
  wire _50417 = _50412 ^ _50416;
  wire _50418 = uncoded_block[226] ^ uncoded_block[232];
  wire _50419 = _50418 ^ _10289;
  wire _50420 = _8032 ^ _11954;
  wire _50421 = _50419 ^ _50420;
  wire _50422 = _1785 ^ _20023;
  wire _50423 = _6185 ^ _40341;
  wire _50424 = _50422 ^ _50423;
  wire _50425 = _50421 ^ _50424;
  wire _50426 = _50417 ^ _50425;
  wire _50427 = _44842 ^ _10303;
  wire _50428 = uncoded_block[283] ^ uncoded_block[291];
  wire _50429 = _5515 ^ _50428;
  wire _50430 = _50427 ^ _50429;
  wire _50431 = _13615 ^ _4111;
  wire _50432 = _6846 ^ _3340;
  wire _50433 = _50431 ^ _50432;
  wire _50434 = _50430 ^ _50433;
  wire _50435 = _18147 ^ _26021;
  wire _50436 = _28074 ^ _50435;
  wire _50437 = _18621 ^ _162;
  wire _50438 = _30994 ^ _50437;
  wire _50439 = _50436 ^ _50438;
  wire _50440 = _50434 ^ _50439;
  wire _50441 = _50426 ^ _50440;
  wire _50442 = _50409 ^ _50441;
  wire _50443 = _2601 ^ _6864;
  wire _50444 = _21955 ^ _16664;
  wire _50445 = _50443 ^ _50444;
  wire _50446 = uncoded_block[381] ^ uncoded_block[388];
  wire _50447 = _4143 ^ _50446;
  wire _50448 = _4152 ^ _1048;
  wire _50449 = _50447 ^ _50448;
  wire _50450 = _50445 ^ _50449;
  wire _50451 = _10341 ^ _44872;
  wire _50452 = _3394 ^ _19612;
  wire _50453 = _50451 ^ _50452;
  wire _50454 = _15197 ^ _14160;
  wire _50455 = _38788 ^ _14689;
  wire _50456 = _50454 ^ _50455;
  wire _50457 = _50453 ^ _50456;
  wire _50458 = _50450 ^ _50457;
  wire _50459 = _16187 ^ _206;
  wire _50460 = _16191 ^ _41909;
  wire _50461 = _50459 ^ _50460;
  wire _50462 = _2653 ^ _4185;
  wire _50463 = _1874 ^ _8686;
  wire _50464 = _50462 ^ _50463;
  wire _50465 = _50461 ^ _50464;
  wire _50466 = _49724 ^ _15212;
  wire _50467 = _7515 ^ _1093;
  wire _50468 = _50466 ^ _50467;
  wire _50469 = _6921 ^ _7529;
  wire _50470 = _26952 ^ _50469;
  wire _50471 = _50468 ^ _50470;
  wire _50472 = _50465 ^ _50471;
  wire _50473 = _50458 ^ _50472;
  wire _50474 = uncoded_block[514] ^ uncoded_block[519];
  wire _50475 = _6285 ^ _50474;
  wire _50476 = _1107 ^ _20602;
  wire _50477 = _50475 ^ _50476;
  wire _50478 = _4925 ^ _16215;
  wire _50479 = uncoded_block[548] ^ uncoded_block[555];
  wire _50480 = _10959 ^ _50479;
  wire _50481 = _50478 ^ _50480;
  wire _50482 = _50477 ^ _50481;
  wire _50483 = _1123 ^ _9319;
  wire _50484 = _5635 ^ _1931;
  wire _50485 = _50483 ^ _50484;
  wire _50486 = _13705 ^ _2701;
  wire _50487 = _46653 ^ _50486;
  wire _50488 = _50485 ^ _50487;
  wire _50489 = _50482 ^ _50488;
  wire _50490 = _19163 ^ _4240;
  wire _50491 = _50490 ^ _36432;
  wire _50492 = uncoded_block[616] ^ uncoded_block[621];
  wire _50493 = _50492 ^ _35228;
  wire _50494 = _5658 ^ _14228;
  wire _50495 = _50493 ^ _50494;
  wire _50496 = _50491 ^ _50495;
  wire _50497 = _5661 ^ _5665;
  wire _50498 = uncoded_block[641] ^ uncoded_block[646];
  wire _50499 = _50498 ^ _2730;
  wire _50500 = _50497 ^ _50499;
  wire _50501 = _40796 ^ _3515;
  wire _50502 = _50500 ^ _50501;
  wire _50503 = _50496 ^ _50502;
  wire _50504 = _50489 ^ _50503;
  wire _50505 = _50473 ^ _50504;
  wire _50506 = _50442 ^ _50505;
  wire _50507 = _1173 ^ _312;
  wire _50508 = _17745 ^ _12634;
  wire _50509 = _50507 ^ _50508;
  wire _50510 = _6983 ^ _325;
  wire _50511 = _22490 ^ _50510;
  wire _50512 = _50509 ^ _50511;
  wire _50513 = _326 ^ _3529;
  wire _50514 = _13740 ^ _6361;
  wire _50515 = _50513 ^ _50514;
  wire _50516 = uncoded_block[707] ^ uncoded_block[715];
  wire _50517 = _50516 ^ _4281;
  wire _50518 = uncoded_block[729] ^ uncoded_block[732];
  wire _50519 = _344 ^ _50518;
  wire _50520 = _50517 ^ _50519;
  wire _50521 = _50515 ^ _50520;
  wire _50522 = _50512 ^ _50521;
  wire _50523 = _5006 ^ _8775;
  wire _50524 = _3550 ^ _36873;
  wire _50525 = _50523 ^ _50524;
  wire _50526 = _43026 ^ _360;
  wire _50527 = _31542 ^ _12117;
  wire _50528 = _50526 ^ _50527;
  wire _50529 = _50525 ^ _50528;
  wire _50530 = _9384 ^ _5033;
  wire _50531 = _2799 ^ _6391;
  wire _50532 = _50530 ^ _50531;
  wire _50533 = _5039 ^ _12127;
  wire _50534 = _50533 ^ _22523;
  wire _50535 = _50532 ^ _50534;
  wire _50536 = _50529 ^ _50535;
  wire _50537 = _50522 ^ _50536;
  wire _50538 = _14802 ^ _5734;
  wire _50539 = _42380 ^ _50538;
  wire _50540 = uncoded_block[837] ^ uncoded_block[844];
  wire _50541 = _4331 ^ _50540;
  wire _50542 = _50541 ^ _40834;
  wire _50543 = _50539 ^ _50542;
  wire _50544 = _11048 ^ _413;
  wire _50545 = uncoded_block[875] ^ uncoded_block[882];
  wire _50546 = _5071 ^ _50545;
  wire _50547 = _50544 ^ _50546;
  wire _50548 = _17811 ^ _19735;
  wire _50549 = _5089 ^ _1281;
  wire _50550 = _50548 ^ _50549;
  wire _50551 = _50547 ^ _50550;
  wire _50552 = _50543 ^ _50551;
  wire _50553 = _25731 ^ _17820;
  wire _50554 = _1286 ^ _50553;
  wire _50555 = _31995 ^ _446;
  wire _50556 = _449 ^ _453;
  wire _50557 = _50555 ^ _50556;
  wire _50558 = _50554 ^ _50557;
  wire _50559 = _9433 ^ _11642;
  wire _50560 = _47863 ^ _9981;
  wire _50561 = _50559 ^ _50560;
  wire _50562 = _5113 ^ _37734;
  wire _50563 = _50561 ^ _50562;
  wire _50564 = _50558 ^ _50563;
  wire _50565 = _50552 ^ _50564;
  wire _50566 = _50537 ^ _50565;
  wire _50567 = uncoded_block[982] ^ uncoded_block[986];
  wire _50568 = _50567 ^ _8856;
  wire _50569 = _8859 ^ _19275;
  wire _50570 = _50568 ^ _50569;
  wire _50571 = _7691 ^ _22122;
  wire _50572 = _50571 ^ _32843;
  wire _50573 = _50570 ^ _50572;
  wire _50574 = _40113 ^ _45001;
  wire _50575 = uncoded_block[1035] ^ uncoded_block[1038];
  wire _50576 = _50575 ^ _512;
  wire _50577 = _50574 ^ _50576;
  wire _50578 = _7712 ^ _3682;
  wire _50579 = uncoded_block[1056] ^ uncoded_block[1061];
  wire _50580 = _50579 ^ _3685;
  wire _50581 = _50578 ^ _50580;
  wire _50582 = _50577 ^ _50581;
  wire _50583 = _50573 ^ _50582;
  wire _50584 = _2921 ^ _8892;
  wire _50585 = _5158 ^ _19301;
  wire _50586 = _50584 ^ _50585;
  wire _50587 = uncoded_block[1092] ^ uncoded_block[1096];
  wire _50588 = _8906 ^ _50587;
  wire _50589 = _43110 ^ _50588;
  wire _50590 = _50586 ^ _50589;
  wire _50591 = _13316 ^ _546;
  wire _50592 = _46063 ^ _4451;
  wire _50593 = _50591 ^ _50592;
  wire _50594 = _19313 ^ _3718;
  wire _50595 = _5854 ^ _14887;
  wire _50596 = _50594 ^ _50595;
  wire _50597 = _50593 ^ _50596;
  wire _50598 = _50590 ^ _50597;
  wire _50599 = _50583 ^ _50598;
  wire _50600 = uncoded_block[1138] ^ uncoded_block[1145];
  wire _50601 = _564 ^ _50600;
  wire _50602 = _27532 ^ _8937;
  wire _50603 = _50601 ^ _50602;
  wire _50604 = _2188 ^ _6511;
  wire _50605 = _5193 ^ _14901;
  wire _50606 = _50604 ^ _50605;
  wire _50607 = _50603 ^ _50606;
  wire _50608 = _5872 ^ _17892;
  wire _50609 = uncoded_block[1186] ^ uncoded_block[1196];
  wire _50610 = _4486 ^ _50609;
  wire _50611 = _50608 ^ _50610;
  wire _50612 = uncoded_block[1197] ^ uncoded_block[1204];
  wire _50613 = _50612 ^ _44674;
  wire _50614 = uncoded_block[1214] ^ uncoded_block[1225];
  wire _50615 = _2981 ^ _50614;
  wire _50616 = _50613 ^ _50615;
  wire _50617 = _50611 ^ _50616;
  wire _50618 = _50607 ^ _50617;
  wire _50619 = _1436 ^ _23548;
  wire _50620 = _50619 ^ _5222;
  wire _50621 = _11734 ^ _2232;
  wire _50622 = _6543 ^ _19358;
  wire _50623 = _50621 ^ _50622;
  wire _50624 = _50620 ^ _50623;
  wire _50625 = _12825 ^ _3003;
  wire _50626 = _50625 ^ _33763;
  wire _50627 = uncoded_block[1283] ^ uncoded_block[1292];
  wire _50628 = _50627 ^ _9547;
  wire _50629 = _19364 ^ _50628;
  wire _50630 = _50626 ^ _50629;
  wire _50631 = _50624 ^ _50630;
  wire _50632 = _50618 ^ _50631;
  wire _50633 = _50599 ^ _50632;
  wire _50634 = _50566 ^ _50633;
  wire _50635 = _50506 ^ _50634;
  wire _50636 = _31666 ^ _13918;
  wire _50637 = _3032 ^ _3820;
  wire _50638 = _38193 ^ _50637;
  wire _50639 = _50636 ^ _50638;
  wire _50640 = _3034 ^ _5261;
  wire _50641 = _7815 ^ _9003;
  wire _50642 = _50640 ^ _50641;
  wire _50643 = _5269 ^ _670;
  wire _50644 = uncoded_block[1354] ^ uncoded_block[1358];
  wire _50645 = _50644 ^ _6588;
  wire _50646 = _50643 ^ _50645;
  wire _50647 = _50642 ^ _50646;
  wire _50648 = _50639 ^ _50647;
  wire _50649 = uncoded_block[1361] ^ uncoded_block[1367];
  wire _50650 = _50649 ^ _24954;
  wire _50651 = _4564 ^ _3059;
  wire _50652 = _50650 ^ _50651;
  wire _50653 = _45074 ^ _4569;
  wire _50654 = _13938 ^ _12315;
  wire _50655 = _50653 ^ _50654;
  wire _50656 = _50652 ^ _50655;
  wire _50657 = _5296 ^ _33375;
  wire _50658 = _43559 ^ _50657;
  wire _50659 = _709 ^ _7844;
  wire _50660 = _50659 ^ _41356;
  wire _50661 = _50658 ^ _50660;
  wire _50662 = _50656 ^ _50661;
  wire _50663 = _50648 ^ _50662;
  wire _50664 = _2314 ^ _14469;
  wire _50665 = _20357 ^ _26763;
  wire _50666 = _50664 ^ _50665;
  wire _50667 = uncoded_block[1463] ^ uncoded_block[1470];
  wire _50668 = _3093 ^ _50667;
  wire _50669 = _47977 ^ _50668;
  wire _50670 = _50666 ^ _50669;
  wire _50671 = uncoded_block[1475] ^ uncoded_block[1493];
  wire _50672 = _50671 ^ _43955;
  wire _50673 = _47603 ^ _6637;
  wire _50674 = _50672 ^ _50673;
  wire _50675 = _7265 ^ _16988;
  wire _50676 = uncoded_block[1530] ^ uncoded_block[1536];
  wire _50677 = _1582 ^ _50676;
  wire _50678 = _50675 ^ _50677;
  wire _50679 = _50674 ^ _50678;
  wire _50680 = _50670 ^ _50679;
  wire _50681 = _6650 ^ _7274;
  wire _50682 = _50681 ^ _16502;
  wire _50683 = uncoded_block[1562] ^ uncoded_block[1568];
  wire _50684 = _4640 ^ _50683;
  wire _50685 = _7892 ^ _15535;
  wire _50686 = _50684 ^ _50685;
  wire _50687 = _50682 ^ _50686;
  wire _50688 = _1609 ^ _46487;
  wire _50689 = _12934 ^ _11292;
  wire _50690 = _50688 ^ _50689;
  wire _50691 = _8502 ^ _800;
  wire _50692 = uncoded_block[1613] ^ uncoded_block[1622];
  wire _50693 = _50692 ^ _5386;
  wire _50694 = _50691 ^ _50693;
  wire _50695 = _50690 ^ _50694;
  wire _50696 = _50687 ^ _50695;
  wire _50697 = _50680 ^ _50696;
  wire _50698 = _50663 ^ _50697;
  wire _50699 = _31749 ^ _20900;
  wire _50700 = _1642 ^ _6689;
  wire _50701 = _50699 ^ _50700;
  wire _50702 = _5394 ^ _819;
  wire _50703 = _50702 ^ _33009;
  wire _50704 = _50701 ^ _50703;
  wire _50705 = _3175 ^ _13511;
  wire _50706 = _25476 ^ _3183;
  wire _50707 = _50705 ^ _50706;
  wire _50708 = uncoded_block[1685] ^ uncoded_block[1692];
  wire _50709 = _5406 ^ _50708;
  wire _50710 = uncoded_block[1693] ^ uncoded_block[1712];
  wire _50711 = _50710 ^ _2441;
  wire _50712 = _50709 ^ _50711;
  wire _50713 = _50707 ^ _50712;
  wire _50714 = _50704 ^ _50713;
  wire _50715 = _50714 ^ uncoded_block[1722];
  wire _50716 = _50698 ^ _50715;
  wire _50717 = _50635 ^ _50716;
  wire _50718 = _4710 ^ _3212;
  wire _50719 = _4 ^ _15075;
  wire _50720 = _50718 ^ _50719;
  wire _50721 = _9692 ^ _1690;
  wire _50722 = _50721 ^ _22791;
  wire _50723 = _50720 ^ _50722;
  wire _50724 = uncoded_block[44] ^ uncoded_block[49];
  wire _50725 = _20457 ^ _50724;
  wire _50726 = _19969 ^ _50725;
  wire _50727 = _4014 ^ _38299;
  wire _50728 = _7364 ^ _9705;
  wire _50729 = _50727 ^ _50728;
  wire _50730 = _50726 ^ _50729;
  wire _50731 = _50723 ^ _50730;
  wire _50732 = _11357 ^ _7367;
  wire _50733 = _897 ^ _5443;
  wire _50734 = _50732 ^ _50733;
  wire _50735 = uncoded_block[83] ^ uncoded_block[93];
  wire _50736 = _50735 ^ _4026;
  wire _50737 = _50736 ^ _29608;
  wire _50738 = _50734 ^ _50737;
  wire _50739 = _33474 ^ _36309;
  wire _50740 = _914 ^ _54;
  wire _50741 = _9721 ^ _56;
  wire _50742 = _50740 ^ _50741;
  wire _50743 = _50739 ^ _50742;
  wire _50744 = _50738 ^ _50743;
  wire _50745 = _50731 ^ _50744;
  wire _50746 = _2502 ^ _22817;
  wire _50747 = _46173 ^ _927;
  wire _50748 = _50746 ^ _50747;
  wire _50749 = _18099 ^ _8000;
  wire _50750 = _9186 ^ _9188;
  wire _50751 = _50749 ^ _50750;
  wire _50752 = _50748 ^ _50751;
  wire _50753 = _16108 ^ _9737;
  wire _50754 = _15123 ^ _42607;
  wire _50755 = _5483 ^ _3284;
  wire _50756 = _50754 ^ _50755;
  wire _50757 = _50753 ^ _50756;
  wire _50758 = _50752 ^ _50757;
  wire _50759 = _16116 ^ _9745;
  wire _50760 = uncoded_block[204] ^ uncoded_block[213];
  wire _50761 = _6805 ^ _50760;
  wire _50762 = _50759 ^ _50761;
  wire _50763 = _8606 ^ _14105;
  wire _50764 = _50763 ^ _12486;
  wire _50765 = _50762 ^ _50764;
  wire _50766 = _8029 ^ _1778;
  wire _50767 = _27299 ^ _50766;
  wire _50768 = _4797 ^ _116;
  wire _50769 = _3309 ^ _13609;
  wire _50770 = _50768 ^ _50769;
  wire _50771 = _50767 ^ _50770;
  wire _50772 = _50765 ^ _50771;
  wire _50773 = _50758 ^ _50772;
  wire _50774 = _50745 ^ _50773;
  wire _50775 = _6831 ^ _7440;
  wire _50776 = _16636 ^ _10872;
  wire _50777 = _50775 ^ _50776;
  wire _50778 = _4103 ^ _4105;
  wire _50779 = _50778 ^ _36771;
  wire _50780 = _50777 ^ _50779;
  wire _50781 = _9776 ^ _1000;
  wire _50782 = _8055 ^ _21017;
  wire _50783 = _50781 ^ _50782;
  wire _50784 = _145 ^ _13624;
  wire _50785 = _3347 ^ _152;
  wire _50786 = _50784 ^ _50785;
  wire _50787 = _50783 ^ _50786;
  wire _50788 = _50780 ^ _50787;
  wire _50789 = _11444 ^ _4125;
  wire _50790 = _3352 ^ _41887;
  wire _50791 = _50789 ^ _50790;
  wire _50792 = _161 ^ _11990;
  wire _50793 = _3356 ^ _50792;
  wire _50794 = _50791 ^ _50793;
  wire _50795 = _6221 ^ _6227;
  wire _50796 = _4851 ^ _15183;
  wire _50797 = _50795 ^ _50796;
  wire _50798 = _8076 ^ _4140;
  wire _50799 = _8079 ^ _13101;
  wire _50800 = _50798 ^ _50799;
  wire _50801 = _50797 ^ _50800;
  wire _50802 = _50794 ^ _50801;
  wire _50803 = _50788 ^ _50802;
  wire _50804 = _31005 ^ _18633;
  wire _50805 = _10910 ^ _2623;
  wire _50806 = _50804 ^ _50805;
  wire _50807 = _34766 ^ _9266;
  wire _50808 = _31452 ^ _50807;
  wire _50809 = _50806 ^ _50808;
  wire _50810 = uncoded_block[416] ^ uncoded_block[424];
  wire _50811 = _50810 ^ _197;
  wire _50812 = uncoded_block[433] ^ uncoded_block[438];
  wire _50813 = _13115 ^ _50812;
  wire _50814 = _50811 ^ _50813;
  wire _50815 = _3408 ^ _9275;
  wire _50816 = _2645 ^ _1870;
  wire _50817 = _50815 ^ _50816;
  wire _50818 = _50814 ^ _50817;
  wire _50819 = _50809 ^ _50818;
  wire _50820 = _13127 ^ _13662;
  wire _50821 = _50820 ^ _35974;
  wire _50822 = _8687 ^ _17687;
  wire _50823 = _50821 ^ _50822;
  wire _50824 = _8115 ^ _3432;
  wire _50825 = _33149 ^ _50824;
  wire _50826 = _1887 ^ _4908;
  wire _50827 = _39595 ^ _50826;
  wire _50828 = _50825 ^ _50827;
  wire _50829 = _50823 ^ _50828;
  wire _50830 = _50819 ^ _50829;
  wire _50831 = _50803 ^ _50830;
  wire _50832 = _50774 ^ _50831;
  wire _50833 = _3439 ^ _4208;
  wire _50834 = uncoded_block[519] ^ uncoded_block[527];
  wire _50835 = _50834 ^ _4925;
  wire _50836 = _50833 ^ _50835;
  wire _50837 = _18208 ^ _14197;
  wire _50838 = _14198 ^ _244;
  wire _50839 = _50837 ^ _50838;
  wire _50840 = _50836 ^ _50839;
  wire _50841 = _246 ^ _25182;
  wire _50842 = _17710 ^ _19153;
  wire _50843 = _50841 ^ _50842;
  wire _50844 = _10399 ^ _265;
  wire _50845 = _9325 ^ _18222;
  wire _50846 = _50844 ^ _50845;
  wire _50847 = _50843 ^ _50846;
  wire _50848 = _50840 ^ _50847;
  wire _50849 = _8149 ^ _4953;
  wire _50850 = _28516 ^ _50849;
  wire _50851 = uncoded_block[602] ^ uncoded_block[606];
  wire _50852 = _50851 ^ _6323;
  wire _50853 = _50852 ^ _13712;
  wire _50854 = _50850 ^ _50853;
  wire _50855 = _4246 ^ _6966;
  wire _50856 = _34421 ^ _50855;
  wire _50857 = _290 ^ _3502;
  wire _50858 = _50857 ^ _28528;
  wire _50859 = _50856 ^ _50858;
  wire _50860 = _50854 ^ _50859;
  wire _50861 = _50848 ^ _50860;
  wire _50862 = _296 ^ _6973;
  wire _50863 = _12080 ^ _12630;
  wire _50864 = _50862 ^ _50863;
  wire _50865 = _4978 ^ _1177;
  wire _50866 = _8176 ^ _3521;
  wire _50867 = _50865 ^ _50866;
  wire _50868 = _50864 ^ _50867;
  wire _50869 = _1971 ^ _13194;
  wire _50870 = _50869 ^ _34035;
  wire _50871 = _19195 ^ _14250;
  wire _50872 = _19685 ^ _50871;
  wire _50873 = _50870 ^ _50872;
  wire _50874 = _50868 ^ _50873;
  wire _50875 = _14255 ^ _4996;
  wire _50876 = _4998 ^ _17266;
  wire _50877 = _50875 ^ _50876;
  wire _50878 = _1984 ^ _8198;
  wire _50879 = _6999 ^ _2768;
  wire _50880 = _50878 ^ _50879;
  wire _50881 = _50877 ^ _50880;
  wire _50882 = _4287 ^ _1206;
  wire _50883 = uncoded_block[738] ^ uncoded_block[746];
  wire _50884 = _50883 ^ _1210;
  wire _50885 = _50882 ^ _50884;
  wire _50886 = _4295 ^ _2003;
  wire _50887 = _4299 ^ _43792;
  wire _50888 = _50886 ^ _50887;
  wire _50889 = _50885 ^ _50888;
  wire _50890 = _50881 ^ _50889;
  wire _50891 = _50874 ^ _50890;
  wire _50892 = _50861 ^ _50891;
  wire _50893 = _13215 ^ _1221;
  wire _50894 = _50893 ^ _26146;
  wire _50895 = _5715 ^ _1224;
  wire _50896 = _12675 ^ _374;
  wire _50897 = _50895 ^ _50896;
  wire _50898 = _50894 ^ _50897;
  wire _50899 = uncoded_block[802] ^ uncoded_block[807];
  wire _50900 = _375 ^ _50899;
  wire _50901 = _5041 ^ _2806;
  wire _50902 = _50900 ^ _50901;
  wire _50903 = _5046 ^ _12131;
  wire _50904 = _3587 ^ _26160;
  wire _50905 = _50903 ^ _50904;
  wire _50906 = _50902 ^ _50905;
  wire _50907 = _50898 ^ _50906;
  wire _50908 = _15329 ^ _7049;
  wire _50909 = _22080 ^ _50908;
  wire _50910 = _14300 ^ _413;
  wire _50911 = _5071 ^ _416;
  wire _50912 = _50910 ^ _50911;
  wire _50913 = _50909 ^ _50912;
  wire _50914 = _11620 ^ _420;
  wire _50915 = _8820 ^ _2059;
  wire _50916 = _50914 ^ _50915;
  wire _50917 = _2061 ^ _3614;
  wire _50918 = _14829 ^ _2843;
  wire _50919 = _50917 ^ _50918;
  wire _50920 = _50916 ^ _50919;
  wire _50921 = _50913 ^ _50920;
  wire _50922 = _50907 ^ _50921;
  wire _50923 = _11062 ^ _16821;
  wire _50924 = _50923 ^ _40845;
  wire _50925 = uncoded_block[919] ^ uncoded_block[926];
  wire _50926 = _2852 ^ _50925;
  wire _50927 = _2857 ^ _3637;
  wire _50928 = _50926 ^ _50927;
  wire _50929 = _50924 ^ _50928;
  wire _50930 = uncoded_block[939] ^ uncoded_block[944];
  wire _50931 = _35688 ^ _50930;
  wire _50932 = _1302 ^ _12175;
  wire _50933 = _50931 ^ _50932;
  wire _50934 = _32422 ^ _36515;
  wire _50935 = _34095 ^ _50934;
  wire _50936 = _50933 ^ _50935;
  wire _50937 = _50929 ^ _50936;
  wire _50938 = _4390 ^ _5789;
  wire _50939 = _5790 ^ _8855;
  wire _50940 = _50938 ^ _50939;
  wire _50941 = _2102 ^ _1318;
  wire _50942 = _19275 ^ _32431;
  wire _50943 = _50941 ^ _50942;
  wire _50944 = _50940 ^ _50943;
  wire _50945 = _38930 ^ _27879;
  wire _50946 = _2894 ^ _9454;
  wire _50947 = _9455 ^ _4417;
  wire _50948 = _50946 ^ _50947;
  wire _50949 = _50945 ^ _50948;
  wire _50950 = _50944 ^ _50949;
  wire _50951 = _50937 ^ _50950;
  wire _50952 = _50922 ^ _50951;
  wire _50953 = _50892 ^ _50952;
  wire _50954 = _50832 ^ _50953;
  wire _50955 = uncoded_block[1037] ^ uncoded_block[1044];
  wire _50956 = _501 ^ _50955;
  wire _50957 = _8309 ^ _13846;
  wire _50958 = _50956 ^ _50957;
  wire _50959 = _2917 ^ _526;
  wire _50960 = _9474 ^ _50959;
  wire _50961 = _50958 ^ _50960;
  wire _50962 = _5156 ^ _2924;
  wire _50963 = _50962 ^ _23971;
  wire _50964 = _17866 ^ _19789;
  wire _50965 = _50963 ^ _50964;
  wire _50966 = _50961 ^ _50965;
  wire _50967 = _25318 ^ _546;
  wire _50968 = uncoded_block[1109] ^ uncoded_block[1117];
  wire _50969 = _50968 ^ _8920;
  wire _50970 = _50967 ^ _50969;
  wire _50971 = _12232 ^ _6499;
  wire _50972 = uncoded_block[1134] ^ uncoded_block[1138];
  wire _50973 = _560 ^ _50972;
  wire _50974 = _50971 ^ _50973;
  wire _50975 = _50970 ^ _50974;
  wire _50976 = _10597 ^ _15902;
  wire _50977 = _40144 ^ _50976;
  wire _50978 = _49869 ^ _578;
  wire _50979 = _32884 ^ _4476;
  wire _50980 = _50978 ^ _50979;
  wire _50981 = _50977 ^ _50980;
  wire _50982 = _50975 ^ _50981;
  wire _50983 = _50966 ^ _50982;
  wire _50984 = _37391 ^ _591;
  wire _50985 = _592 ^ _3746;
  wire _50986 = _2971 ^ _15431;
  wire _50987 = _50985 ^ _50986;
  wire _50988 = _50984 ^ _50987;
  wire _50989 = _2210 ^ _26694;
  wire _50990 = _50989 ^ _24914;
  wire _50991 = _38574 ^ _13357;
  wire _50992 = _50991 ^ _22643;
  wire _50993 = _50990 ^ _50992;
  wire _50994 = _50988 ^ _50993;
  wire _50995 = _3771 ^ _31231;
  wire _50996 = _50995 ^ _48303;
  wire _50997 = _11186 ^ _3002;
  wire _50998 = _50996 ^ _50997;
  wire _50999 = _3003 ^ _627;
  wire _51000 = _3008 ^ _49897;
  wire _51001 = _50999 ^ _51000;
  wire _51002 = uncoded_block[1276] ^ uncoded_block[1279];
  wire _51003 = _51002 ^ _6560;
  wire _51004 = _1468 ^ _5916;
  wire _51005 = _51003 ^ _51004;
  wire _51006 = _51001 ^ _51005;
  wire _51007 = _50998 ^ _51006;
  wire _51008 = _50994 ^ _51007;
  wire _51009 = _50983 ^ _51008;
  wire _51010 = _8991 ^ _3808;
  wire _51011 = _23569 ^ _51010;
  wire _51012 = _5919 ^ _9552;
  wire _51013 = _7805 ^ _656;
  wire _51014 = _51012 ^ _51013;
  wire _51015 = _51011 ^ _51014;
  wire _51016 = _28672 ^ _35781;
  wire _51017 = _4553 ^ _7815;
  wire _51018 = _4556 ^ _3826;
  wire _51019 = _51017 ^ _51018;
  wire _51020 = _51016 ^ _51019;
  wire _51021 = _51015 ^ _51020;
  wire _51022 = _16443 ^ _6590;
  wire _51023 = _10101 ^ _16449;
  wire _51024 = uncoded_block[1379] ^ uncoded_block[1381];
  wire _51025 = _15966 ^ _51024;
  wire _51026 = _51023 ^ _51025;
  wire _51027 = _51022 ^ _51026;
  wire _51028 = _3059 ^ _12867;
  wire _51029 = _51028 ^ _33795;
  wire _51030 = _9016 ^ _701;
  wire _51031 = _21316 ^ _51030;
  wire _51032 = _51029 ^ _51031;
  wire _51033 = _51027 ^ _51032;
  wire _51034 = _51021 ^ _51033;
  wire _51035 = _5961 ^ _15492;
  wire _51036 = _26301 ^ _9588;
  wire _51037 = _51035 ^ _51036;
  wire _51038 = _13429 ^ _1531;
  wire _51039 = _1533 ^ _1540;
  wire _51040 = _51038 ^ _51039;
  wire _51041 = _51037 ^ _51040;
  wire _51042 = _4590 ^ _5305;
  wire _51043 = _2322 ^ _3865;
  wire _51044 = _51042 ^ _51043;
  wire _51045 = _719 ^ _3089;
  wire _51046 = _3870 ^ _2336;
  wire _51047 = _51045 ^ _51046;
  wire _51048 = _51044 ^ _51047;
  wire _51049 = _51041 ^ _51048;
  wire _51050 = _16977 ^ _1555;
  wire _51051 = _14988 ^ _51050;
  wire _51052 = _12342 ^ _27184;
  wire _51053 = _51052 ^ _9045;
  wire _51054 = _51051 ^ _51053;
  wire _51055 = uncoded_block[1501] ^ uncoded_block[1508];
  wire _51056 = _51055 ^ _4617;
  wire _51057 = _9047 ^ _51056;
  wire _51058 = _9055 ^ _6643;
  wire _51059 = _51058 ^ _24993;
  wire _51060 = _51057 ^ _51059;
  wire _51061 = _51054 ^ _51060;
  wire _51062 = _51049 ^ _51061;
  wire _51063 = _51034 ^ _51062;
  wire _51064 = _51009 ^ _51063;
  wire _51065 = _6005 ^ _5348;
  wire _51066 = _9627 ^ _51065;
  wire _51067 = _7883 ^ _2367;
  wire _51068 = _8482 ^ _24094;
  wire _51069 = _51067 ^ _51068;
  wire _51070 = _51066 ^ _51069;
  wire _51071 = _776 ^ _5363;
  wire _51072 = _9080 ^ _46485;
  wire _51073 = _51071 ^ _51072;
  wire _51074 = _6031 ^ _25008;
  wire _51075 = _51074 ^ _10174;
  wire _51076 = _51073 ^ _51075;
  wire _51077 = _51070 ^ _51076;
  wire _51078 = uncoded_block[1601] ^ uncoded_block[1606];
  wire _51079 = _51078 ^ _5380;
  wire _51080 = _18504 ^ _51079;
  wire _51081 = _16031 ^ _29999;
  wire _51082 = _51081 ^ _43985;
  wire _51083 = _51080 ^ _51082;
  wire _51084 = _10754 ^ _3948;
  wire _51085 = _24121 ^ _51084;
  wire _51086 = _7312 ^ _24578;
  wire _51087 = uncoded_block[1653] ^ uncoded_block[1660];
  wire _51088 = _51087 ^ _3175;
  wire _51089 = _51086 ^ _51088;
  wire _51090 = _51085 ^ _51089;
  wire _51091 = _51083 ^ _51090;
  wire _51092 = _51077 ^ _51091;
  wire _51093 = _9666 ^ _7322;
  wire _51094 = _7323 ^ _11870;
  wire _51095 = _51093 ^ _51094;
  wire _51096 = uncoded_block[1695] ^ uncoded_block[1700];
  wire _51097 = _6066 ^ _51096;
  wire _51098 = _11873 ^ _51097;
  wire _51099 = _51095 ^ _51098;
  wire _51100 = uncoded_block[1707] ^ uncoded_block[1714];
  wire _51101 = _24137 ^ _51100;
  wire _51102 = _51101 ^ _23679;
  wire _51103 = _51102 ^ uncoded_block[1720];
  wire _51104 = _51099 ^ _51103;
  wire _51105 = _51092 ^ _51104;
  wire _51106 = _51064 ^ _51105;
  wire _51107 = _50954 ^ _51106;
  wire _51108 = _1683 ^ _6724;
  wire _51109 = _49999 ^ _1687;
  wire _51110 = _51108 ^ _51109;
  wire _51111 = _21865 ^ _40665;
  wire _51112 = _51110 ^ _51111;
  wire _51113 = _20941 ^ _23;
  wire _51114 = _19969 ^ _51113;
  wire _51115 = _10238 ^ _7969;
  wire _51116 = _19973 ^ _51115;
  wire _51117 = _51114 ^ _51116;
  wire _51118 = _51112 ^ _51117;
  wire _51119 = _6742 ^ _12435;
  wire _51120 = uncoded_block[70] ^ uncoded_block[78];
  wire _51121 = _16085 ^ _51120;
  wire _51122 = _51119 ^ _51121;
  wire _51123 = uncoded_block[84] ^ uncoded_block[90];
  wire _51124 = _51123 ^ _14591;
  wire _51125 = _39111 ^ _51124;
  wire _51126 = _51122 ^ _51125;
  wire _51127 = _6758 ^ _7986;
  wire _51128 = _17584 ^ _9720;
  wire _51129 = _51127 ^ _51128;
  wire _51130 = uncoded_block[116] ^ uncoded_block[121];
  wire _51131 = _10816 ^ _51130;
  wire _51132 = _51131 ^ _45564;
  wire _51133 = _51129 ^ _51132;
  wire _51134 = _51126 ^ _51133;
  wire _51135 = _51118 ^ _51134;
  wire _51136 = _8581 ^ _11918;
  wire _51137 = _20964 ^ _51136;
  wire _51138 = _33909 ^ _14082;
  wire _51139 = _932 ^ _21906;
  wire _51140 = _51138 ^ _51139;
  wire _51141 = _51137 ^ _51140;
  wire _51142 = _48071 ^ _29626;
  wire _51143 = _4062 ^ _19544;
  wire _51144 = _34715 ^ _51143;
  wire _51145 = _51142 ^ _51144;
  wire _51146 = _51141 ^ _51145;
  wire _51147 = uncoded_block[197] ^ uncoded_block[205];
  wire _51148 = _3284 ^ _51147;
  wire _51149 = uncoded_block[209] ^ uncoded_block[214];
  wire _51150 = _51149 ^ _6811;
  wire _51151 = _51148 ^ _51150;
  wire _51152 = _109 ^ _1775;
  wire _51153 = _25100 ^ _51152;
  wire _51154 = _51151 ^ _51153;
  wire _51155 = _28051 ^ _26433;
  wire _51156 = _116 ^ _13053;
  wire _51157 = _9761 ^ _10864;
  wire _51158 = _51156 ^ _51157;
  wire _51159 = _51155 ^ _51158;
  wire _51160 = _51154 ^ _51159;
  wire _51161 = _51146 ^ _51160;
  wire _51162 = _51135 ^ _51161;
  wire _51163 = _6831 ^ _127;
  wire _51164 = _2566 ^ _7445;
  wire _51165 = _51163 ^ _51164;
  wire _51166 = _3327 ^ _17635;
  wire _51167 = _11425 ^ _51166;
  wire _51168 = _51165 ^ _51167;
  wire _51169 = _12511 ^ _33949;
  wire _51170 = _145 ^ _152;
  wire _51171 = _12521 ^ _2586;
  wire _51172 = _51170 ^ _51171;
  wire _51173 = _51169 ^ _51172;
  wire _51174 = _51168 ^ _51173;
  wire _51175 = _10323 ^ _1021;
  wire _51176 = _10321 ^ _51175;
  wire _51177 = _16161 ^ _4132;
  wire _51178 = _6863 ^ _33119;
  wire _51179 = _51177 ^ _51178;
  wire _51180 = _51176 ^ _51179;
  wire _51181 = _8076 ^ _173;
  wire _51182 = _42932 ^ _51181;
  wire _51183 = _19599 ^ _4151;
  wire _51184 = _20058 ^ _51183;
  wire _51185 = _51182 ^ _51184;
  wire _51186 = _51180 ^ _51185;
  wire _51187 = _51174 ^ _51186;
  wire _51188 = _3384 ^ _181;
  wire _51189 = _41525 ^ _4867;
  wire _51190 = _51188 ^ _51189;
  wire _51191 = _11473 ^ _9266;
  wire _51192 = _4871 ^ _1059;
  wire _51193 = _51191 ^ _51192;
  wire _51194 = _51190 ^ _51193;
  wire _51195 = _24248 ^ _32297;
  wire _51196 = _19115 ^ _1864;
  wire _51197 = _51195 ^ _51196;
  wire _51198 = uncoded_block[456] ^ uncoded_block[462];
  wire _51199 = _2650 ^ _51198;
  wire _51200 = _47378 ^ _51199;
  wire _51201 = _51197 ^ _51200;
  wire _51202 = _51194 ^ _51201;
  wire _51203 = _10927 ^ _6906;
  wire _51204 = _1083 ^ _49724;
  wire _51205 = _51203 ^ _51204;
  wire _51206 = _4897 ^ _24727;
  wire _51207 = _51206 ^ _17202;
  wire _51208 = _51205 ^ _51207;
  wire _51209 = _10375 ^ _4908;
  wire _51210 = _3435 ^ _51209;
  wire _51211 = _4910 ^ _3444;
  wire _51212 = _26080 ^ _16711;
  wire _51213 = _51211 ^ _51212;
  wire _51214 = _51210 ^ _51213;
  wire _51215 = _51208 ^ _51214;
  wire _51216 = _51202 ^ _51215;
  wire _51217 = _51187 ^ _51216;
  wire _51218 = _51162 ^ _51217;
  wire _51219 = _24279 ^ _14198;
  wire _51220 = _20605 ^ _51219;
  wire _51221 = _4933 ^ _15236;
  wire _51222 = _6299 ^ _51221;
  wire _51223 = _51220 ^ _51222;
  wire _51224 = _1916 ^ _8725;
  wire _51225 = _51224 ^ _21557;
  wire _51226 = _25186 ^ _8731;
  wire _51227 = _11526 ^ _4946;
  wire _51228 = _51226 ^ _51227;
  wire _51229 = _51225 ^ _51228;
  wire _51230 = _51223 ^ _51229;
  wire _51231 = uncoded_block[586] ^ uncoded_block[590];
  wire _51232 = _51231 ^ _2700;
  wire _51233 = _15247 ^ _25640;
  wire _51234 = _51232 ^ _51233;
  wire _51235 = _2707 ^ _11535;
  wire _51236 = _51235 ^ _279;
  wire _51237 = _51234 ^ _51236;
  wire _51238 = _20125 ^ _12618;
  wire _51239 = _7565 ^ _51238;
  wire _51240 = _6966 ^ _43761;
  wire _51241 = _1161 ^ _16241;
  wire _51242 = _51240 ^ _51241;
  wire _51243 = _51239 ^ _51242;
  wire _51244 = _51237 ^ _51243;
  wire _51245 = _51230 ^ _51244;
  wire _51246 = _2729 ^ _35630;
  wire _51247 = _304 ^ _18705;
  wire _51248 = _51246 ^ _51247;
  wire _51249 = uncoded_block[665] ^ uncoded_block[671];
  wire _51250 = _4262 ^ _51249;
  wire _51251 = uncoded_block[672] ^ uncoded_block[676];
  wire _51252 = _51251 ^ _6352;
  wire _51253 = _51250 ^ _51252;
  wire _51254 = _51248 ^ _51253;
  wire _51255 = _12092 ^ _13740;
  wire _51256 = _34035 ^ _51255;
  wire _51257 = _6361 ^ _46294;
  wire _51258 = uncoded_block[718] ^ uncoded_block[725];
  wire _51259 = _10452 ^ _51258;
  wire _51260 = _51257 ^ _51259;
  wire _51261 = _51256 ^ _51260;
  wire _51262 = _51254 ^ _51261;
  wire _51263 = _11006 ^ _1206;
  wire _51264 = _4289 ^ _15301;
  wire _51265 = _51263 ^ _51264;
  wire _51266 = _21139 ^ _25685;
  wire _51267 = uncoded_block[761] ^ uncoded_block[767];
  wire _51268 = _3559 ^ _51267;
  wire _51269 = _51266 ^ _51268;
  wire _51270 = _51265 ^ _51269;
  wire _51271 = _7617 ^ _1221;
  wire _51272 = _31545 ^ _2794;
  wire _51273 = _51271 ^ _51272;
  wire _51274 = uncoded_block[784] ^ uncoded_block[790];
  wire _51275 = _51274 ^ _374;
  wire _51276 = uncoded_block[795] ^ uncoded_block[801];
  wire _51277 = _2799 ^ _51276;
  wire _51278 = _51275 ^ _51277;
  wire _51279 = _51273 ^ _51278;
  wire _51280 = _51270 ^ _51279;
  wire _51281 = _51262 ^ _51280;
  wire _51282 = _51245 ^ _51281;
  wire _51283 = _3577 ^ _1238;
  wire _51284 = _8228 ^ _11030;
  wire _51285 = _51283 ^ _51284;
  wire _51286 = _3587 ^ _24350;
  wire _51287 = _2030 ^ _51286;
  wire _51288 = _51285 ^ _51287;
  wire _51289 = _7043 ^ _8808;
  wire _51290 = _47457 ^ _51289;
  wire _51291 = _1257 ^ _7643;
  wire _51292 = _21165 ^ _5742;
  wire _51293 = _51291 ^ _51292;
  wire _51294 = _51290 ^ _51293;
  wire _51295 = _51288 ^ _51294;
  wire _51296 = _5069 ^ _2828;
  wire _51297 = _9953 ^ _11620;
  wire _51298 = _51296 ^ _51297;
  wire _51299 = _11621 ^ _35678;
  wire _51300 = _2061 ^ _1277;
  wire _51301 = _51299 ^ _51300;
  wire _51302 = _51298 ^ _51301;
  wire _51303 = _4361 ^ _3629;
  wire _51304 = _33684 ^ _7670;
  wire _51305 = _51303 ^ _51304;
  wire _51306 = _23914 ^ _51305;
  wire _51307 = _51302 ^ _51306;
  wire _51308 = _51295 ^ _51307;
  wire _51309 = _2084 ^ _2086;
  wire _51310 = _9975 ^ _4381;
  wire _51311 = _51309 ^ _51310;
  wire _51312 = _5779 ^ _5105;
  wire _51313 = _1310 ^ _10531;
  wire _51314 = _51312 ^ _51313;
  wire _51315 = _51311 ^ _51314;
  wire _51316 = _13821 ^ _5789;
  wire _51317 = _46738 ^ _51316;
  wire _51318 = _8856 ^ _12737;
  wire _51319 = _10538 ^ _51318;
  wire _51320 = _51317 ^ _51319;
  wire _51321 = _51315 ^ _51320;
  wire _51322 = _8293 ^ _2107;
  wire _51323 = _40109 ^ _2886;
  wire _51324 = _51322 ^ _51323;
  wire _51325 = _2890 ^ _9996;
  wire _51326 = uncoded_block[1019] ^ uncoded_block[1024];
  wire _51327 = _2893 ^ _51326;
  wire _51328 = _51325 ^ _51327;
  wire _51329 = _51324 ^ _51328;
  wire _51330 = uncoded_block[1027] ^ uncoded_block[1033];
  wire _51331 = _495 ^ _51330;
  wire _51332 = _51331 ^ _2131;
  wire _51333 = uncoded_block[1045] ^ uncoded_block[1056];
  wire _51334 = _51333 ^ _1363;
  wire _51335 = _4433 ^ _2917;
  wire _51336 = _51334 ^ _51335;
  wire _51337 = _51332 ^ _51336;
  wire _51338 = _51329 ^ _51337;
  wire _51339 = _51321 ^ _51338;
  wire _51340 = _51308 ^ _51339;
  wire _51341 = _51282 ^ _51340;
  wire _51342 = _51218 ^ _51341;
  wire _51343 = _2921 ^ _13851;
  wire _51344 = _2924 ^ _5162;
  wire _51345 = _51343 ^ _51344;
  wire _51346 = _3696 ^ _10021;
  wire _51347 = _25777 ^ _51346;
  wire _51348 = _51345 ^ _51347;
  wire _51349 = _11138 ^ _8332;
  wire _51350 = _550 ^ _552;
  wire _51351 = _51350 ^ _1390;
  wire _51352 = _51349 ^ _51351;
  wire _51353 = _51348 ^ _51352;
  wire _51354 = _13869 ^ _20269;
  wire _51355 = _47526 ^ _51354;
  wire _51356 = _46389 ^ _4466;
  wire _51357 = _4468 ^ _46391;
  wire _51358 = _51356 ^ _51357;
  wire _51359 = _51355 ^ _51358;
  wire _51360 = _13335 ^ _1408;
  wire _51361 = _16892 ^ _51360;
  wire _51362 = _1410 ^ _13339;
  wire _51363 = uncoded_block[1183] ^ uncoded_block[1191];
  wire _51364 = _31637 ^ _51363;
  wire _51365 = _51362 ^ _51364;
  wire _51366 = _51361 ^ _51365;
  wire _51367 = _51359 ^ _51366;
  wire _51368 = _51353 ^ _51367;
  wire _51369 = uncoded_block[1193] ^ uncoded_block[1199];
  wire _51370 = uncoded_block[1200] ^ uncoded_block[1205];
  wire _51371 = _51369 ^ _51370;
  wire _51372 = _51371 ^ _36983;
  wire _51373 = _12813 ^ _606;
  wire _51374 = _19347 ^ _612;
  wire _51375 = _51373 ^ _51374;
  wire _51376 = _51372 ^ _51375;
  wire _51377 = _1439 ^ _31228;
  wire _51378 = _2226 ^ _2230;
  wire _51379 = _51377 ^ _51378;
  wire _51380 = _23550 ^ _2997;
  wire _51381 = _51380 ^ _7779;
  wire _51382 = _51379 ^ _51381;
  wire _51383 = _51376 ^ _51382;
  wire _51384 = uncoded_block[1261] ^ uncoded_block[1270];
  wire _51385 = _12825 ^ _51384;
  wire _51386 = _1463 ^ _23123;
  wire _51387 = _51385 ^ _51386;
  wire _51388 = _638 ^ _11195;
  wire _51389 = _5916 ^ _4536;
  wire _51390 = _51388 ^ _51389;
  wire _51391 = _51387 ^ _51390;
  wire _51392 = _14430 ^ _1486;
  wire _51393 = _51392 ^ _20820;
  wire _51394 = _44316 ^ _4550;
  wire _51395 = uncoded_block[1336] ^ uncoded_block[1342];
  wire _51396 = _4551 ^ _51395;
  wire _51397 = _51394 ^ _51396;
  wire _51398 = _51393 ^ _51397;
  wire _51399 = _51391 ^ _51398;
  wire _51400 = _51383 ^ _51399;
  wire _51401 = _51368 ^ _51400;
  wire _51402 = _17938 ^ _15473;
  wire _51403 = _15477 ^ _5275;
  wire _51404 = _51402 ^ _51403;
  wire _51405 = _677 ^ _2289;
  wire _51406 = _5285 ^ _10108;
  wire _51407 = _51405 ^ _51406;
  wire _51408 = _51404 ^ _51407;
  wire _51409 = _17953 ^ _5952;
  wire _51410 = _13416 ^ _2299;
  wire _51411 = _51409 ^ _51410;
  wire _51412 = _43559 ^ _47587;
  wire _51413 = _51411 ^ _51412;
  wire _51414 = _51408 ^ _51413;
  wire _51415 = uncoded_block[1426] ^ uncoded_block[1431];
  wire _51416 = _51415 ^ _14978;
  wire _51417 = _51416 ^ _18913;
  wire _51418 = _46843 ^ _42513;
  wire _51419 = _51417 ^ _51418;
  wire _51420 = _7241 ^ _20361;
  wire _51421 = _51420 ^ _42519;
  wire _51422 = _23179 ^ _1558;
  wire _51423 = _22711 ^ _15510;
  wire _51424 = _51422 ^ _51423;
  wire _51425 = _51421 ^ _51424;
  wire _51426 = _51419 ^ _51425;
  wire _51427 = _51414 ^ _51426;
  wire _51428 = _1571 ^ _3894;
  wire _51429 = _7257 ^ _51428;
  wire _51430 = _4616 ^ _750;
  wire _51431 = _9055 ^ _7265;
  wire _51432 = _51430 ^ _51431;
  wire _51433 = _51429 ^ _51432;
  wire _51434 = _24993 ^ _16991;
  wire _51435 = uncoded_block[1533] ^ uncoded_block[1539];
  wire _51436 = _6002 ^ _51435;
  wire _51437 = _51436 ^ _51067;
  wire _51438 = _51434 ^ _51437;
  wire _51439 = _51433 ^ _51438;
  wire _51440 = _6013 ^ _3131;
  wire _51441 = _51440 ^ _43592;
  wire _51442 = uncoded_block[1565] ^ uncoded_block[1572];
  wire _51443 = _51442 ^ _6028;
  wire _51444 = _1609 ^ _11838;
  wire _51445 = _51443 ^ _51444;
  wire _51446 = _51441 ^ _51445;
  wire _51447 = _49119 ^ _46490;
  wire _51448 = _46491 ^ _16030;
  wire _51449 = _51447 ^ _51448;
  wire _51450 = _51446 ^ _51449;
  wire _51451 = _51439 ^ _51450;
  wire _51452 = _51427 ^ _51451;
  wire _51453 = _51401 ^ _51452;
  wire _51454 = _47635 ^ _11307;
  wire _51455 = _39847 ^ _51454;
  wire _51456 = uncoded_block[1636] ^ uncoded_block[1640];
  wire _51457 = _51456 ^ _13500;
  wire _51458 = _24121 ^ _51457;
  wire _51459 = _51455 ^ _51458;
  wire _51460 = _7312 ^ _3172;
  wire _51461 = _9106 ^ _12390;
  wire _51462 = _51460 ^ _51461;
  wire _51463 = _22761 ^ _4687;
  wire _51464 = _19939 ^ _11319;
  wire _51465 = _51463 ^ _51464;
  wire _51466 = _51462 ^ _51465;
  wire _51467 = _51459 ^ _51466;
  wire _51468 = uncoded_block[1680] ^ uncoded_block[1685];
  wire _51469 = _51468 ^ _3189;
  wire _51470 = uncoded_block[1693] ^ uncoded_block[1699];
  wire _51471 = _3190 ^ _51470;
  wire _51472 = _51469 ^ _51471;
  wire _51473 = _6068 ^ _22314;
  wire _51474 = _2438 ^ _854;
  wire _51475 = _51473 ^ _51474;
  wire _51476 = _51472 ^ _51475;
  wire _51477 = _51476 ^ _861;
  wire _51478 = _51467 ^ _51477;
  wire _51479 = _51453 ^ _51478;
  wire _51480 = _51342 ^ _51479;
  wire _51481 = _2454 ^ _46150;
  wire _51482 = _46148 ^ _51481;
  wire _51483 = _19963 ^ _11344;
  wire _51484 = _51483 ^ _26847;
  wire _51485 = _51482 ^ _51484;
  wire _51486 = _886 ^ _10238;
  wire _51487 = _38296 ^ _51486;
  wire _51488 = _901 ^ _6750;
  wire _51489 = _11356 ^ _51488;
  wire _51490 = _51487 ^ _51489;
  wire _51491 = _51485 ^ _51490;
  wire _51492 = _45555 ^ _41045;
  wire _51493 = _12447 ^ _7986;
  wire _51494 = _50 ^ _6769;
  wire _51495 = _51493 ^ _51494;
  wire _51496 = _51492 ^ _51495;
  wire _51497 = _6771 ^ _13017;
  wire _51498 = _51497 ^ _46174;
  wire _51499 = uncoded_block[147] ^ uncoded_block[155];
  wire _51500 = _51499 ^ _4764;
  wire _51501 = _48065 ^ _51500;
  wire _51502 = _51498 ^ _51501;
  wire _51503 = _51496 ^ _51502;
  wire _51504 = _51491 ^ _51503;
  wire _51505 = _2521 ^ _85;
  wire _51506 = _48071 ^ _51505;
  wire _51507 = uncoded_block[180] ^ uncoded_block[186];
  wire _51508 = _51507 ^ _18111;
  wire _51509 = _33077 ^ _18583;
  wire _51510 = _51508 ^ _51509;
  wire _51511 = _51506 ^ _51510;
  wire _51512 = _17112 ^ _6805;
  wire _51513 = _4070 ^ _10852;
  wire _51514 = _51512 ^ _51513;
  wire _51515 = _6811 ^ _104;
  wire _51516 = _20990 ^ _1775;
  wire _51517 = _51515 ^ _51516;
  wire _51518 = _51514 ^ _51517;
  wire _51519 = _51511 ^ _51518;
  wire _51520 = _26441 ^ _26000;
  wire _51521 = _13607 ^ _51520;
  wire _51522 = _46197 ^ _51521;
  wire _51523 = _44843 ^ _24211;
  wire _51524 = _48092 ^ _42917;
  wire _51525 = _51523 ^ _51524;
  wire _51526 = _51522 ^ _51525;
  wire _51527 = _51519 ^ _51526;
  wire _51528 = _51504 ^ _51527;
  wire _51529 = _8636 ^ _4111;
  wire _51530 = _1000 ^ _31847;
  wire _51531 = _51529 ^ _51530;
  wire _51532 = _145 ^ _5530;
  wire _51533 = _51532 ^ _11982;
  wire _51534 = _51531 ^ _51533;
  wire _51535 = _11983 ^ _4126;
  wire _51536 = _51535 ^ _6215;
  wire _51537 = _6217 ^ _18151;
  wire _51538 = _6220 ^ _2602;
  wire _51539 = _51537 ^ _51538;
  wire _51540 = _51536 ^ _51539;
  wire _51541 = _51534 ^ _51540;
  wire _51542 = _21030 ^ _1835;
  wire _51543 = _51542 ^ _50798;
  wire _51544 = _21504 ^ _49229;
  wire _51545 = _26474 ^ _51544;
  wire _51546 = _51543 ^ _51545;
  wire _51547 = _2625 ^ _16177;
  wire _51548 = uncoded_block[417] ^ uncoded_block[424];
  wire _51549 = _12547 ^ _51548;
  wire _51550 = _51547 ^ _51549;
  wire _51551 = _46234 ^ _35578;
  wire _51552 = _51550 ^ _51551;
  wire _51553 = _51546 ^ _51552;
  wire _51554 = _51541 ^ _51553;
  wire _51555 = _46239 ^ _46241;
  wire _51556 = _4186 ^ _4188;
  wire _51557 = _28493 ^ _51556;
  wire _51558 = _51555 ^ _51557;
  wire _51559 = uncoded_block[476] ^ uncoded_block[481];
  wire _51560 = _11494 ^ _51559;
  wire _51561 = _5598 ^ _12577;
  wire _51562 = _51560 ^ _51561;
  wire _51563 = _21536 ^ _13674;
  wire _51564 = _1095 ^ _51563;
  wire _51565 = _51562 ^ _51564;
  wire _51566 = _51558 ^ _51565;
  wire _51567 = _4908 ^ _23370;
  wire _51568 = _51567 ^ _48889;
  wire _51569 = _48892 ^ _15231;
  wire _51570 = _51568 ^ _51569;
  wire _51571 = _49268 ^ _3472;
  wire _51572 = _46260 ^ _51571;
  wire _51573 = _46259 ^ _51572;
  wire _51574 = _51570 ^ _51573;
  wire _51575 = _51566 ^ _51574;
  wire _51576 = _51554 ^ _51575;
  wire _51577 = _51528 ^ _51576;
  wire _51578 = _10399 ^ _15747;
  wire _51579 = _51578 ^ _48163;
  wire _51580 = _1939 ^ _4953;
  wire _51581 = _40409 ^ _51580;
  wire _51582 = _51579 ^ _51581;
  wire _51583 = _47041 ^ _19165;
  wire _51584 = uncoded_block[615] ^ uncoded_block[621];
  wire _51585 = _5652 ^ _51584;
  wire _51586 = _15261 ^ _1156;
  wire _51587 = _51585 ^ _51586;
  wire _51588 = _51583 ^ _51587;
  wire _51589 = _51582 ^ _51588;
  wire _51590 = _12075 ^ _5665;
  wire _51591 = _51590 ^ _14749;
  wire _51592 = _297 ^ _302;
  wire _51593 = _51592 ^ _36021;
  wire _51594 = _51591 ^ _51593;
  wire _51595 = _3514 ^ _10431;
  wire _51596 = _16752 ^ _21586;
  wire _51597 = _51595 ^ _51596;
  wire _51598 = _32764 ^ _1974;
  wire _51599 = uncoded_block[693] ^ uncoded_block[702];
  wire _51600 = _326 ^ _51599;
  wire _51601 = _51598 ^ _51600;
  wire _51602 = _51597 ^ _51601;
  wire _51603 = _51594 ^ _51602;
  wire _51604 = _51589 ^ _51603;
  wire _51605 = _51257 ^ _28171;
  wire _51606 = _6367 ^ _48933;
  wire _51607 = _51606 ^ _38862;
  wire _51608 = _51605 ^ _51607;
  wire _51609 = _33213 ^ _356;
  wire _51610 = _51609 ^ _46306;
  wire _51611 = _5019 ^ _365;
  wire _51612 = _51611 ^ _51271;
  wire _51613 = _51610 ^ _51612;
  wire _51614 = _51608 ^ _51613;
  wire _51615 = _49309 ^ _2019;
  wire _51616 = _14279 ^ _51615;
  wire _51617 = _4316 ^ _7629;
  wire _51618 = _1234 ^ _51617;
  wire _51619 = _51616 ^ _51618;
  wire _51620 = _1238 ^ _392;
  wire _51621 = uncoded_block[817] ^ uncoded_block[821];
  wire _51622 = _11030 ^ _51621;
  wire _51623 = _51620 ^ _51622;
  wire _51624 = _3587 ^ _12138;
  wire _51625 = _51624 ^ _47095;
  wire _51626 = _51623 ^ _51625;
  wire _51627 = _51619 ^ _51626;
  wire _51628 = _51614 ^ _51627;
  wire _51629 = _51604 ^ _51628;
  wire _51630 = _11609 ^ _1262;
  wire _51631 = _30680 ^ _5747;
  wire _51632 = _51630 ^ _51631;
  wire _51633 = _48222 ^ _46332;
  wire _51634 = _51632 ^ _51633;
  wire _51635 = _11621 ^ _2058;
  wire _51636 = _51635 ^ _50917;
  wire _51637 = _5085 ^ _5759;
  wire _51638 = _1280 ^ _7070;
  wire _51639 = _51637 ^ _51638;
  wire _51640 = _51636 ^ _51639;
  wire _51641 = _51634 ^ _51640;
  wire _51642 = _46723 ^ _438;
  wire _51643 = _51642 ^ _51304;
  wire _51644 = _48235 ^ _45368;
  wire _51645 = _51643 ^ _51644;
  wire _51646 = _5783 ^ _11646;
  wire _51647 = _49344 ^ _51646;
  wire _51648 = _8847 ^ _13821;
  wire _51649 = _471 ^ _10537;
  wire _51650 = _51648 ^ _51649;
  wire _51651 = _51647 ^ _51650;
  wire _51652 = _51645 ^ _51651;
  wire _51653 = _51641 ^ _51652;
  wire _51654 = _7093 ^ _8856;
  wire _51655 = _18333 ^ _5798;
  wire _51656 = _51654 ^ _51655;
  wire _51657 = _4409 ^ _5131;
  wire _51658 = _37740 ^ _51657;
  wire _51659 = _51656 ^ _51658;
  wire _51660 = _11663 ^ _7108;
  wire _51661 = _9455 ^ _30306;
  wire _51662 = _51660 ^ _51661;
  wire _51663 = _38937 ^ _46364;
  wire _51664 = _51663 ^ _21681;
  wire _51665 = _51662 ^ _51664;
  wire _51666 = _51659 ^ _51665;
  wire _51667 = _2924 ^ _20251;
  wire _51668 = _20753 ^ _20253;
  wire _51669 = _51667 ^ _51668;
  wire _51670 = _49849 ^ _51669;
  wire _51671 = _5840 ^ _5166;
  wire _51672 = _5169 ^ _15405;
  wire _51673 = _51671 ^ _51672;
  wire _51674 = uncoded_block[1109] ^ uncoded_block[1115];
  wire _51675 = _51674 ^ _1388;
  wire _51676 = uncoded_block[1127] ^ uncoded_block[1134];
  wire _51677 = _14376 ^ _51676;
  wire _51678 = _51675 ^ _51677;
  wire _51679 = _51673 ^ _51678;
  wire _51680 = _51670 ^ _51679;
  wire _51681 = _51666 ^ _51680;
  wire _51682 = _51653 ^ _51681;
  wire _51683 = _51629 ^ _51682;
  wire _51684 = _51577 ^ _51683;
  wire _51685 = _9496 ^ _46389;
  wire _51686 = _51685 ^ _34541;
  wire _51687 = _13335 ^ _9506;
  wire _51688 = _47532 ^ _51687;
  wire _51689 = _51686 ^ _51688;
  wire _51690 = _5872 ^ _4482;
  wire _51691 = _5200 ^ _49028;
  wire _51692 = _51690 ^ _51691;
  wire _51693 = _24910 ^ _2206;
  wire _51694 = _7163 ^ _49882;
  wire _51695 = _51693 ^ _51694;
  wire _51696 = _51692 ^ _51695;
  wire _51697 = _51689 ^ _51696;
  wire _51698 = _28298 ^ _32488;
  wire _51699 = uncoded_block[1233] ^ uncoded_block[1240];
  wire _51700 = _14919 ^ _51699;
  wire _51701 = _49399 ^ _51700;
  wire _51702 = _51698 ^ _51701;
  wire _51703 = _19829 ^ _8385;
  wire _51704 = _5231 ^ _32082;
  wire _51705 = _51703 ^ _51704;
  wire _51706 = _5234 ^ _34563;
  wire _51707 = _2239 ^ _3010;
  wire _51708 = _51706 ^ _51707;
  wire _51709 = _51705 ^ _51708;
  wire _51710 = _51702 ^ _51709;
  wire _51711 = _51697 ^ _51710;
  wire _51712 = _29468 ^ _16924;
  wire _51713 = _18866 ^ _642;
  wire _51714 = _51712 ^ _51713;
  wire _51715 = _23131 ^ _8407;
  wire _51716 = _39385 ^ _51715;
  wire _51717 = _51714 ^ _51716;
  wire _51718 = _49909 ^ _43163;
  wire _51719 = _5260 ^ _43922;
  wire _51720 = _51718 ^ _51719;
  wire _51721 = _51717 ^ _51720;
  wire _51722 = _21303 ^ _23581;
  wire _51723 = _51722 ^ _33365;
  wire _51724 = uncoded_block[1365] ^ uncoded_block[1369];
  wire _51725 = _51724 ^ _2289;
  wire _51726 = _7824 ^ _10108;
  wire _51727 = _51725 ^ _51726;
  wire _51728 = _51723 ^ _51727;
  wire _51729 = _46446 ^ _9015;
  wire _51730 = _5955 ^ _2299;
  wire _51731 = _51730 ^ _48340;
  wire _51732 = _51729 ^ _51731;
  wire _51733 = _51728 ^ _51732;
  wire _51734 = _51721 ^ _51733;
  wire _51735 = _51711 ^ _51734;
  wire _51736 = uncoded_block[1411] ^ uncoded_block[1421];
  wire _51737 = _51736 ^ _1527;
  wire _51738 = _15498 ^ _2314;
  wire _51739 = _51737 ^ _51738;
  wire _51740 = _45085 ^ _2322;
  wire _51741 = _21785 ^ _51740;
  wire _51742 = _51739 ^ _51741;
  wire _51743 = uncoded_block[1452] ^ uncoded_block[1461];
  wire _51744 = _3865 ^ _51743;
  wire _51745 = _51744 ^ _17973;
  wire _51746 = uncoded_block[1474] ^ uncoded_block[1478];
  wire _51747 = _1550 ^ _51746;
  wire _51748 = _12342 ^ _739;
  wire _51749 = _51747 ^ _51748;
  wire _51750 = _51745 ^ _51749;
  wire _51751 = _51742 ^ _51750;
  wire _51752 = _740 ^ _13967;
  wire _51753 = _51752 ^ _7257;
  wire _51754 = _5333 ^ _9055;
  wire _51755 = _49098 ^ _51754;
  wire _51756 = _51753 ^ _51755;
  wire _51757 = _9058 ^ _2357;
  wire _51758 = _51757 ^ _49459;
  wire _51759 = _39050 ^ _1589;
  wire _51760 = _32972 ^ _51759;
  wire _51761 = _51758 ^ _51760;
  wire _51762 = _51756 ^ _51761;
  wire _51763 = _51751 ^ _51762;
  wire _51764 = _48368 ^ _48370;
  wire _51765 = _15022 ^ _2376;
  wire _51766 = _5363 ^ _10163;
  wire _51767 = _51765 ^ _51766;
  wire _51768 = _51764 ^ _51767;
  wire _51769 = _3145 ^ _2394;
  wire _51770 = _50688 ^ _51769;
  wire _51771 = _13486 ^ _5373;
  wire _51772 = _51771 ^ _40994;
  wire _51773 = _51770 ^ _51772;
  wire _51774 = _51768 ^ _51773;
  wire _51775 = _4662 ^ _29997;
  wire _51776 = _18020 ^ _7912;
  wire _51777 = _51775 ^ _51776;
  wire _51778 = _46497 ^ _19929;
  wire _51779 = _12949 ^ _7309;
  wire _51780 = _51778 ^ _51779;
  wire _51781 = _51777 ^ _51780;
  wire _51782 = _7921 ^ _10757;
  wire _51783 = _51782 ^ _4679;
  wire _51784 = _10760 ^ _12960;
  wire _51785 = _3180 ^ _6059;
  wire _51786 = _51784 ^ _51785;
  wire _51787 = _51783 ^ _51786;
  wire _51788 = _51781 ^ _51787;
  wire _51789 = _51774 ^ _51788;
  wire _51790 = _51763 ^ _51789;
  wire _51791 = _51735 ^ _51790;
  wire _51792 = _35081 ^ _3189;
  wire _51793 = _51792 ^ _47648;
  wire _51794 = _3973 ^ _35477;
  wire _51795 = _51794 ^ _46519;
  wire _51796 = _51793 ^ _51795;
  wire _51797 = _51796 ^ _21402;
  wire _51798 = _51791 ^ _51797;
  wire _51799 = _51684 ^ _51798;
  wire _51800 = _19963 ^ _14565;
  wire _51801 = _49152 ^ _19501;
  wire _51802 = _51800 ^ _51801;
  wire _51803 = _51482 ^ _51802;
  wire _51804 = uncoded_block[66] ^ uncoded_block[75];
  wire _51805 = _51804 ^ _2481;
  wire _51806 = _51119 ^ _51805;
  wire _51807 = _51487 ^ _51806;
  wire _51808 = _51803 ^ _51807;
  wire _51809 = _6755 ^ _41044;
  wire _51810 = _35502 ^ _51809;
  wire _51811 = _46167 ^ _20477;
  wire _51812 = _51810 ^ _51811;
  wire _51813 = _6769 ^ _13016;
  wire _51814 = _51813 ^ _49174;
  wire _51815 = _46173 ^ _6136;
  wire _51816 = _10830 ^ _51499;
  wire _51817 = _51815 ^ _51816;
  wire _51818 = _51814 ^ _51817;
  wire _51819 = _51812 ^ _51818;
  wire _51820 = _51808 ^ _51819;
  wire _51821 = _24182 ^ _39128;
  wire _51822 = _51821 ^ _46183;
  wire _51823 = _34715 ^ _4063;
  wire _51824 = _51822 ^ _51823;
  wire _51825 = _46185 ^ _46188;
  wire _51826 = _33082 ^ _3296;
  wire _51827 = _51826 ^ _14106;
  wire _51828 = _51825 ^ _51827;
  wire _51829 = _51824 ^ _51828;
  wire _51830 = _963 ^ _7422;
  wire _51831 = _10289 ^ _10860;
  wire _51832 = _51830 ^ _51831;
  wire _51833 = _32258 ^ _13607;
  wire _51834 = _51832 ^ _51833;
  wire _51835 = uncoded_block[271] ^ uncoded_block[278];
  wire _51836 = _985 ^ _51835;
  wire _51837 = _51520 ^ _51836;
  wire _51838 = _49687 ^ _17635;
  wire _51839 = _12507 ^ _51838;
  wire _51840 = _51837 ^ _51839;
  wire _51841 = _51834 ^ _51840;
  wire _51842 = _51829 ^ _51841;
  wire _51843 = _51820 ^ _51842;
  wire _51844 = _46206 ^ _13618;
  wire _51845 = _8642 ^ _1014;
  wire _51846 = _46212 ^ _51845;
  wire _51847 = _51844 ^ _51846;
  wire _51848 = _48105 ^ _6858;
  wire _51849 = _46219 ^ _49222;
  wire _51850 = _51848 ^ _51849;
  wire _51851 = _51847 ^ _51850;
  wire _51852 = _33119 ^ _40360;
  wire _51853 = _51852 ^ _22415;
  wire _51854 = _48114 ^ _4858;
  wire _51855 = _10907 ^ _3383;
  wire _51856 = _51854 ^ _51855;
  wire _51857 = _51853 ^ _51856;
  wire _51858 = _24701 ^ _5559;
  wire _51859 = _7487 ^ _4867;
  wire _51860 = _51858 ^ _51859;
  wire _51861 = uncoded_block[413] ^ uncoded_block[417];
  wire _51862 = _11473 ^ _51861;
  wire _51863 = _24248 ^ _13115;
  wire _51864 = _51862 ^ _51863;
  wire _51865 = _51860 ^ _51864;
  wire _51866 = _51857 ^ _51865;
  wire _51867 = _51851 ^ _51866;
  wire _51868 = _13117 ^ _205;
  wire _51869 = _51868 ^ _48878;
  wire _51870 = _212 ^ _4181;
  wire _51871 = _10362 ^ _1878;
  wire _51872 = _51870 ^ _51871;
  wire _51873 = _51869 ^ _51872;
  wire _51874 = _51559 ^ _5598;
  wire _51875 = _19127 ^ _51874;
  wire _51876 = _12577 ^ _1093;
  wire _51877 = _1094 ^ _228;
  wire _51878 = _51876 ^ _51877;
  wire _51879 = _51875 ^ _51878;
  wire _51880 = _51873 ^ _51879;
  wire _51881 = _1887 ^ _9294;
  wire _51882 = _4908 ^ _4208;
  wire _51883 = _51881 ^ _51882;
  wire _51884 = _8709 ^ _30173;
  wire _51885 = _51883 ^ _51884;
  wire _51886 = _8132 ^ _1117;
  wire _51887 = _48149 ^ _51886;
  wire _51888 = _46258 ^ _33594;
  wire _51889 = _51887 ^ _51888;
  wire _51890 = _51885 ^ _51889;
  wire _51891 = _51880 ^ _51890;
  wire _51892 = _51867 ^ _51891;
  wire _51893 = _51843 ^ _51892;
  wire _51894 = _8725 ^ _24745;
  wire _51895 = _51894 ^ _3473;
  wire _51896 = _31915 ^ _18222;
  wire _51897 = _51227 ^ _51896;
  wire _51898 = _51895 ^ _51897;
  wire _51899 = _3481 ^ _46272;
  wire _51900 = _8154 ^ _5652;
  wire _51901 = _14219 ^ _51900;
  wire _51902 = _51899 ^ _51901;
  wire _51903 = _51898 ^ _51902;
  wire _51904 = _51584 ^ _3499;
  wire _51905 = _7576 ^ _4249;
  wire _51906 = _51904 ^ _51905;
  wire _51907 = _48916 ^ _49285;
  wire _51908 = _51906 ^ _51907;
  wire _51909 = _51249 ^ _1178;
  wire _51910 = _3515 ^ _51909;
  wire _51911 = _43774 ^ _22965;
  wire _51912 = _51910 ^ _51911;
  wire _51913 = _51908 ^ _51912;
  wire _51914 = _51903 ^ _51913;
  wire _51915 = _4272 ^ _1975;
  wire _51916 = _51915 ^ _51257;
  wire _51917 = _28171 ^ _51606;
  wire _51918 = _51916 ^ _51917;
  wire _51919 = _38862 ^ _51609;
  wire _51920 = _5019 ^ _28933;
  wire _51921 = _46306 ^ _51920;
  wire _51922 = _51919 ^ _51921;
  wire _51923 = _51918 ^ _51922;
  wire _51924 = _51271 ^ _26146;
  wire _51925 = _12673 ^ _2019;
  wire _51926 = _51925 ^ _1234;
  wire _51927 = _51924 ^ _51926;
  wire _51928 = _30669 ^ _46315;
  wire _51929 = uncoded_block[810] ^ uncoded_block[814];
  wire _51930 = _51929 ^ _5046;
  wire _51931 = _12131 ^ _3587;
  wire _51932 = _51930 ^ _51931;
  wire _51933 = _51928 ^ _51932;
  wire _51934 = _51927 ^ _51933;
  wire _51935 = _51923 ^ _51934;
  wire _51936 = _51914 ^ _51935;
  wire _51937 = _401 ^ _2035;
  wire _51938 = _51937 ^ _17301;
  wire _51939 = _1257 ^ _49326;
  wire _51940 = _51939 ^ _5067;
  wire _51941 = _51938 ^ _51940;
  wire _51942 = _49330 ^ _2828;
  wire _51943 = _9412 ^ _3608;
  wire _51944 = _51942 ^ _51943;
  wire _51945 = _11056 ^ _3613;
  wire _51946 = _51945 ^ _47103;
  wire _51947 = _51944 ^ _51946;
  wire _51948 = _51941 ^ _51947;
  wire _51949 = _23913 ^ _51638;
  wire _51950 = _6428 ^ _5092;
  wire _51951 = _15350 ^ _16315;
  wire _51952 = _51950 ^ _51951;
  wire _51953 = _51949 ^ _51952;
  wire _51954 = _2857 ^ _46344;
  wire _51955 = _51954 ^ _9976;
  wire _51956 = _49826 ^ _20717;
  wire _51957 = _51955 ^ _51956;
  wire _51958 = _51953 ^ _51957;
  wire _51959 = _51948 ^ _51958;
  wire _51960 = _51646 ^ _38510;
  wire _51961 = _51316 ^ _26641;
  wire _51962 = _51960 ^ _51961;
  wire _51963 = _50941 ^ _33277;
  wire _51964 = _51323 ^ _47132;
  wire _51965 = _51963 ^ _51964;
  wire _51966 = _51962 ^ _51965;
  wire _51967 = _7108 ^ _9455;
  wire _51968 = _30303 ^ _51967;
  wire _51969 = _30306 ^ _12199;
  wire _51970 = uncoded_block[1049] ^ uncoded_block[1056];
  wire _51971 = _2910 ^ _51970;
  wire _51972 = _51969 ^ _51971;
  wire _51973 = _51968 ^ _51972;
  wire _51974 = _49005 ^ _10570;
  wire _51975 = _13851 ^ _2924;
  wire _51976 = _20251 ^ _10575;
  wire _51977 = _51975 ^ _51976;
  wire _51978 = _51974 ^ _51977;
  wire _51979 = _51973 ^ _51978;
  wire _51980 = _51966 ^ _51979;
  wire _51981 = _51959 ^ _51980;
  wire _51982 = _51936 ^ _51981;
  wire _51983 = _51893 ^ _51982;
  wire _51984 = _1373 ^ _10021;
  wire _51985 = _11137 ^ _1380;
  wire _51986 = _51984 ^ _51985;
  wire _51987 = _545 ^ _20761;
  wire _51988 = _10585 ^ _1388;
  wire _51989 = _51987 ^ _51988;
  wire _51990 = _51986 ^ _51989;
  wire _51991 = _13869 ^ _43121;
  wire _51992 = _48272 ^ _51991;
  wire _51993 = _27533 ^ _46392;
  wire _51994 = _51992 ^ _51993;
  wire _51995 = _51990 ^ _51994;
  wire _51996 = uncoded_block[1166] ^ uncoded_block[1170];
  wire _51997 = _3734 ^ _51996;
  wire _51998 = _1410 ^ _5872;
  wire _51999 = _51997 ^ _51998;
  wire _52000 = _4482 ^ _35354;
  wire _52001 = _52000 ^ _49392;
  wire _52002 = _51999 ^ _52001;
  wire _52003 = _2206 ^ _7163;
  wire _52004 = _52003 ^ _27122;
  wire _52005 = _606 ^ _19347;
  wire _52006 = _21720 ^ _52005;
  wire _52007 = _52004 ^ _52006;
  wire _52008 = _52002 ^ _52007;
  wire _52009 = _51995 ^ _52008;
  wire _52010 = _31228 ^ _31231;
  wire _52011 = _46409 ^ _52010;
  wire _52012 = _17911 ^ _7778;
  wire _52013 = _3780 ^ _7780;
  wire _52014 = _52012 ^ _52013;
  wire _52015 = _52011 ^ _52014;
  wire _52016 = _10071 ^ _46419;
  wire _52017 = _52016 ^ _51386;
  wire _52018 = _639 ^ _45826;
  wire _52019 = _52018 ^ _39385;
  wire _52020 = _52017 ^ _52019;
  wire _52021 = _52015 ^ _52020;
  wire _52022 = _1486 ^ _40190;
  wire _52023 = _51715 ^ _52022;
  wire _52024 = _44316 ^ _660;
  wire _52025 = _3034 ^ _7815;
  wire _52026 = _52024 ^ _52025;
  wire _52027 = _52023 ^ _52026;
  wire _52028 = _20327 ^ _10097;
  wire _52029 = _7821 ^ _677;
  wire _52030 = _52028 ^ _52029;
  wire _52031 = uncoded_block[1365] ^ uncoded_block[1374];
  wire _52032 = _52031 ^ _12305;
  wire _52033 = _32935 ^ _6596;
  wire _52034 = _52032 ^ _52033;
  wire _52035 = _52030 ^ _52034;
  wire _52036 = _52027 ^ _52035;
  wire _52037 = _52021 ^ _52036;
  wire _52038 = _52009 ^ _52037;
  wire _52039 = _1513 ^ _5952;
  wire _52040 = _52039 ^ _46447;
  wire _52041 = _2300 ^ _3849;
  wire _52042 = _46449 ^ _52041;
  wire _52043 = _52040 ^ _52042;
  wire _52044 = _51736 ^ _24058;
  wire _52045 = _52044 ^ _51738;
  wire _52046 = _45085 ^ _3084;
  wire _52047 = _21785 ^ _52046;
  wire _52048 = _52045 ^ _52047;
  wire _52049 = _52043 ^ _52048;
  wire _52050 = _51743 ^ _2336;
  wire _52051 = _3866 ^ _52050;
  wire _52052 = _733 ^ _3100;
  wire _52053 = _42519 ^ _52052;
  wire _52054 = _52051 ^ _52053;
  wire _52055 = _19887 ^ _2349;
  wire _52056 = _52055 ^ _39039;
  wire _52057 = _45099 ^ _28370;
  wire _52058 = _52056 ^ _52057;
  wire _52059 = _52054 ^ _52058;
  wire _52060 = _52049 ^ _52059;
  wire _52061 = _19429 ^ _11267;
  wire _52062 = _52061 ^ _24993;
  wire _52063 = _16991 ^ _21349;
  wire _52064 = _52062 ^ _52063;
  wire _52065 = _7274 ^ _13472;
  wire _52066 = _49461 ^ _52065;
  wire _52067 = _22731 ^ _4638;
  wire _52068 = _26794 ^ _2376;
  wire _52069 = _52067 ^ _52068;
  wire _52070 = _52066 ^ _52069;
  wire _52071 = _52064 ^ _52070;
  wire _52072 = _16020 ^ _1609;
  wire _52073 = _46487 ^ _25454;
  wire _52074 = _52072 ^ _52073;
  wire _52075 = _37878 ^ _1626;
  wire _52076 = _52074 ^ _52075;
  wire _52077 = _3154 ^ _16031;
  wire _52078 = _52077 ^ _806;
  wire _52079 = _46497 ^ _5388;
  wire _52080 = _18965 ^ _3948;
  wire _52081 = _52079 ^ _52080;
  wire _52082 = _52078 ^ _52081;
  wire _52083 = _52076 ^ _52082;
  wire _52084 = _52071 ^ _52083;
  wire _52085 = _52060 ^ _52084;
  wire _52086 = _52038 ^ _52085;
  wire _52087 = _13501 ^ _17029;
  wire _52088 = uncoded_block[1663] ^ uncoded_block[1668];
  wire _52089 = _52088 ^ _19939;
  wire _52090 = _25024 ^ _52089;
  wire _52091 = _52087 ^ _52090;
  wire _52092 = _11319 ^ _35081;
  wire _52093 = _52092 ^ _3191;
  wire _52094 = _6066 ^ _3973;
  wire _52095 = _35477 ^ _7335;
  wire _52096 = _52094 ^ _52095;
  wire _52097 = _52093 ^ _52096;
  wire _52098 = _52091 ^ _52097;
  wire _52099 = _41018 ^ uncoded_block[1721];
  wire _52100 = _52098 ^ _52099;
  wire _52101 = _52086 ^ _52100;
  wire _52102 = _51983 ^ _52101;
  wire _52103 = _51483 ^ _19969;
  wire _52104 = _51482 ^ _52103;
  wire _52105 = uncoded_block[43] ^ uncoded_block[51];
  wire _52106 = _3230 ^ _52105;
  wire _52107 = _52106 ^ _49159;
  wire _52108 = _12435 ^ _51804;
  wire _52109 = _52108 ^ _51488;
  wire _52110 = _52107 ^ _52109;
  wire _52111 = _52104 ^ _52110;
  wire _52112 = _12451 ^ _1730;
  wire _52113 = _52112 ^ _925;
  wire _52114 = _2510 ^ _11918;
  wire _52115 = _33909 ^ _932;
  wire _52116 = _52114 ^ _52115;
  wire _52117 = _52113 ^ _52116;
  wire _52118 = _51496 ^ _52117;
  wire _52119 = _52111 ^ _52118;
  wire _52120 = _8591 ^ _48823;
  wire _52121 = _16108 ^ _52120;
  wire _52122 = _49186 ^ _48077;
  wire _52123 = _52121 ^ _52122;
  wire _52124 = _10278 ^ _33082;
  wire _52125 = _48078 ^ _52124;
  wire _52126 = _52125 ^ _51517;
  wire _52127 = _52123 ^ _52126;
  wire _52128 = _51836 ^ _12507;
  wire _52129 = uncoded_block[290] ^ uncoded_block[295];
  wire _52130 = _49687 ^ _52129;
  wire _52131 = _52130 ^ _15162;
  wire _52132 = _52128 ^ _52131;
  wire _52133 = _51522 ^ _52132;
  wire _52134 = _52127 ^ _52133;
  wire _52135 = _52119 ^ _52134;
  wire _52136 = _31847 ^ _145;
  wire _52137 = _22400 ^ _52136;
  wire _52138 = _5530 ^ _152;
  wire _52139 = _52138 ^ _16153;
  wire _52140 = _52137 ^ _52139;
  wire _52141 = _20544 ^ _30994;
  wire _52142 = _15686 ^ _40360;
  wire _52143 = _37980 ^ _52142;
  wire _52144 = _52141 ^ _52143;
  wire _52145 = _52140 ^ _52144;
  wire _52146 = _22415 ^ _51854;
  wire _52147 = _49229 ^ _2625;
  wire _52148 = _51855 ^ _52147;
  wire _52149 = _52146 ^ _52148;
  wire _52150 = _16177 ^ _12547;
  wire _52151 = _51548 ^ _14163;
  wire _52152 = _52150 ^ _52151;
  wire _52153 = _48126 ^ _49241;
  wire _52154 = _52152 ^ _52153;
  wire _52155 = _52149 ^ _52154;
  wire _52156 = _52145 ^ _52155;
  wire _52157 = _2650 ^ _9280;
  wire _52158 = _52157 ^ _27763;
  wire _52159 = _8687 ^ _9286;
  wire _52160 = _52158 ^ _52159;
  wire _52161 = _46246 ^ _24728;
  wire _52162 = _4905 ^ _1887;
  wire _52163 = _52162 ^ _13149;
  wire _52164 = _52161 ^ _52163;
  wire _52165 = _52160 ^ _52164;
  wire _52166 = _4208 ^ _8708;
  wire _52167 = _52166 ^ _46254;
  wire _52168 = _16711 ^ _1905;
  wire _52169 = _14197 ^ _8132;
  wire _52170 = _52168 ^ _52169;
  wire _52171 = _52167 ^ _52170;
  wire _52172 = _1909 ^ _1118;
  wire _52173 = _52172 ^ _43371;
  wire _52174 = _3472 ^ _10399;
  wire _52175 = _49269 ^ _52174;
  wire _52176 = _52173 ^ _52175;
  wire _52177 = _52171 ^ _52176;
  wire _52178 = _52165 ^ _52177;
  wire _52179 = _52156 ^ _52178;
  wire _52180 = _52135 ^ _52179;
  wire _52181 = _28513 ^ _51896;
  wire _52182 = _52181 ^ _51899;
  wire _52183 = _51584 ^ _15261;
  wire _52184 = _1156 ^ _12075;
  wire _52185 = _52183 ^ _52184;
  wire _52186 = _51901 ^ _52185;
  wire _52187 = _52182 ^ _52186;
  wire _52188 = _5665 ^ _4972;
  wire _52189 = _52188 ^ _298;
  wire _52190 = _6974 ^ _40030;
  wire _52191 = _52190 ^ _46283;
  wire _52192 = _52189 ^ _52191;
  wire _52193 = _21586 ^ _32764;
  wire _52194 = _21117 ^ _52193;
  wire _52195 = _51599 ^ _6361;
  wire _52196 = _34035 ^ _52195;
  wire _52197 = _52194 ^ _52196;
  wire _52198 = _52192 ^ _52197;
  wire _52199 = _52187 ^ _52198;
  wire _52200 = _46295 ^ _22972;
  wire _52201 = _1996 ^ _2774;
  wire _52202 = _48934 ^ _52201;
  wire _52203 = _52200 ^ _52202;
  wire _52204 = _1999 ^ _1210;
  wire _52205 = _52204 ^ _49788;
  wire _52206 = _43792 ^ _17776;
  wire _52207 = _52206 ^ _46309;
  wire _52208 = _52205 ^ _52207;
  wire _52209 = _52203 ^ _52208;
  wire _52210 = _368 ^ _3568;
  wire _52211 = _52210 ^ _51615;
  wire _52212 = _52211 ^ _51618;
  wire _52213 = _3587 ^ _401;
  wire _52214 = _52213 ^ _46322;
  wire _52215 = _51623 ^ _52214;
  wire _52216 = _52212 ^ _52215;
  wire _52217 = _52209 ^ _52216;
  wire _52218 = _52199 ^ _52217;
  wire _52219 = _8808 ^ _33239;
  wire _52220 = _2046 ^ _5066;
  wire _52221 = _52219 ^ _52220;
  wire _52222 = _3603 ^ _49330;
  wire _52223 = _2828 ^ _9412;
  wire _52224 = _52222 ^ _52223;
  wire _52225 = _52221 ^ _52224;
  wire _52226 = _17308 ^ _46336;
  wire _52227 = _8251 ^ _25728;
  wire _52228 = _52226 ^ _52227;
  wire _52229 = _52225 ^ _52228;
  wire _52230 = uncoded_block[910] ^ uncoded_block[914];
  wire _52231 = _2070 ^ _52230;
  wire _52232 = _438 ^ _33684;
  wire _52233 = _52231 ^ _52232;
  wire _52234 = _1302 ^ _5777;
  wire _52235 = _49341 ^ _52234;
  wire _52236 = _52233 ^ _52235;
  wire _52237 = _11646 ^ _1314;
  wire _52238 = _2877 ^ _5114;
  wire _52239 = _52237 ^ _52238;
  wire _52240 = _46349 ^ _52239;
  wire _52241 = _52236 ^ _52240;
  wire _52242 = _52229 ^ _52241;
  wire _52243 = _26641 ^ _50941;
  wire _52244 = _33277 ^ _51323;
  wire _52245 = _52243 ^ _52244;
  wire _52246 = _51657 ^ _51660;
  wire _52247 = _51661 ^ _51663;
  wire _52248 = _52246 ^ _52247;
  wire _52249 = _52245 ^ _52248;
  wire _52250 = _21681 ^ _3686;
  wire _52251 = _49848 ^ _51667;
  wire _52252 = _52250 ^ _52251;
  wire _52253 = _51668 ^ _51671;
  wire _52254 = _550 ^ _19313;
  wire _52255 = _51672 ^ _52254;
  wire _52256 = _52253 ^ _52255;
  wire _52257 = _52252 ^ _52256;
  wire _52258 = _52249 ^ _52257;
  wire _52259 = _52242 ^ _52258;
  wire _52260 = _52218 ^ _52259;
  wire _52261 = _52180 ^ _52260;
  wire _52262 = _51676 ^ _9496;
  wire _52263 = _49380 ^ _52262;
  wire _52264 = _46389 ^ _2185;
  wire _52265 = _8937 ^ _11711;
  wire _52266 = _52264 ^ _52265;
  wire _52267 = _52263 ^ _52266;
  wire _52268 = _2958 ^ _13335;
  wire _52269 = _9506 ^ _5872;
  wire _52270 = _52268 ^ _52269;
  wire _52271 = _10612 ^ _25805;
  wire _52272 = _52000 ^ _52271;
  wire _52273 = _52270 ^ _52272;
  wire _52274 = _52267 ^ _52273;
  wire _52275 = _23541 ^ _1429;
  wire _52276 = _6532 ^ _12819;
  wire _52277 = _31643 ^ _52276;
  wire _52278 = _52275 ^ _52277;
  wire _52279 = _31231 ^ _47551;
  wire _52280 = _51377 ^ _52279;
  wire _52281 = _7779 ^ _34564;
  wire _52282 = _52280 ^ _52281;
  wire _52283 = _52278 ^ _52282;
  wire _52284 = _52274 ^ _52283;
  wire _52285 = _51707 ^ _51712;
  wire _52286 = _51713 ^ _39385;
  wire _52287 = _52285 ^ _52286;
  wire _52288 = _51715 ^ _49909;
  wire _52289 = _20321 ^ _660;
  wire _52290 = _52289 ^ _46432;
  wire _52291 = _52288 ^ _52290;
  wire _52292 = _52287 ^ _52291;
  wire _52293 = _17938 ^ _37427;
  wire _52294 = _52293 ^ _46437;
  wire _52295 = _2289 ^ _7824;
  wire _52296 = _46438 ^ _52295;
  wire _52297 = _52294 ^ _52296;
  wire _52298 = _10108 ^ _11782;
  wire _52299 = _52298 ^ _48333;
  wire _52300 = _7226 ^ _29501;
  wire _52301 = _52299 ^ _52300;
  wire _52302 = _52297 ^ _52301;
  wire _52303 = _52292 ^ _52302;
  wire _52304 = _52284 ^ _52303;
  wire _52305 = _701 ^ _51736;
  wire _52306 = _52305 ^ _43945;
  wire _52307 = _52306 ^ _49443;
  wire _52308 = _42512 ^ _726;
  wire _52309 = _40962 ^ _52308;
  wire _52310 = _40603 ^ _2342;
  wire _52311 = _47599 ^ _52310;
  wire _52312 = _52309 ^ _52311;
  wire _52313 = _52307 ^ _52312;
  wire _52314 = _51748 ^ _51752;
  wire _52315 = _7257 ^ _49098;
  wire _52316 = _52314 ^ _52315;
  wire _52317 = _51754 ^ _51757;
  wire _52318 = _49459 ^ _32972;
  wire _52319 = _52317 ^ _52318;
  wire _52320 = _52316 ^ _52319;
  wire _52321 = _52313 ^ _52320;
  wire _52322 = _51759 ^ _48368;
  wire _52323 = _48370 ^ _51765;
  wire _52324 = _52322 ^ _52323;
  wire _52325 = _51766 ^ _50688;
  wire _52326 = _51769 ^ _51771;
  wire _52327 = _52325 ^ _52326;
  wire _52328 = _52324 ^ _52327;
  wire _52329 = _40994 ^ _51775;
  wire _52330 = _51776 ^ _52079;
  wire _52331 = _52329 ^ _52330;
  wire _52332 = _13500 ^ _6691;
  wire _52333 = _52080 ^ _52332;
  wire _52334 = _14011 ^ _2414;
  wire _52335 = _19463 ^ _52334;
  wire _52336 = _52333 ^ _52335;
  wire _52337 = _52331 ^ _52336;
  wire _52338 = _52328 ^ _52337;
  wire _52339 = _52321 ^ _52338;
  wire _52340 = _52304 ^ _52339;
  wire _52341 = _17032 ^ _2422;
  wire _52342 = _6059 ^ _35081;
  wire _52343 = _52341 ^ _52342;
  wire _52344 = _3191 ^ _52094;
  wire _52345 = _52343 ^ _52344;
  wire _52346 = _52095 ^ _41018;
  wire _52347 = _52346 ^ uncoded_block[1721];
  wire _52348 = _52345 ^ _52347;
  wire _52349 = _52340 ^ _52348;
  wire _52350 = _52261 ^ _52349;
  wire _52351 = _0 ^ _3212;
  wire _52352 = _52351 ^ _51481;
  wire _52353 = _1690 ^ _35096;
  wire _52354 = _11890 ^ _16;
  wire _52355 = _52353 ^ _52354;
  wire _52356 = _52352 ^ _52355;
  wire _52357 = _44419 ^ _51486;
  wire _52358 = _13552 ^ _12435;
  wire _52359 = _52358 ^ _33046;
  wire _52360 = _52357 ^ _52359;
  wire _52361 = _52356 ^ _52360;
  wire _52362 = _51488 ^ _31377;
  wire _52363 = _48807 ^ _34297;
  wire _52364 = _52362 ^ _52363;
  wire _52365 = _911 ^ _914;
  wire _52366 = _52365 ^ _46935;
  wire _52367 = _925 ^ _29199;
  wire _52368 = _52366 ^ _52367;
  wire _52369 = _52364 ^ _52368;
  wire _52370 = _52361 ^ _52369;
  wire _52371 = uncoded_block[149] ^ uncoded_block[155];
  wire _52372 = _18099 ^ _52371;
  wire _52373 = _24182 ^ _6785;
  wire _52374 = _52372 ^ _52373;
  wire _52375 = _4054 ^ _5473;
  wire _52376 = _2521 ^ _5476;
  wire _52377 = _52375 ^ _52376;
  wire _52378 = _52374 ^ _52377;
  wire _52379 = _5477 ^ _22368;
  wire _52380 = _52379 ^ _50755;
  wire _52381 = _52380 ^ _49669;
  wire _52382 = _52378 ^ _52381;
  wire _52383 = uncoded_block[205] ^ uncoded_block[215];
  wire _52384 = _52383 ^ _8606;
  wire _52385 = _52384 ^ _28799;
  wire _52386 = _11410 ^ _4081;
  wire _52387 = _52386 ^ _12489;
  wire _52388 = _52385 ^ _52387;
  wire _52389 = _16622 ^ _4797;
  wire _52390 = _116 ^ _3309;
  wire _52391 = _52389 ^ _52390;
  wire _52392 = _3311 ^ _26441;
  wire _52393 = _52392 ^ _10871;
  wire _52394 = _52391 ^ _52393;
  wire _52395 = _52388 ^ _52394;
  wire _52396 = _52382 ^ _52395;
  wire _52397 = _52370 ^ _52396;
  wire _52398 = uncoded_block[272] ^ uncoded_block[278];
  wire _52399 = _52398 ^ _1796;
  wire _52400 = _11428 ^ _135;
  wire _52401 = _52399 ^ _52400;
  wire _52402 = _49689 ^ _49691;
  wire _52403 = _52401 ^ _52402;
  wire _52404 = _6845 ^ _15668;
  wire _52405 = _145 ^ _6849;
  wire _52406 = _52404 ^ _52405;
  wire _52407 = _1821 ^ _5536;
  wire _52408 = _17152 ^ _52407;
  wire _52409 = _52406 ^ _52408;
  wire _52410 = _52403 ^ _52409;
  wire _52411 = _18151 ^ _30123;
  wire _52412 = _43325 ^ _52411;
  wire _52413 = _43705 ^ _8076;
  wire _52414 = _3363 ^ _52413;
  wire _52415 = _52412 ^ _52414;
  wire _52416 = _6873 ^ _13101;
  wire _52417 = _14677 ^ _3383;
  wire _52418 = _52416 ^ _52417;
  wire _52419 = _49229 ^ _7487;
  wire _52420 = _52419 ^ _14680;
  wire _52421 = _52418 ^ _52420;
  wire _52422 = _52415 ^ _52421;
  wire _52423 = _52410 ^ _52422;
  wire _52424 = _51191 ^ _52151;
  wire _52425 = uncoded_block[431] ^ uncoded_block[438];
  wire _52426 = _52425 ^ _3408;
  wire _52427 = _1864 ^ _1075;
  wire _52428 = _52426 ^ _52427;
  wire _52429 = _52424 ^ _52428;
  wire _52430 = _8686 ^ _221;
  wire _52431 = _52430 ^ _48137;
  wire _52432 = _51872 ^ _52431;
  wire _52433 = _52429 ^ _52432;
  wire _52434 = _24727 ^ _9837;
  wire _52435 = _52434 ^ _8702;
  wire _52436 = _1108 ^ _4921;
  wire _52437 = _49254 ^ _52436;
  wire _52438 = _52435 ^ _52437;
  wire _52439 = _52168 ^ _4928;
  wire _52440 = _8133 ^ _26085;
  wire _52441 = _52439 ^ _52440;
  wire _52442 = _52438 ^ _52441;
  wire _52443 = _52433 ^ _52442;
  wire _52444 = _52423 ^ _52443;
  wire _52445 = _52397 ^ _52444;
  wire _52446 = _8721 ^ _6940;
  wire _52447 = uncoded_block[569] ^ uncoded_block[575];
  wire _52448 = _2690 ^ _52447;
  wire _52449 = _52446 ^ _52448;
  wire _52450 = uncoded_block[583] ^ uncoded_block[590];
  wire _52451 = _4946 ^ _52450;
  wire _52452 = _15748 ^ _52451;
  wire _52453 = _52449 ^ _52452;
  wire _52454 = _2700 ^ _6316;
  wire _52455 = _52454 ^ _51580;
  wire _52456 = _2709 ^ _277;
  wire _52457 = _278 ^ _23400;
  wire _52458 = _52456 ^ _52457;
  wire _52459 = _52455 ^ _52458;
  wire _52460 = _52453 ^ _52459;
  wire _52461 = _16238 ^ _2719;
  wire _52462 = _6966 ^ _8161;
  wire _52463 = _52461 ^ _52462;
  wire _52464 = _17735 ^ _12077;
  wire _52465 = _52463 ^ _52464;
  wire _52466 = _40030 ^ _3514;
  wire _52467 = _25207 ^ _52466;
  wire _52468 = _51249 ^ _51251;
  wire _52469 = uncoded_block[686] ^ uncoded_block[690];
  wire _52470 = _23412 ^ _52469;
  wire _52471 = _52468 ^ _52470;
  wire _52472 = _52467 ^ _52471;
  wire _52473 = _52465 ^ _52472;
  wire _52474 = _52460 ^ _52473;
  wire _52475 = uncoded_block[693] ^ uncoded_block[699];
  wire _52476 = _326 ^ _52475;
  wire _52477 = _14250 ^ _11564;
  wire _52478 = _52476 ^ _52477;
  wire _52479 = _49778 ^ _342;
  wire _52480 = _52478 ^ _52479;
  wire _52481 = _27417 ^ _12104;
  wire _52482 = _34048 ^ _353;
  wire _52483 = _1210 ^ _5017;
  wire _52484 = _52482 ^ _52483;
  wire _52485 = _52481 ^ _52484;
  wire _52486 = _52480 ^ _52485;
  wire _52487 = _5020 ^ _17776;
  wire _52488 = _20162 ^ _52487;
  wire _52489 = _1221 ^ _14278;
  wire _52490 = _13219 ^ _12673;
  wire _52491 = _52489 ^ _52490;
  wire _52492 = _52488 ^ _52491;
  wire _52493 = _51276 ^ _5726;
  wire _52494 = _15806 ^ _52493;
  wire _52495 = _18755 ^ _48209;
  wire _52496 = _52494 ^ _52495;
  wire _52497 = _52492 ^ _52496;
  wire _52498 = _52486 ^ _52497;
  wire _52499 = _52474 ^ _52498;
  wire _52500 = uncoded_block[823] ^ uncoded_block[829];
  wire _52501 = _12131 ^ _52500;
  wire _52502 = _52501 ^ _34873;
  wire _52503 = _15329 ^ _2046;
  wire _52504 = _17301 ^ _52503;
  wire _52505 = _52502 ^ _52504;
  wire _52506 = uncoded_block[861] ^ uncoded_block[867];
  wire _52507 = _5066 ^ _52506;
  wire _52508 = _52507 ^ _52223;
  wire _52509 = _3608 ^ _4351;
  wire _52510 = _33249 ^ _14827;
  wire _52511 = _52509 ^ _52510;
  wire _52512 = _52508 ^ _52511;
  wire _52513 = _52505 ^ _52512;
  wire _52514 = _4355 ^ _1278;
  wire _52515 = _429 ^ _1280;
  wire _52516 = _52514 ^ _52515;
  wire _52517 = _16821 ^ _6428;
  wire _52518 = _5762 ^ _3629;
  wire _52519 = _52517 ^ _52518;
  wire _52520 = _52516 ^ _52519;
  wire _52521 = _2857 ^ _23475;
  wire _52522 = _3633 ^ _52521;
  wire _52523 = _2865 ^ _1302;
  wire _52524 = _52523 ^ _45368;
  wire _52525 = _52522 ^ _52524;
  wire _52526 = _52520 ^ _52525;
  wire _52527 = _52513 ^ _52526;
  wire _52528 = _4382 ^ _12726;
  wire _52529 = _11643 ^ _11646;
  wire _52530 = _52528 ^ _52529;
  wire _52531 = _15363 ^ _2877;
  wire _52532 = _5114 ^ _10537;
  wire _52533 = _52531 ^ _52532;
  wire _52534 = _52530 ^ _52533;
  wire _52535 = _23939 ^ _8293;
  wire _52536 = _51654 ^ _52535;
  wire _52537 = _5798 ^ _40109;
  wire _52538 = _2886 ^ _4409;
  wire _52539 = _52537 ^ _52538;
  wire _52540 = _52536 ^ _52539;
  wire _52541 = _52534 ^ _52540;
  wire _52542 = _26211 ^ _43854;
  wire _52543 = _27496 ^ _6474;
  wire _52544 = _29846 ^ _514;
  wire _52545 = _52543 ^ _52544;
  wire _52546 = _52542 ^ _52545;
  wire _52547 = _42039 ^ _12762;
  wire _52548 = _52547 ^ _42043;
  wire _52549 = _3689 ^ _21685;
  wire _52550 = _23502 ^ _52549;
  wire _52551 = _52548 ^ _52550;
  wire _52552 = _52546 ^ _52551;
  wire _52553 = _52541 ^ _52552;
  wire _52554 = _52527 ^ _52553;
  wire _52555 = _52499 ^ _52554;
  wire _52556 = _52445 ^ _52555;
  wire _52557 = uncoded_block[1076] ^ uncoded_block[1080];
  wire _52558 = _52557 ^ _10575;
  wire _52559 = _52558 ^ _49369;
  wire _52560 = _5840 ^ _33305;
  wire _52561 = _18365 ^ _19794;
  wire _52562 = _52560 ^ _52561;
  wire _52563 = _52559 ^ _52562;
  wire _52564 = _8339 ^ _5854;
  wire _52565 = _22154 ^ _52564;
  wire _52566 = _23523 ^ _14887;
  wire _52567 = _16380 ^ _46389;
  wire _52568 = _52566 ^ _52567;
  wire _52569 = _52565 ^ _52568;
  wire _52570 = _52563 ^ _52569;
  wire _52571 = _40149 ^ _47532;
  wire _52572 = _13339 ^ _4481;
  wire _52573 = _51687 ^ _52572;
  wire _52574 = _52571 ^ _52573;
  wire _52575 = _24910 ^ _11721;
  wire _52576 = _49029 ^ _52575;
  wire _52577 = _5207 ^ _1427;
  wire _52578 = _52577 ^ _21720;
  wire _52579 = _52576 ^ _52578;
  wire _52580 = _52574 ^ _52579;
  wire _52581 = _52570 ^ _52580;
  wire _52582 = _46406 ^ _46409;
  wire _52583 = _51699 ^ _19829;
  wire _52584 = _52583 ^ _39372;
  wire _52585 = _52582 ^ _52584;
  wire _52586 = _5232 ^ _40556;
  wire _52587 = _26271 ^ _45826;
  wire _52588 = _1464 ^ _52587;
  wire _52589 = _52586 ^ _52588;
  wire _52590 = _52585 ^ _52589;
  wire _52591 = uncoded_block[1293] ^ uncoded_block[1298];
  wire _52592 = _52591 ^ _8984;
  wire _52593 = _52592 ^ _46426;
  wire _52594 = _20816 ^ _21293;
  wire _52595 = _52594 ^ _34997;
  wire _52596 = _52593 ^ _52595;
  wire _52597 = _52024 ^ _46432;
  wire _52598 = _17938 ^ _10097;
  wire _52599 = _52598 ^ _35396;
  wire _52600 = _52597 ^ _52599;
  wire _52601 = _52596 ^ _52600;
  wire _52602 = _52590 ^ _52601;
  wire _52603 = _52581 ^ _52602;
  wire _52604 = _1504 ^ _6594;
  wire _52605 = _7824 ^ _11781;
  wire _52606 = _52604 ^ _52605;
  wire _52607 = _45074 ^ _5952;
  wire _52608 = _52607 ^ _46447;
  wire _52609 = _52606 ^ _52608;
  wire _52610 = _3066 ^ _3846;
  wire _52611 = _3847 ^ _3849;
  wire _52612 = _52610 ^ _52611;
  wire _52613 = _3069 ^ _3850;
  wire _52614 = _24058 ^ _5968;
  wire _52615 = _52613 ^ _52614;
  wire _52616 = _52612 ^ _52615;
  wire _52617 = _52609 ^ _52616;
  wire _52618 = _9591 ^ _2314;
  wire _52619 = _52618 ^ _21785;
  wire _52620 = _28354 ^ _5305;
  wire _52621 = _52620 ^ _51043;
  wire _52622 = _52619 ^ _52621;
  wire _52623 = _2326 ^ _2329;
  wire _52624 = _52623 ^ _18467;
  wire _52625 = _18919 ^ _733;
  wire _52626 = _35808 ^ _52625;
  wire _52627 = _52624 ^ _52626;
  wire _52628 = _52622 ^ _52627;
  wire _52629 = _52617 ^ _52628;
  wire _52630 = _7251 ^ _8462;
  wire _52631 = _24982 ^ _52630;
  wire _52632 = _52631 ^ _51429;
  wire _52633 = _4618 ^ _51058;
  wire _52634 = _24993 ^ _10720;
  wire _52635 = _52633 ^ _52634;
  wire _52636 = _52632 ^ _52635;
  wire _52637 = _39050 ^ _32975;
  wire _52638 = _32972 ^ _52637;
  wire _52639 = _16501 ^ _22731;
  wire _52640 = _7276 ^ _52639;
  wire _52641 = _52638 ^ _52640;
  wire _52642 = _24102 ^ _4647;
  wire _52643 = _19909 ^ _52642;
  wire _52644 = _3921 ^ _6031;
  wire _52645 = _52644 ^ _15032;
  wire _52646 = _52643 ^ _52645;
  wire _52647 = _52641 ^ _52646;
  wire _52648 = _52636 ^ _52647;
  wire _52649 = _52629 ^ _52648;
  wire _52650 = _52603 ^ _52649;
  wire _52651 = _11295 ^ _1624;
  wire _52652 = _46490 ^ _52651;
  wire _52653 = _29997 ^ _18020;
  wire _52654 = _44760 ^ _52653;
  wire _52655 = _52652 ^ _52654;
  wire _52656 = _33847 ^ _1639;
  wire _52657 = _812 ^ _51456;
  wire _52658 = _52656 ^ _52657;
  wire _52659 = _52658 ^ _52087;
  wire _52660 = _52655 ^ _52659;
  wire _52661 = _12960 ^ _5399;
  wire _52662 = _18032 ^ _52661;
  wire _52663 = _2422 ^ _830;
  wire _52664 = _52663 ^ _51792;
  wire _52665 = _52662 ^ _52664;
  wire _52666 = _3967 ^ _9675;
  wire _52667 = _32189 ^ _6068;
  wire _52668 = _52666 ^ _52667;
  wire _52669 = _1672 ^ _851;
  wire _52670 = _52669 ^ _41018;
  wire _52671 = _52668 ^ _52670;
  wire _52672 = _52665 ^ _52671;
  wire _52673 = _52660 ^ _52672;
  wire _52674 = _52673 ^ uncoded_block[1720];
  wire _52675 = _52650 ^ _52674;
  wire _52676 = _52556 ^ _52675;
  wire _52677 = _18539 ^ _4712;
  wire _52678 = _6724 ^ _3213;
  wire _52679 = _52677 ^ _52678;
  wire _52680 = _3219 ^ _2459;
  wire _52681 = _28748 ^ _52680;
  wire _52682 = _52679 ^ _52681;
  wire _52683 = _5429 ^ _6095;
  wire _52684 = uncoded_block[37] ^ uncoded_block[42];
  wire _52685 = _879 ^ _52684;
  wire _52686 = _52683 ^ _52685;
  wire _52687 = uncoded_block[48] ^ uncoded_block[60];
  wire _52688 = _4009 ^ _52687;
  wire _52689 = _13553 ^ _34;
  wire _52690 = _52688 ^ _52689;
  wire _52691 = _52686 ^ _52690;
  wire _52692 = _52682 ^ _52691;
  wire _52693 = uncoded_block[68] ^ uncoded_block[77];
  wire _52694 = _52693 ^ _28765;
  wire _52695 = _52694 ^ _17078;
  wire _52696 = _8568 ^ _14593;
  wire _52697 = _52695 ^ _52696;
  wire _52698 = _4031 ^ _20957;
  wire _52699 = _4034 ^ _54;
  wire _52700 = _52698 ^ _52699;
  wire _52701 = _10819 ^ _923;
  wire _52702 = _52701 ^ _11917;
  wire _52703 = _52700 ^ _52702;
  wire _52704 = _52697 ^ _52703;
  wire _52705 = _52692 ^ _52704;
  wire _52706 = _2511 ^ _8000;
  wire _52707 = _30066 ^ _52706;
  wire _52708 = _3271 ^ _73;
  wire _52709 = _52708 ^ _20976;
  wire _52710 = _52707 ^ _52709;
  wire _52711 = uncoded_block[170] ^ uncoded_block[175];
  wire _52712 = _6788 ^ _52711;
  wire _52713 = _52712 ^ _25981;
  wire _52714 = _14616 ^ _10277;
  wire _52715 = _6158 ^ _1764;
  wire _52716 = _52714 ^ _52715;
  wire _52717 = _52713 ^ _52716;
  wire _52718 = _52710 ^ _52717;
  wire _52719 = _29220 ^ _43297;
  wire _52720 = uncoded_block[235] ^ uncoded_block[240];
  wire _52721 = _2550 ^ _52720;
  wire _52722 = _10858 ^ _52721;
  wire _52723 = _52719 ^ _52722;
  wire _52724 = uncoded_block[241] ^ uncoded_block[248];
  wire _52725 = _52724 ^ _14116;
  wire _52726 = _11419 ^ _2559;
  wire _52727 = _52725 ^ _52726;
  wire _52728 = _10297 ^ _984;
  wire _52729 = uncoded_block[277] ^ uncoded_block[284];
  wire _52730 = _21479 ^ _52729;
  wire _52731 = _52728 ^ _52730;
  wire _52732 = _52727 ^ _52731;
  wire _52733 = _52723 ^ _52732;
  wire _52734 = _52718 ^ _52733;
  wire _52735 = _52705 ^ _52734;
  wire _52736 = _134 ^ _14128;
  wire _52737 = uncoded_block[307] ^ uncoded_block[311];
  wire _52738 = _14133 ^ _52737;
  wire _52739 = _52736 ^ _52738;
  wire _52740 = uncoded_block[326] ^ uncoded_block[331];
  wire _52741 = _13625 ^ _52740;
  wire _52742 = _32681 ^ _52741;
  wire _52743 = _52739 ^ _52742;
  wire _52744 = uncoded_block[340] ^ uncoded_block[345];
  wire _52745 = _6857 ^ _52744;
  wire _52746 = _1023 ^ _4132;
  wire _52747 = _52745 ^ _52746;
  wire _52748 = _162 ^ _36370;
  wire _52749 = _7470 ^ _3369;
  wire _52750 = _52748 ^ _52749;
  wire _52751 = _52747 ^ _52750;
  wire _52752 = _52743 ^ _52751;
  wire _52753 = _1838 ^ _10899;
  wire _52754 = _1038 ^ _3381;
  wire _52755 = _52753 ^ _52754;
  wire _52756 = uncoded_block[396] ^ uncoded_block[406];
  wire _52757 = _12541 ^ _52756;
  wire _52758 = _8091 ^ _13110;
  wire _52759 = _52757 ^ _52758;
  wire _52760 = _52755 ^ _52759;
  wire _52761 = _19613 ^ _4164;
  wire _52762 = _2633 ^ _201;
  wire _52763 = _52761 ^ _52762;
  wire _52764 = _5574 ^ _205;
  wire _52765 = _5580 ^ _3411;
  wire _52766 = _52764 ^ _52765;
  wire _52767 = _52763 ^ _52766;
  wire _52768 = _52760 ^ _52767;
  wire _52769 = _52752 ^ _52768;
  wire _52770 = _39197 ^ _3415;
  wire _52771 = _11491 ^ _3418;
  wire _52772 = _52770 ^ _52771;
  wire _52773 = _19127 ^ _21984;
  wire _52774 = _52772 ^ _52773;
  wire _52775 = _4895 ^ _8111;
  wire _52776 = _52775 ^ _43731;
  wire _52777 = _30605 ^ _13676;
  wire _52778 = _41544 ^ _52777;
  wire _52779 = _52776 ^ _52778;
  wire _52780 = _52774 ^ _52779;
  wire _52781 = uncoded_block[516] ^ uncoded_block[524];
  wire _52782 = _52781 ^ _4921;
  wire _52783 = _16711 ^ _9309;
  wire _52784 = _52782 ^ _52783;
  wire _52785 = uncoded_block[536] ^ uncoded_block[543];
  wire _52786 = uncoded_block[552] ^ uncoded_block[555];
  wire _52787 = _52785 ^ _52786;
  wire _52788 = _12051 ^ _9319;
  wire _52789 = _52787 ^ _52788;
  wire _52790 = _52784 ^ _52789;
  wire _52791 = _9320 ^ _1126;
  wire _52792 = _7550 ^ _4223;
  wire _52793 = _52791 ^ _52792;
  wire _52794 = uncoded_block[575] ^ uncoded_block[579];
  wire _52795 = _4224 ^ _52794;
  wire _52796 = _11527 ^ _8733;
  wire _52797 = _52795 ^ _52796;
  wire _52798 = _52793 ^ _52797;
  wire _52799 = _52790 ^ _52798;
  wire _52800 = _52780 ^ _52799;
  wire _52801 = _52769 ^ _52800;
  wire _52802 = _52735 ^ _52801;
  wire _52803 = _3478 ^ _2700;
  wire _52804 = _52803 ^ _13174;
  wire _52805 = _20626 ^ _5652;
  wire _52806 = _9335 ^ _52805;
  wire _52807 = _52804 ^ _52806;
  wire _52808 = _5653 ^ _20125;
  wire _52809 = _10979 ^ _17238;
  wire _52810 = _52808 ^ _52809;
  wire _52811 = _6969 ^ _40023;
  wire _52812 = _15763 ^ _52811;
  wire _52813 = _52810 ^ _52812;
  wire _52814 = _52807 ^ _52813;
  wire _52815 = _26112 ^ _3507;
  wire _52816 = _3514 ^ _9885;
  wire _52817 = _52815 ^ _52816;
  wire _52818 = _13731 ^ _319;
  wire _52819 = _3520 ^ _52818;
  wire _52820 = _52817 ^ _52819;
  wire _52821 = _3526 ^ _6983;
  wire _52822 = uncoded_block[689] ^ uncoded_block[694];
  wire _52823 = _52822 ^ _4989;
  wire _52824 = _52821 ^ _52823;
  wire _52825 = _334 ^ _4995;
  wire _52826 = _52825 ^ _36035;
  wire _52827 = _52824 ^ _52826;
  wire _52828 = _52820 ^ _52827;
  wire _52829 = _52814 ^ _52828;
  wire _52830 = _1983 ^ _340;
  wire _52831 = _30221 ^ _6374;
  wire _52832 = _52830 ^ _52831;
  wire _52833 = _10457 ^ _7605;
  wire _52834 = _1996 ^ _17272;
  wire _52835 = _52833 ^ _52834;
  wire _52836 = _52832 ^ _52835;
  wire _52837 = uncoded_block[750] ^ uncoded_block[763];
  wire _52838 = _3554 ^ _52837;
  wire _52839 = _13762 ^ _5027;
  wire _52840 = _52838 ^ _52839;
  wire _52841 = _33217 ^ _3562;
  wire _52842 = _52841 ^ _48582;
  wire _52843 = _52840 ^ _52842;
  wire _52844 = _52836 ^ _52843;
  wire _52845 = _8791 ^ _6391;
  wire _52846 = _48203 ^ _52845;
  wire _52847 = _7029 ^ _1235;
  wire _52848 = _52847 ^ _22523;
  wire _52849 = _52846 ^ _52848;
  wire _52850 = _4324 ^ _2029;
  wire _52851 = _52850 ^ _46705;
  wire _52852 = _2033 ^ _1253;
  wire _52853 = _5057 ^ _2820;
  wire _52854 = _52852 ^ _52853;
  wire _52855 = _52851 ^ _52854;
  wire _52856 = _52849 ^ _52855;
  wire _52857 = _52844 ^ _52856;
  wire _52858 = _52829 ^ _52857;
  wire _52859 = _8809 ^ _9945;
  wire _52860 = _5066 ^ _9949;
  wire _52861 = _52859 ^ _52860;
  wire _52862 = uncoded_block[873] ^ uncoded_block[877];
  wire _52863 = _52862 ^ _2053;
  wire _52864 = _20195 ^ _52863;
  wire _52865 = _52861 ^ _52864;
  wire _52866 = _12704 ^ _13251;
  wire _52867 = _21173 ^ _52866;
  wire _52868 = _15345 ^ _16312;
  wire _52869 = _21641 ^ _52868;
  wire _52870 = _52867 ^ _52869;
  wire _52871 = _52865 ^ _52870;
  wire _52872 = uncoded_block[914] ^ uncoded_block[920];
  wire _52873 = _52872 ^ _4370;
  wire _52874 = _10517 ^ _8839;
  wire _52875 = _52873 ^ _52874;
  wire _52876 = _8842 ^ _1310;
  wire _52877 = _13814 ^ _52876;
  wire _52878 = _52875 ^ _52877;
  wire _52879 = _11646 ^ _7088;
  wire _52880 = _38915 ^ _4391;
  wire _52881 = _52879 ^ _52880;
  wire _52882 = _8853 ^ _50567;
  wire _52883 = uncoded_block[987] ^ uncoded_block[995];
  wire _52884 = _52883 ^ _480;
  wire _52885 = _52882 ^ _52884;
  wire _52886 = _52881 ^ _52885;
  wire _52887 = _52878 ^ _52886;
  wire _52888 = _52871 ^ _52887;
  wire _52889 = _22122 ^ _2886;
  wire _52890 = uncoded_block[1008] ^ uncoded_block[1012];
  wire _52891 = _52890 ^ _2117;
  wire _52892 = _52889 ^ _52891;
  wire _52893 = _8299 ^ _5138;
  wire _52894 = _48252 ^ _52893;
  wire _52895 = _52892 ^ _52894;
  wire _52896 = _45001 ^ _1345;
  wire _52897 = _52896 ^ _11115;
  wire _52898 = _22135 ^ _1359;
  wire _52899 = _52898 ^ _17858;
  wire _52900 = _52897 ^ _52899;
  wire _52901 = _52895 ^ _52900;
  wire _52902 = _12213 ^ _12217;
  wire _52903 = _34932 ^ _52902;
  wire _52904 = _2148 ^ _30315;
  wire _52905 = _52903 ^ _52904;
  wire _52906 = uncoded_block[1088] ^ uncoded_block[1091];
  wire _52907 = _11687 ^ _52906;
  wire _52908 = _23071 ^ _545;
  wire _52909 = _52907 ^ _52908;
  wire _52910 = _19794 ^ _29426;
  wire _52911 = _8917 ^ _12782;
  wire _52912 = _52910 ^ _52911;
  wire _52913 = _52909 ^ _52912;
  wire _52914 = _52905 ^ _52913;
  wire _52915 = _52901 ^ _52914;
  wire _52916 = _52888 ^ _52915;
  wire _52917 = _52858 ^ _52916;
  wire _52918 = _52802 ^ _52917;
  wire _52919 = uncoded_block[1123] ^ uncoded_block[1128];
  wire _52920 = _5853 ^ _52919;
  wire _52921 = _4460 ^ _30329;
  wire _52922 = _52920 ^ _52921;
  wire _52923 = _18377 ^ _2185;
  wire _52924 = _3727 ^ _2958;
  wire _52925 = _52923 ^ _52924;
  wire _52926 = _52922 ^ _52925;
  wire _52927 = _2964 ^ _5193;
  wire _52928 = uncoded_block[1171] ^ uncoded_block[1174];
  wire _52929 = _52928 ^ _5872;
  wire _52930 = _52927 ^ _52929;
  wire _52931 = uncoded_block[1184] ^ uncoded_block[1190];
  wire _52932 = _592 ^ _52931;
  wire _52933 = _43886 ^ _52932;
  wire _52934 = _52930 ^ _52933;
  wire _52935 = _52926 ^ _52934;
  wire _52936 = _10612 ^ _5882;
  wire _52937 = _52936 ^ _14910;
  wire _52938 = _2982 ^ _2220;
  wire _52939 = _47172 ^ _52938;
  wire _52940 = _52937 ^ _52939;
  wire _52941 = _3766 ^ _1435;
  wire _52942 = _52941 ^ _29457;
  wire _52943 = _49401 ^ _6538;
  wire _52944 = _52943 ^ _31234;
  wire _52945 = _52942 ^ _52944;
  wire _52946 = _52940 ^ _52945;
  wire _52947 = _52935 ^ _52946;
  wire _52948 = _8388 ^ _1455;
  wire _52949 = _4514 ^ _9530;
  wire _52950 = _52948 ^ _52949;
  wire _52951 = uncoded_block[1266] ^ uncoded_block[1272];
  wire _52952 = _52951 ^ _631;
  wire _52953 = _52952 ^ _12275;
  wire _52954 = _52950 ^ _52953;
  wire _52955 = _43909 ^ _15947;
  wire _52956 = _21292 ^ _9555;
  wire _52957 = _41327 ^ _52956;
  wire _52958 = _52955 ^ _52957;
  wire _52959 = _52954 ^ _52958;
  wire _52960 = uncoded_block[1322] ^ uncoded_block[1331];
  wire _52961 = _52960 ^ _8413;
  wire _52962 = _52961 ^ _9565;
  wire _52963 = _5937 ^ _670;
  wire _52964 = _2280 ^ _1504;
  wire _52965 = _52963 ^ _52964;
  wire _52966 = _52962 ^ _52965;
  wire _52967 = _51724 ^ _3832;
  wire _52968 = _2290 ^ _18896;
  wire _52969 = _52967 ^ _52968;
  wire _52970 = _5950 ^ _4568;
  wire _52971 = _52970 ^ _46447;
  wire _52972 = _52969 ^ _52971;
  wire _52973 = _52966 ^ _52972;
  wire _52974 = _52959 ^ _52973;
  wire _52975 = _52947 ^ _52974;
  wire _52976 = _3066 ^ _16954;
  wire _52977 = _52976 ^ _2307;
  wire _52978 = _13429 ^ _14977;
  wire _52979 = _18456 ^ _52978;
  wire _52980 = _52977 ^ _52979;
  wire _52981 = _3857 ^ _24065;
  wire _52982 = _1535 ^ _52981;
  wire _52983 = _38626 ^ _1543;
  wire _52984 = _3088 ^ _3870;
  wire _52985 = _52983 ^ _52984;
  wire _52986 = _52982 ^ _52985;
  wire _52987 = _52980 ^ _52986;
  wire _52988 = _2336 ^ _10136;
  wire _52989 = _6627 ^ _1556;
  wire _52990 = _52988 ^ _52989;
  wire _52991 = _1558 ^ _50324;
  wire _52992 = _4610 ^ _25430;
  wire _52993 = _52991 ^ _52992;
  wire _52994 = _52990 ^ _52993;
  wire _52995 = uncoded_block[1500] ^ uncoded_block[1506];
  wire _52996 = _52995 ^ _4616;
  wire _52997 = _16488 ^ _9621;
  wire _52998 = _52996 ^ _52997;
  wire _52999 = _3118 ^ _6647;
  wire _53000 = _10150 ^ _52999;
  wire _53001 = _52998 ^ _53000;
  wire _53002 = _52994 ^ _53001;
  wire _53003 = _52987 ^ _53002;
  wire _53004 = _1586 ^ _1589;
  wire _53005 = _3129 ^ _22731;
  wire _53006 = _53004 ^ _53005;
  wire _53007 = _774 ^ _17007;
  wire _53008 = _31315 ^ _53007;
  wire _53009 = _53006 ^ _53008;
  wire _53010 = uncoded_block[1577] ^ uncoded_block[1588];
  wire _53011 = _4648 ^ _53010;
  wire _53012 = _53011 ^ _10174;
  wire _53013 = _33839 ^ _8502;
  wire _53014 = uncoded_block[1613] ^ uncoded_block[1619];
  wire _53015 = _3154 ^ _53014;
  wire _53016 = _53013 ^ _53015;
  wire _53017 = _53012 ^ _53016;
  wire _53018 = _53009 ^ _53017;
  wire _53019 = _6684 ^ _5386;
  wire _53020 = _808 ^ _7914;
  wire _53021 = _53019 ^ _53020;
  wire _53022 = _3169 ^ _36684;
  wire _53023 = _45903 ^ _53022;
  wire _53024 = _53021 ^ _53023;
  wire _53025 = uncoded_block[1649] ^ uncoded_block[1655];
  wire _53026 = uncoded_block[1658] ^ uncoded_block[1663];
  wire _53027 = _53025 ^ _53026;
  wire _53028 = _3179 ^ _5399;
  wire _53029 = _53027 ^ _53028;
  wire _53030 = _830 ^ _11321;
  wire _53031 = _12962 ^ _53030;
  wire _53032 = _53029 ^ _53031;
  wire _53033 = _53024 ^ _53032;
  wire _53034 = _53018 ^ _53033;
  wire _53035 = _53003 ^ _53034;
  wire _53036 = _52975 ^ _53035;
  wire _53037 = _17040 ^ _14543;
  wire _53038 = uncoded_block[1696] ^ uncoded_block[1701];
  wire _53039 = _18041 ^ _53038;
  wire _53040 = _53037 ^ _53039;
  wire _53041 = _44408 ^ _3200;
  wire _53042 = _45531 ^ _53041;
  wire _53043 = _53040 ^ _53042;
  wire _53044 = _2441 ^ _20923;
  wire _53045 = _53044 ^ uncoded_block[1720];
  wire _53046 = _53043 ^ _53045;
  wire _53047 = _53036 ^ _53046;
  wire _53048 = _52918 ^ _53047;
  wire _53049 = uncoded_block[5] ^ uncoded_block[9];
  wire _53050 = _1683 ^ _53049;
  wire _53051 = _15075 ^ _13537;
  wire _53052 = _53050 ^ _53051;
  wire _53053 = _44793 ^ _19969;
  wire _53054 = _53052 ^ _53053;
  wire _53055 = _20941 ^ _885;
  wire _53056 = _53055 ^ _51486;
  wire _53057 = _21881 ^ _4735;
  wire _53058 = _14581 ^ _53057;
  wire _53059 = _53056 ^ _53058;
  wire _53060 = _53054 ^ _53059;
  wire _53061 = _41044 ^ _1719;
  wire _53062 = _12441 ^ _53061;
  wire _53063 = _11911 ^ _32225;
  wire _53064 = _53062 ^ _53063;
  wire _53065 = _6769 ^ _12451;
  wire _53066 = _1730 ^ _923;
  wire _53067 = _53065 ^ _53066;
  wire _53068 = _33065 ^ _39515;
  wire _53069 = _53067 ^ _53068;
  wire _53070 = _53064 ^ _53069;
  wire _53071 = _53060 ^ _53070;
  wire _53072 = _4046 ^ _932;
  wire _53073 = _21906 ^ _4054;
  wire _53074 = _53072 ^ _53073;
  wire _53075 = uncoded_block[175] ^ uncoded_block[179];
  wire _53076 = _2521 ^ _53075;
  wire _53077 = _941 ^ _4062;
  wire _53078 = _53076 ^ _53077;
  wire _53079 = _53074 ^ _53078;
  wire _53080 = uncoded_block[189] ^ uncoded_block[194];
  wire _53081 = _53080 ^ _18583;
  wire _53082 = _53081 ^ _51512;
  wire _53083 = _4070 ^ _46189;
  wire _53084 = _8606 ^ _962;
  wire _53085 = _53083 ^ _53084;
  wire _53086 = _53082 ^ _53085;
  wire _53087 = _53079 ^ _53086;
  wire _53088 = _51830 ^ _5504;
  wire _53089 = _6180 ^ _39154;
  wire _53090 = _53089 ^ _33934;
  wire _53091 = _53088 ^ _53090;
  wire _53092 = _16636 ^ _9222;
  wire _53093 = _46199 ^ _53092;
  wire _53094 = uncoded_block[288] ^ uncoded_block[295];
  wire _53095 = _4105 ^ _53094;
  wire _53096 = _24211 ^ _53095;
  wire _53097 = _53093 ^ _53096;
  wire _53098 = _53091 ^ _53097;
  wire _53099 = _53087 ^ _53098;
  wire _53100 = _53071 ^ _53099;
  wire _53101 = _15162 ^ _22400;
  wire _53102 = _20536 ^ _4117;
  wire _53103 = _32274 ^ _13625;
  wire _53104 = _53102 ^ _53103;
  wire _53105 = _53101 ^ _53104;
  wire _53106 = _11982 ^ _51535;
  wire _53107 = _12526 ^ _11454;
  wire _53108 = _43325 ^ _53107;
  wire _53109 = _53106 ^ _53108;
  wire _53110 = _53105 ^ _53109;
  wire _53111 = _1028 ^ _2602;
  wire _53112 = _40360 ^ _19590;
  wire _53113 = _53111 ^ _53112;
  wire _53114 = _48114 ^ _6876;
  wire _53115 = _53114 ^ _51183;
  wire _53116 = _53113 ^ _53115;
  wire _53117 = _8661 ^ _181;
  wire _53118 = _2625 ^ _4867;
  wire _53119 = _53117 ^ _53118;
  wire _53120 = _11473 ^ _4871;
  wire _53121 = _53120 ^ _51863;
  wire _53122 = _53119 ^ _53121;
  wire _53123 = _53116 ^ _53122;
  wire _53124 = _53110 ^ _53123;
  wire _53125 = _10352 ^ _205;
  wire _53126 = _53125 ^ _39587;
  wire _53127 = _51870 ^ _51203;
  wire _53128 = _53126 ^ _53127;
  wire _53129 = _19127 ^ _15720;
  wire _53130 = _8694 ^ _35592;
  wire _53131 = _53130 ^ _5605;
  wire _53132 = _53129 ^ _53131;
  wire _53133 = _53128 ^ _53132;
  wire _53134 = _21536 ^ _12034;
  wire _53135 = _9294 ^ _11508;
  wire _53136 = _53134 ^ _53135;
  wire _53137 = _53136 ^ _51884;
  wire _53138 = _1118 ^ _3459;
  wire _53139 = _25631 ^ _4937;
  wire _53140 = _53138 ^ _53139;
  wire _53141 = _48150 ^ _53140;
  wire _53142 = _53137 ^ _53141;
  wire _53143 = _53133 ^ _53142;
  wire _53144 = _53124 ^ _53143;
  wire _53145 = _53100 ^ _53144;
  wire _53146 = _21555 ^ _24745;
  wire _53147 = _53146 ^ _47035;
  wire _53148 = _20116 ^ _9330;
  wire _53149 = _47405 ^ _53148;
  wire _53150 = _53147 ^ _53149;
  wire _53151 = _6316 ^ _25640;
  wire _53152 = _53151 ^ _7559;
  wire _53153 = _8154 ^ _8744;
  wire _53154 = _14219 ^ _53153;
  wire _53155 = _53152 ^ _53154;
  wire _53156 = _53150 ^ _53155;
  wire _53157 = _3499 ^ _7576;
  wire _53158 = _53157 ^ _46279;
  wire _53159 = _2729 ^ _6341;
  wire _53160 = _53159 ^ _36021;
  wire _53161 = _53158 ^ _53160;
  wire _53162 = _5670 ^ _312;
  wire _53163 = _19185 ^ _21586;
  wire _53164 = _53162 ^ _53163;
  wire _53165 = _34834 ^ _2754;
  wire _53166 = _2755 ^ _1188;
  wire _53167 = _53165 ^ _53166;
  wire _53168 = _53164 ^ _53167;
  wire _53169 = _53161 ^ _53168;
  wire _53170 = _53156 ^ _53169;
  wire _53171 = _11564 ^ _2762;
  wire _53172 = _10452 ^ _18726;
  wire _53173 = _53171 ^ _53172;
  wire _53174 = _46297 ^ _47068;
  wire _53175 = _1206 ^ _34048;
  wire _53176 = _53174 ^ _53175;
  wire _53177 = _53173 ^ _53176;
  wire _53178 = _25685 ^ _5019;
  wire _53179 = _18736 ^ _53178;
  wire _53180 = _2783 ^ _7617;
  wire _53181 = _53180 ^ _31105;
  wire _53182 = _53179 ^ _53181;
  wire _53183 = _53177 ^ _53182;
  wire _53184 = _52210 ^ _51275;
  wire _53185 = _4316 ^ _390;
  wire _53186 = _36474 ^ _53185;
  wire _53187 = _53184 ^ _53186;
  wire _53188 = uncoded_block[824] ^ uncoded_block[835];
  wire _53189 = _1241 ^ _53188;
  wire _53190 = _49316 ^ _53189;
  wire _53191 = _53190 ^ _46324;
  wire _53192 = _53187 ^ _53191;
  wire _53193 = _53183 ^ _53192;
  wire _53194 = _53170 ^ _53193;
  wire _53195 = _7643 ^ _8237;
  wire _53196 = _5747 ^ _13244;
  wire _53197 = _53195 ^ _53196;
  wire _53198 = uncoded_block[869] ^ uncoded_block[875];
  wire _53199 = _1266 ^ _53198;
  wire _53200 = _3608 ^ _2058;
  wire _53201 = _53199 ^ _53200;
  wire _53202 = _53197 ^ _53201;
  wire _53203 = _15345 ^ _2070;
  wire _53204 = _52230 ^ _3629;
  wire _53205 = _53203 ^ _53204;
  wire _53206 = _49336 ^ _53205;
  wire _53207 = _53202 ^ _53206;
  wire _53208 = _8259 ^ _31141;
  wire _53209 = uncoded_block[936] ^ uncoded_block[943];
  wire _53210 = _3637 ^ _53209;
  wire _53211 = _53208 ^ _53210;
  wire _53212 = _17829 ^ _52528;
  wire _53213 = _53211 ^ _53212;
  wire _53214 = _2871 ^ _1310;
  wire _53215 = _11646 ^ _15363;
  wire _53216 = _53214 ^ _53215;
  wire _53217 = _11089 ^ _8854;
  wire _53218 = _53216 ^ _53217;
  wire _53219 = _53213 ^ _53218;
  wire _53220 = _53207 ^ _53219;
  wire _53221 = _3659 ^ _8856;
  wire _53222 = _23939 ^ _479;
  wire _53223 = _53221 ^ _53222;
  wire _53224 = _20730 ^ _2886;
  wire _53225 = _25756 ^ _53224;
  wire _53226 = _53223 ^ _53225;
  wire _53227 = _47132 ^ _30303;
  wire _53228 = uncoded_block[1025] ^ uncoded_block[1028];
  wire _53229 = _7108 ^ _53228;
  wire _53230 = _30306 ^ _38937;
  wire _53231 = _53229 ^ _53230;
  wire _53232 = _53227 ^ _53231;
  wire _53233 = _53226 ^ _53232;
  wire _53234 = _46364 ^ _37755;
  wire _53235 = _1363 ^ _3684;
  wire _53236 = _53234 ^ _53235;
  wire _53237 = _527 ^ _2924;
  wire _53238 = _46370 ^ _53237;
  wire _53239 = _53236 ^ _53238;
  wire _53240 = _4440 ^ _5840;
  wire _53241 = _49010 ^ _53240;
  wire _53242 = uncoded_block[1100] ^ uncoded_block[1109];
  wire _53243 = _53242 ^ _10585;
  wire _53244 = _34527 ^ _53243;
  wire _53245 = _53241 ^ _53244;
  wire _53246 = _53239 ^ _53245;
  wire _53247 = _53233 ^ _53246;
  wire _53248 = _53220 ^ _53247;
  wire _53249 = _53194 ^ _53248;
  wire _53250 = _53145 ^ _53249;
  wire _53251 = _14376 ^ _23523;
  wire _53252 = _18830 ^ _53251;
  wire _53253 = _13866 ^ _13869;
  wire _53254 = _53253 ^ _38158;
  wire _53255 = _53252 ^ _53254;
  wire _53256 = _27533 ^ _47532;
  wire _53257 = _3736 ^ _1408;
  wire _53258 = _53257 ^ _48289;
  wire _53259 = _53256 ^ _53258;
  wire _53260 = _53255 ^ _53259;
  wire _53261 = _1417 ^ _9508;
  wire _53262 = _10612 ^ _14398;
  wire _53263 = _53261 ^ _53262;
  wire _53264 = _2216 ^ _18395;
  wire _53265 = _52003 ^ _53264;
  wire _53266 = _53263 ^ _53265;
  wire _53267 = _4498 ^ _606;
  wire _53268 = _19347 ^ _4504;
  wire _53269 = _53267 ^ _53268;
  wire _53270 = _31231 ^ _17911;
  wire _53271 = _49039 ^ _53270;
  wire _53272 = _53269 ^ _53271;
  wire _53273 = _53266 ^ _53272;
  wire _53274 = _53260 ^ _53273;
  wire _53275 = _8385 ^ _623;
  wire _53276 = _7780 ^ _2239;
  wire _53277 = _53275 ^ _53276;
  wire _53278 = _10075 ^ _2247;
  wire _53279 = _23123 ^ _639;
  wire _53280 = _53278 ^ _53279;
  wire _53281 = _53277 ^ _53280;
  wire _53282 = _13380 ^ _645;
  wire _53283 = _53282 ^ _15459;
  wire _53284 = uncoded_block[1312] ^ uncoded_block[1317];
  wire _53285 = _7802 ^ _53284;
  wire _53286 = _12287 ^ _40190;
  wire _53287 = _53285 ^ _53286;
  wire _53288 = _53283 ^ _53287;
  wire _53289 = _53281 ^ _53288;
  wire _53290 = uncoded_block[1335] ^ uncoded_block[1342];
  wire _53291 = _53290 ^ _17938;
  wire _53292 = _52024 ^ _53291;
  wire _53293 = _6588 ^ _25393;
  wire _53294 = _49916 ^ _53293;
  wire _53295 = _53292 ^ _53294;
  wire _53296 = _2283 ^ _4563;
  wire _53297 = _3054 ^ _29939;
  wire _53298 = _53296 ^ _53297;
  wire _53299 = _2293 ^ _694;
  wire _53300 = _52298 ^ _53299;
  wire _53301 = _53298 ^ _53300;
  wire _53302 = _53295 ^ _53301;
  wire _53303 = _53289 ^ _53302;
  wire _53304 = _53274 ^ _53303;
  wire _53305 = _13938 ^ _29090;
  wire _53306 = _53305 ^ _29946;
  wire _53307 = _3849 ^ _9021;
  wire _53308 = _24058 ^ _1530;
  wire _53309 = _53307 ^ _53308;
  wire _53310 = _53306 ^ _53309;
  wire _53311 = _3081 ^ _2314;
  wire _53312 = _24521 ^ _4590;
  wire _53313 = _53311 ^ _53312;
  wire _53314 = _5305 ^ _2322;
  wire _53315 = _53314 ^ _28356;
  wire _53316 = _53313 ^ _53315;
  wire _53317 = _53310 ^ _53316;
  wire _53318 = _11255 ^ _733;
  wire _53319 = _44350 ^ _53318;
  wire _53320 = _24982 ^ _46464;
  wire _53321 = _53319 ^ _53320;
  wire _53322 = _15512 ^ _22720;
  wire _53323 = _9055 ^ _9058;
  wire _53324 = _32142 ^ _53323;
  wire _53325 = _53322 ^ _53324;
  wire _53326 = _53321 ^ _53325;
  wire _53327 = _53317 ^ _53326;
  wire _53328 = _29122 ^ _23198;
  wire _53329 = _13979 ^ _1589;
  wire _53330 = _16499 ^ _13472;
  wire _53331 = _53329 ^ _53330;
  wire _53332 = _53328 ^ _53331;
  wire _53333 = _7889 ^ _24102;
  wire _53334 = _52067 ^ _53333;
  wire _53335 = uncoded_block[1573] ^ uncoded_block[1579];
  wire _53336 = _53335 ^ _18952;
  wire _53337 = _53336 ^ _15032;
  wire _53338 = _53334 ^ _53337;
  wire _53339 = _53332 ^ _53338;
  wire _53340 = _793 ^ _29551;
  wire _53341 = _35452 ^ _806;
  wire _53342 = _53340 ^ _53341;
  wire _53343 = _6046 ^ _1639;
  wire _53344 = _812 ^ _12949;
  wire _53345 = _53343 ^ _53344;
  wire _53346 = _6689 ^ _3169;
  wire _53347 = _53346 ^ _49479;
  wire _53348 = _53345 ^ _53347;
  wire _53349 = _53342 ^ _53348;
  wire _53350 = _53339 ^ _53349;
  wire _53351 = _53327 ^ _53350;
  wire _53352 = _53304 ^ _53351;
  wire _53353 = uncoded_block[1656] ^ uncoded_block[1663];
  wire _53354 = _53353 ^ _2422;
  wire _53355 = _22758 ^ _53354;
  wire _53356 = _6059 ^ _10766;
  wire _53357 = _3187 ^ _3189;
  wire _53358 = _53356 ^ _53357;
  wire _53359 = _53355 ^ _53358;
  wire _53360 = _47648 ^ _49992;
  wire _53361 = _2435 ^ _27671;
  wire _53362 = _53361 ^ _41018;
  wire _53363 = _53360 ^ _53362;
  wire _53364 = _53359 ^ _53363;
  wire _53365 = _53364 ^ uncoded_block[1721];
  wire _53366 = _53352 ^ _53365;
  wire _53367 = _53250 ^ _53366;
  wire _53368 = _5443 ^ _11363;
  wire _53369 = _14581 ^ _53368;
  wire _53370 = _52107 ^ _53369;
  wire _53371 = _52104 ^ _53370;
  wire _53372 = _9713 ^ _4026;
  wire _53373 = _12441 ^ _53372;
  wire _53374 = uncoded_block[108] ^ uncoded_block[114];
  wire _53375 = _6120 ^ _53374;
  wire _53376 = _28016 ^ _53375;
  wire _53377 = _53373 ^ _53376;
  wire _53378 = _48812 ^ _49174;
  wire _53379 = _53378 ^ _51817;
  wire _53380 = _53377 ^ _53379;
  wire _53381 = _53371 ^ _53380;
  wire _53382 = _4054 ^ _8591;
  wire _53383 = _52373 ^ _53382;
  wire _53384 = _48823 ^ _5477;
  wire _53385 = _53384 ^ _4063;
  wire _53386 = _53383 ^ _53385;
  wire _53387 = _51826 ^ _48081;
  wire _53388 = _51825 ^ _53387;
  wire _53389 = _53386 ^ _53388;
  wire _53390 = _4081 ^ _7422;
  wire _53391 = _53390 ^ _51831;
  wire _53392 = _53391 ^ _51833;
  wire _53393 = _53392 ^ _51840;
  wire _53394 = _53389 ^ _53393;
  wire _53395 = _53381 ^ _53394;
  wire _53396 = _6846 ^ _32274;
  wire _53397 = _53396 ^ _51845;
  wire _53398 = _51844 ^ _53397;
  wire _53399 = _48105 ^ _49218;
  wire _53400 = _3359 ^ _13089;
  wire _53401 = _51537 ^ _53400;
  wire _53402 = _53399 ^ _53401;
  wire _53403 = _53398 ^ _53402;
  wire _53404 = _52142 ^ _22415;
  wire _53405 = _53404 ^ _51856;
  wire _53406 = _16177 ^ _2629;
  wire _53407 = _52147 ^ _53406;
  wire _53408 = _51861 ^ _24248;
  wire _53409 = _53408 ^ _26937;
  wire _53410 = _53407 ^ _53409;
  wire _53411 = _53405 ^ _53410;
  wire _53412 = _53403 ^ _53411;
  wire _53413 = _50094 ^ _33566;
  wire _53414 = _4181 ^ _10362;
  wire _53415 = _53414 ^ _8687;
  wire _53416 = _53413 ^ _53415;
  wire _53417 = _9286 ^ _46246;
  wire _53418 = _24728 ^ _52162;
  wire _53419 = _53417 ^ _53418;
  wire _53420 = _53416 ^ _53419;
  wire _53421 = _9294 ^ _4908;
  wire _53422 = _23370 ^ _19638;
  wire _53423 = _53421 ^ _53422;
  wire _53424 = _1900 ^ _15230;
  wire _53425 = _40002 ^ _53424;
  wire _53426 = _53423 ^ _53425;
  wire _53427 = _6932 ^ _6293;
  wire _53428 = _53427 ^ _47398;
  wire _53429 = _31044 ^ _51224;
  wire _53430 = _53428 ^ _53429;
  wire _53431 = _53426 ^ _53430;
  wire _53432 = _53420 ^ _53431;
  wire _53433 = _53412 ^ _53432;
  wire _53434 = _53395 ^ _53433;
  wire _53435 = _24745 ^ _3472;
  wire _53436 = _53435 ^ _51578;
  wire _53437 = _48163 ^ _40409;
  wire _53438 = _53436 ^ _53437;
  wire _53439 = _51580 ^ _47041;
  wire _53440 = _19165 ^ _51585;
  wire _53441 = _53439 ^ _53440;
  wire _53442 = _53438 ^ _53441;
  wire _53443 = _46280 ^ _32755;
  wire _53444 = _53158 ^ _53443;
  wire _53445 = _52193 ^ _34035;
  wire _53446 = _51910 ^ _53445;
  wire _53447 = _53444 ^ _53446;
  wire _53448 = _53442 ^ _53447;
  wire _53449 = _52195 ^ _46295;
  wire _53450 = _22972 ^ _48934;
  wire _53451 = _53449 ^ _53450;
  wire _53452 = _52201 ^ _52204;
  wire _53453 = _43417 ^ _7617;
  wire _53454 = _49788 ^ _53453;
  wire _53455 = _53452 ^ _53454;
  wire _53456 = _53451 ^ _53455;
  wire _53457 = _5722 ^ _9392;
  wire _53458 = _52491 ^ _53457;
  wire _53459 = _385 ^ _34062;
  wire _53460 = _5041 ^ _51929;
  wire _53461 = _53459 ^ _53460;
  wire _53462 = _50903 ^ _52213;
  wire _53463 = _53461 ^ _53462;
  wire _53464 = _53458 ^ _53463;
  wire _53465 = _53456 ^ _53464;
  wire _53466 = _53448 ^ _53465;
  wire _53467 = _46322 ^ _52219;
  wire _53468 = _52220 ^ _52222;
  wire _53469 = _53467 ^ _53468;
  wire _53470 = _52223 ^ _17308;
  wire _53471 = _46336 ^ _8251;
  wire _53472 = _53470 ^ _53471;
  wire _53473 = _53469 ^ _53472;
  wire _53474 = _52515 ^ _7071;
  wire _53475 = _5092 ^ _8259;
  wire _53476 = _53475 ^ _51954;
  wire _53477 = _53474 ^ _53476;
  wire _53478 = _9976 ^ _49826;
  wire _53479 = _20717 ^ _51646;
  wire _53480 = _53478 ^ _53479;
  wire _53481 = _53477 ^ _53480;
  wire _53482 = _53473 ^ _53481;
  wire _53483 = _13271 ^ _8854;
  wire _53484 = _1318 ^ _28985;
  wire _53485 = _3660 ^ _53484;
  wire _53486 = _53483 ^ _53485;
  wire _53487 = _2107 ^ _40109;
  wire _53488 = _53487 ^ _52538;
  wire _53489 = _53488 ^ _52542;
  wire _53490 = _53486 ^ _53489;
  wire _53491 = _46363 ^ _51971;
  wire _53492 = _49005 ^ _23502;
  wire _53493 = _53491 ^ _53492;
  wire _53494 = _52549 ^ _50233;
  wire _53495 = _53494 ^ _52253;
  wire _53496 = _53493 ^ _53495;
  wire _53497 = _53490 ^ _53496;
  wire _53498 = _53482 ^ _53497;
  wire _53499 = _53466 ^ _53498;
  wire _53500 = _53434 ^ _53499;
  wire _53501 = _51676 ^ _43121;
  wire _53502 = _49380 ^ _53501;
  wire _53503 = _52255 ^ _53502;
  wire _53504 = _51997 ^ _48289;
  wire _53505 = _51993 ^ _53504;
  wire _53506 = _53503 ^ _53505;
  wire _53507 = _592 ^ _9508;
  wire _53508 = _53507 ^ _52271;
  wire _53509 = _53508 ^ _52275;
  wire _53510 = _31643 ^ _49399;
  wire _53511 = _51700 ^ _40171;
  wire _53512 = _53510 ^ _53511;
  wire _53513 = _53509 ^ _53512;
  wire _53514 = _53506 ^ _53513;
  wire _53515 = _52281 ^ _52285;
  wire _53516 = _18866 ^ _5916;
  wire _53517 = _53516 ^ _15459;
  wire _53518 = _53517 ^ _53287;
  wire _53519 = _53515 ^ _53518;
  wire _53520 = _19849 ^ _49063;
  wire _53521 = _52028 ^ _53293;
  wire _53522 = _53520 ^ _53521;
  wire _53523 = _2283 ^ _2289;
  wire _53524 = _53523 ^ _51726;
  wire _53525 = _53524 ^ _51729;
  wire _53526 = _53522 ^ _53525;
  wire _53527 = _53519 ^ _53526;
  wire _53528 = _53514 ^ _53527;
  wire _53529 = _5961 ^ _3853;
  wire _53530 = _3075 ^ _21783;
  wire _53531 = _53529 ^ _53530;
  wire _53532 = _51731 ^ _53531;
  wire _53533 = _37038 ^ _51042;
  wire _53534 = _51043 ^ _52050;
  wire _53535 = _53533 ^ _53534;
  wire _53536 = _53532 ^ _53535;
  wire _53537 = _23179 ^ _12342;
  wire _53538 = _42519 ^ _53537;
  wire _53539 = _741 ^ _39039;
  wire _53540 = _53538 ^ _53539;
  wire _53541 = _3894 ^ _4616;
  wire _53542 = _45099 ^ _53541;
  wire _53543 = _47228 ^ _11267;
  wire _53544 = _53543 ^ _24993;
  wire _53545 = _53542 ^ _53544;
  wire _53546 = _53540 ^ _53545;
  wire _53547 = _53536 ^ _53546;
  wire _53548 = _52063 ^ _52066;
  wire _53549 = _46487 ^ _3145;
  wire _53550 = _48374 ^ _53549;
  wire _53551 = _53334 ^ _53550;
  wire _53552 = _53548 ^ _53551;
  wire _53553 = _46494 ^ _52653;
  wire _53554 = _46492 ^ _53553;
  wire _53555 = _7912 ^ _46497;
  wire _53556 = _53555 ^ _33429;
  wire _53557 = _50359 ^ _49479;
  wire _53558 = _53556 ^ _53557;
  wire _53559 = _53554 ^ _53558;
  wire _53560 = _53552 ^ _53559;
  wire _53561 = _53547 ^ _53560;
  wire _53562 = _53528 ^ _53561;
  wire _53563 = _4679 ^ _51784;
  wire _53564 = _49985 ^ _51792;
  wire _53565 = _53563 ^ _53564;
  wire _53566 = _47648 ^ _51794;
  wire _53567 = _53566 ^ _46520;
  wire _53568 = _53565 ^ _53567;
  wire _53569 = _53562 ^ _53568;
  wire _53570 = _53500 ^ _53569;
  wire _53571 = _4710 ^ _21861;
  wire _53572 = _3995 ^ _33031;
  wire _53573 = _53571 ^ _53572;
  wire _53574 = uncoded_block[17] ^ uncoded_block[20];
  wire _53575 = _53574 ^ _4000;
  wire _53576 = _4001 ^ _21412;
  wire _53577 = _53575 ^ _53576;
  wire _53578 = _53573 ^ _53577;
  wire _53579 = _14569 ^ _880;
  wire _53580 = _53579 ^ _26387;
  wire _53581 = uncoded_block[53] ^ uncoded_block[57];
  wire _53582 = _13547 ^ _53581;
  wire _53583 = _20465 ^ _23698;
  wire _53584 = _53582 ^ _53583;
  wire _53585 = _53580 ^ _53584;
  wire _53586 = _53578 ^ _53585;
  wire _53587 = _34 ^ _7367;
  wire _53588 = _897 ^ _19019;
  wire _53589 = _53587 ^ _53588;
  wire _53590 = _19980 ^ _11909;
  wire _53591 = _53590 ^ _17585;
  wire _53592 = _53589 ^ _53591;
  wire _53593 = _915 ^ _13571;
  wire _53594 = _31383 ^ _53593;
  wire _53595 = _20961 ^ _1735;
  wire _53596 = _53595 ^ _17093;
  wire _53597 = _53594 ^ _53596;
  wire _53598 = _53592 ^ _53597;
  wire _53599 = _53586 ^ _53598;
  wire _53600 = uncoded_block[147] ^ uncoded_block[152];
  wire _53601 = _53600 ^ _5469;
  wire _53602 = _25081 ^ _53601;
  wire _53603 = _23281 ^ _21906;
  wire _53604 = uncoded_block[164] ^ uncoded_block[168];
  wire _53605 = _4053 ^ _53604;
  wire _53606 = _53603 ^ _53605;
  wire _53607 = _53602 ^ _53606;
  wire _53608 = _82 ^ _944;
  wire _53609 = _25978 ^ _53608;
  wire _53610 = _20983 ^ _15133;
  wire _53611 = _53609 ^ _53610;
  wire _53612 = _53607 ^ _53611;
  wire _53613 = _6801 ^ _6805;
  wire _53614 = _53613 ^ _21918;
  wire _53615 = _7415 ^ _17116;
  wire _53616 = _35136 ^ _105;
  wire _53617 = _53615 ^ _53616;
  wire _53618 = _53614 ^ _53617;
  wire _53619 = _967 ^ _35141;
  wire _53620 = _4082 ^ _53619;
  wire _53621 = _10292 ^ _21465;
  wire _53622 = _9212 ^ _4803;
  wire _53623 = _53621 ^ _53622;
  wire _53624 = _53620 ^ _53623;
  wire _53625 = _53618 ^ _53624;
  wire _53626 = _53612 ^ _53625;
  wire _53627 = _53599 ^ _53626;
  wire _53628 = uncoded_block[260] ^ uncoded_block[263];
  wire _53629 = _53628 ^ _977;
  wire _53630 = _30098 ^ _53629;
  wire _53631 = _21007 ^ _14124;
  wire _53632 = _1795 ^ _26447;
  wire _53633 = _53631 ^ _53632;
  wire _53634 = _53630 ^ _53633;
  wire _53635 = _6197 ^ _992;
  wire _53636 = _53635 ^ _10313;
  wire _53637 = _999 ^ _12515;
  wire _53638 = uncoded_block[308] ^ uncoded_block[313];
  wire _53639 = _53638 ^ _15168;
  wire _53640 = _53637 ^ _53639;
  wire _53641 = _53636 ^ _53640;
  wire _53642 = _53634 ^ _53641;
  wire _53643 = _6208 ^ _4123;
  wire _53644 = uncoded_block[332] ^ uncoded_block[338];
  wire _53645 = _1819 ^ _53644;
  wire _53646 = _53643 ^ _53645;
  wire _53647 = uncoded_block[339] ^ uncoded_block[343];
  wire _53648 = _53647 ^ _2599;
  wire _53649 = uncoded_block[354] ^ uncoded_block[357];
  wire _53650 = _53649 ^ _6864;
  wire _53651 = _53648 ^ _53650;
  wire _53652 = _53646 ^ _53651;
  wire _53653 = _168 ^ _1035;
  wire _53654 = _8079 ^ _4854;
  wire _53655 = _53653 ^ _53654;
  wire _53656 = _1841 ^ _4149;
  wire _53657 = uncoded_block[393] ^ uncoded_block[397];
  wire _53658 = _5554 ^ _53657;
  wire _53659 = _53656 ^ _53658;
  wire _53660 = _53655 ^ _53659;
  wire _53661 = _53652 ^ _53660;
  wire _53662 = _53642 ^ _53661;
  wire _53663 = _10911 ^ _6244;
  wire _53664 = _53663 ^ _22424;
  wire _53665 = _19612 ^ _13112;
  wire _53666 = _194 ^ _197;
  wire _53667 = _53665 ^ _53666;
  wire _53668 = _53664 ^ _53667;
  wire _53669 = _9820 ^ _21516;
  wire _53670 = _8097 ^ _53669;
  wire _53671 = _27757 ^ _1077;
  wire _53672 = _53670 ^ _53671;
  wire _53673 = _53668 ^ _53672;
  wire _53674 = _15715 ^ _7507;
  wire _53675 = _53674 ^ _1880;
  wire _53676 = _13132 ^ _5593;
  wire _53677 = _1090 ^ _3424;
  wire _53678 = _53676 ^ _53677;
  wire _53679 = _53675 ^ _53678;
  wire _53680 = uncoded_block[494] ^ uncoded_block[501];
  wire _53681 = uncoded_block[502] ^ uncoded_block[511];
  wire _53682 = _53680 ^ _53681;
  wire _53683 = uncoded_block[513] ^ uncoded_block[517];
  wire _53684 = _53683 ^ _4918;
  wire _53685 = _53682 ^ _53684;
  wire _53686 = _13684 ^ _6929;
  wire _53687 = _53686 ^ _24278;
  wire _53688 = _53685 ^ _53687;
  wire _53689 = _53679 ^ _53688;
  wire _53690 = _53673 ^ _53689;
  wire _53691 = _53662 ^ _53690;
  wire _53692 = _53627 ^ _53691;
  wire _53693 = _1908 ^ _1912;
  wire _53694 = _45658 ^ _53693;
  wire _53695 = _41151 ^ _14729;
  wire _53696 = _53694 ^ _53695;
  wire _53697 = _17221 ^ _6945;
  wire _53698 = _1132 ^ _38826;
  wire _53699 = _53697 ^ _53698;
  wire _53700 = _17721 ^ _28519;
  wire _53701 = _1942 ^ _12609;
  wire _53702 = _53700 ^ _53701;
  wire _53703 = _53699 ^ _53702;
  wire _53704 = _53696 ^ _53703;
  wire _53705 = _7570 ^ _22950;
  wire _53706 = _36010 ^ _53705;
  wire _53707 = _25203 ^ _5666;
  wire _53708 = _53706 ^ _53707;
  wire _53709 = _6338 ^ _301;
  wire _53710 = _302 ^ _10987;
  wire _53711 = _53709 ^ _53710;
  wire _53712 = _18705 ^ _7582;
  wire _53713 = _17742 ^ _2744;
  wire _53714 = _53712 ^ _53713;
  wire _53715 = _53711 ^ _53714;
  wire _53716 = _53708 ^ _53715;
  wire _53717 = _53704 ^ _53716;
  wire _53718 = _1968 ^ _321;
  wire _53719 = _34833 ^ _53718;
  wire _53720 = _6983 ^ _52822;
  wire _53721 = _53720 ^ _24778;
  wire _53722 = _53719 ^ _53721;
  wire _53723 = _2762 ^ _18726;
  wire _53724 = _26128 ^ _53723;
  wire _53725 = _12648 ^ _7001;
  wire _53726 = _8201 ^ _7605;
  wire _53727 = _53725 ^ _53726;
  wire _53728 = _53724 ^ _53727;
  wire _53729 = _53722 ^ _53728;
  wire _53730 = _5012 ^ _5704;
  wire _53731 = _38868 ^ _53730;
  wire _53732 = _5016 ^ _2003;
  wire _53733 = _53732 ^ _25230;
  wire _53734 = _53731 ^ _53733;
  wire _53735 = _3561 ^ _11019;
  wire _53736 = _53735 ^ _27016;
  wire _53737 = _19217 ^ _2794;
  wire _53738 = _6388 ^ _4314;
  wire _53739 = _53737 ^ _53738;
  wire _53740 = _53736 ^ _53739;
  wire _53741 = _53734 ^ _53740;
  wire _53742 = _53729 ^ _53741;
  wire _53743 = _53717 ^ _53742;
  wire _53744 = uncoded_block[808] ^ uncoded_block[812];
  wire _53745 = _34062 ^ _53744;
  wire _53746 = _39273 ^ _53745;
  wire _53747 = _4324 ^ _5046;
  wire _53748 = uncoded_block[821] ^ uncoded_block[827];
  wire _53749 = _53748 ^ _26160;
  wire _53750 = _53747 ^ _53749;
  wire _53751 = _53746 ^ _53750;
  wire _53752 = _38481 ^ _1257;
  wire _53753 = _4340 ^ _14814;
  wire _53754 = _53752 ^ _53753;
  wire _53755 = _2821 ^ _14300;
  wire _53756 = _53755 ^ _26166;
  wire _53757 = _53754 ^ _53756;
  wire _53758 = _53751 ^ _53757;
  wire _53759 = _8244 ^ _31131;
  wire _53760 = _32811 ^ _53759;
  wire _53761 = _25262 ^ _2844;
  wire _53762 = _45351 ^ _53761;
  wire _53763 = _53760 ^ _53762;
  wire _53764 = _18311 ^ _1284;
  wire _53765 = _53764 ^ _44213;
  wire _53766 = _439 ^ _9968;
  wire _53767 = _44215 ^ _53766;
  wire _53768 = _53765 ^ _53767;
  wire _53769 = _53763 ^ _53768;
  wire _53770 = _53758 ^ _53769;
  wire _53771 = uncoded_block[932] ^ uncoded_block[938];
  wire _53772 = _53771 ^ _4377;
  wire _53773 = _9433 ^ _5777;
  wire _53774 = _53772 ^ _53773;
  wire _53775 = _4381 ^ _4384;
  wire _53776 = _53775 ^ _28594;
  wire _53777 = _53774 ^ _53776;
  wire _53778 = _12179 ^ _7682;
  wire _53779 = _53778 ^ _38916;
  wire _53780 = _5114 ^ _8855;
  wire _53781 = _43844 ^ _29835;
  wire _53782 = _53780 ^ _53781;
  wire _53783 = _53779 ^ _53782;
  wire _53784 = _53777 ^ _53783;
  wire _53785 = _22584 ^ _2111;
  wire _53786 = _484 ^ _1327;
  wire _53787 = _53785 ^ _53786;
  wire _53788 = _13283 ^ _491;
  wire _53789 = uncoded_block[1021] ^ uncoded_block[1029];
  wire _53790 = _7703 ^ _53789;
  wire _53791 = _53788 ^ _53790;
  wire _53792 = _53787 ^ _53791;
  wire _53793 = _38937 ^ _12761;
  wire _53794 = _41265 ^ _53793;
  wire _53795 = uncoded_block[1057] ^ uncoded_block[1062];
  wire _53796 = _2914 ^ _53795;
  wire _53797 = _53796 ^ _14358;
  wire _53798 = _53794 ^ _53797;
  wire _53799 = _53792 ^ _53798;
  wire _53800 = _53784 ^ _53799;
  wire _53801 = _53770 ^ _53800;
  wire _53802 = _53743 ^ _53801;
  wire _53803 = _53692 ^ _53802;
  wire _53804 = _3691 ^ _8893;
  wire _53805 = _2925 ^ _7724;
  wire _53806 = _53804 ^ _53805;
  wire _53807 = _15401 ^ _1374;
  wire _53808 = _53807 ^ _30320;
  wire _53809 = _53806 ^ _53808;
  wire _53810 = uncoded_block[1101] ^ uncoded_block[1107];
  wire _53811 = _2935 ^ _53810;
  wire _53812 = _53811 ^ _2166;
  wire _53813 = _32044 ^ _47156;
  wire _53814 = _53812 ^ _53813;
  wire _53815 = _53809 ^ _53814;
  wire _53816 = _4460 ^ _15896;
  wire _53817 = _25329 ^ _53816;
  wire _53818 = _564 ^ _27528;
  wire _53819 = uncoded_block[1147] ^ uncoded_block[1150];
  wire _53820 = _574 ^ _53819;
  wire _53821 = _53818 ^ _53820;
  wire _53822 = _53817 ^ _53821;
  wire _53823 = _41690 ^ _22627;
  wire _53824 = _40149 ^ _53823;
  wire _53825 = _6511 ^ _5870;
  wire _53826 = _53825 ^ _3741;
  wire _53827 = _53824 ^ _53826;
  wire _53828 = _53822 ^ _53827;
  wire _53829 = _53815 ^ _53828;
  wire _53830 = _17397 ^ _9508;
  wire _53831 = _2201 ^ _3749;
  wire _53832 = _53830 ^ _53831;
  wire _53833 = _7758 ^ _2207;
  wire _53834 = _24911 ^ _53833;
  wire _53835 = _53832 ^ _53834;
  wire _53836 = _3762 ^ _30352;
  wire _53837 = _32071 ^ _53836;
  wire _53838 = _29045 ^ _612;
  wire _53839 = _5894 ^ _1440;
  wire _53840 = _53838 ^ _53839;
  wire _53841 = _53837 ^ _53840;
  wire _53842 = _53835 ^ _53841;
  wire _53843 = _33758 ^ _4511;
  wire _53844 = _44297 ^ _53843;
  wire _53845 = _15934 ^ _3003;
  wire _53846 = uncoded_block[1264] ^ uncoded_block[1268];
  wire _53847 = _53846 ^ _16419;
  wire _53848 = _53845 ^ _53847;
  wire _53849 = _53844 ^ _53848;
  wire _53850 = _21280 ^ _16924;
  wire _53851 = _11195 ^ _7193;
  wire _53852 = _53850 ^ _53851;
  wire _53853 = _645 ^ _10081;
  wire _53854 = _53853 ^ _34177;
  wire _53855 = _53852 ^ _53854;
  wire _53856 = _53849 ^ _53855;
  wire _53857 = _53842 ^ _53856;
  wire _53858 = _53829 ^ _53857;
  wire _53859 = _3026 ^ _21293;
  wire _53860 = _53859 ^ _31251;
  wire _53861 = uncoded_block[1330] ^ uncoded_block[1336];
  wire _53862 = _53861 ^ _1497;
  wire _53863 = _11215 ^ _1501;
  wire _53864 = _53862 ^ _53863;
  wire _53865 = _53860 ^ _53864;
  wire _53866 = _12857 ^ _48711;
  wire _53867 = _40940 ^ _53866;
  wire _53868 = _12861 ^ _11776;
  wire _53869 = _53868 ^ _10104;
  wire _53870 = _53867 ^ _53869;
  wire _53871 = _53865 ^ _53870;
  wire _53872 = _2290 ^ _29083;
  wire _53873 = _12867 ^ _20340;
  wire _53874 = _53872 ^ _53873;
  wire _53875 = _2296 ^ _9016;
  wire _53876 = _53875 ^ _50304;
  wire _53877 = _53874 ^ _53876;
  wire _53878 = _2308 ^ _5968;
  wire _53879 = _16464 ^ _53878;
  wire _53880 = _2318 ^ _2321;
  wire _53881 = _3858 ^ _53880;
  wire _53882 = _53879 ^ _53881;
  wire _53883 = _53877 ^ _53882;
  wire _53884 = _53871 ^ _53883;
  wire _53885 = _9033 ^ _719;
  wire _53886 = _720 ^ _2335;
  wire _53887 = _53885 ^ _53886;
  wire _53888 = _732 ^ _22707;
  wire _53889 = _42519 ^ _53888;
  wire _53890 = _53887 ^ _53889;
  wire _53891 = _1556 ^ _23181;
  wire _53892 = _17980 ^ _15996;
  wire _53893 = _53891 ^ _53892;
  wire _53894 = uncoded_block[1504] ^ uncoded_block[1508];
  wire _53895 = _747 ^ _53894;
  wire _53896 = _6632 ^ _53895;
  wire _53897 = _53893 ^ _53896;
  wire _53898 = _53890 ^ _53897;
  wire _53899 = _16001 ^ _9056;
  wire _53900 = _19897 ^ _3118;
  wire _53901 = uncoded_block[1529] ^ uncoded_block[1533];
  wire _53902 = _13459 ^ _53901;
  wire _53903 = _53900 ^ _53902;
  wire _53904 = _53899 ^ _53903;
  wire _53905 = uncoded_block[1541] ^ uncoded_block[1546];
  wire _53906 = _4632 ^ _53905;
  wire _53907 = _10157 ^ _22731;
  wire _53908 = _53906 ^ _53907;
  wire _53909 = _6016 ^ _44372;
  wire _53910 = _11284 ^ _7891;
  wire _53911 = _53909 ^ _53910;
  wire _53912 = _53908 ^ _53911;
  wire _53913 = _53904 ^ _53912;
  wire _53914 = _53898 ^ _53913;
  wire _53915 = _53884 ^ _53914;
  wire _53916 = _53858 ^ _53915;
  wire _53917 = uncoded_block[1580] ^ uncoded_block[1589];
  wire _53918 = _782 ^ _53917;
  wire _53919 = _9081 ^ _53918;
  wire _53920 = _1620 ^ _3151;
  wire _53921 = _40991 ^ _53920;
  wire _53922 = _53919 ^ _53921;
  wire _53923 = _1625 ^ _6040;
  wire _53924 = _801 ^ _6042;
  wire _53925 = _53923 ^ _53924;
  wire _53926 = _10181 ^ _7298;
  wire _53927 = _53926 ^ _20899;
  wire _53928 = _53925 ^ _53927;
  wire _53929 = _53922 ^ _53928;
  wire _53930 = _23658 ^ _9659;
  wire _53931 = _15555 ^ _4673;
  wire _53932 = _53930 ^ _53931;
  wire _53933 = _2412 ^ _10757;
  wire _53934 = _8515 ^ _822;
  wire _53935 = _53933 ^ _53934;
  wire _53936 = _53932 ^ _53935;
  wire _53937 = _12960 ^ _7319;
  wire _53938 = _53937 ^ _27659;
  wire _53939 = _10767 ^ _53037;
  wire _53940 = _53938 ^ _53939;
  wire _53941 = _53936 ^ _53940;
  wire _53942 = _53929 ^ _53941;
  wire _53943 = uncoded_block[1705] ^ uncoded_block[1710];
  wire _53944 = _20920 ^ _53943;
  wire _53945 = _9671 ^ _53944;
  wire _53946 = _29581 ^ _19485;
  wire _53947 = _53945 ^ _53946;
  wire _53948 = _53947 ^ _12977;
  wire _53949 = _53942 ^ _53948;
  wire _53950 = _53916 ^ _53949;
  wire _53951 = _53803 ^ _53950;
  wire _53952 = _48790 ^ _53051;
  wire _53953 = _10791 ^ _11344;
  wire _53954 = _53953 ^ _19969;
  wire _53955 = _53952 ^ _53954;
  wire _53956 = uncoded_block[68] ^ uncoded_block[75];
  wire _53957 = _53956 ^ _901;
  wire _53958 = _49636 ^ _53957;
  wire _53959 = _52107 ^ _53958;
  wire _53960 = _53955 ^ _53959;
  wire _53961 = _35502 ^ _30933;
  wire _53962 = _53961 ^ _52363;
  wire _53963 = _53374 ^ _48432;
  wire _53964 = _53963 ^ _13018;
  wire _53965 = _4760 ^ _11918;
  wire _53966 = _46174 ^ _53965;
  wire _53967 = _53964 ^ _53966;
  wire _53968 = _53962 ^ _53967;
  wire _53969 = _53960 ^ _53968;
  wire _53970 = _33909 ^ _52371;
  wire _53971 = _53970 ^ _52373;
  wire _53972 = _52375 ^ _51505;
  wire _53973 = _53971 ^ _53972;
  wire _53974 = _51507 ^ _947;
  wire _53975 = _53974 ^ _12477;
  wire _53976 = _4070 ^ _3296;
  wire _53977 = _51512 ^ _53976;
  wire _53978 = _53975 ^ _53977;
  wire _53979 = _53973 ^ _53978;
  wire _53980 = _28799 ^ _51516;
  wire _53981 = _20510 ^ _37956;
  wire _53982 = _53980 ^ _53981;
  wire _53983 = _39154 ^ _9761;
  wire _53984 = _1786 ^ _37959;
  wire _53985 = _53983 ^ _53984;
  wire _53986 = _16636 ^ _7445;
  wire _53987 = _988 ^ _49687;
  wire _53988 = _53986 ^ _53987;
  wire _53989 = _53985 ^ _53988;
  wire _53990 = _53982 ^ _53989;
  wire _53991 = _53979 ^ _53990;
  wire _53992 = _53969 ^ _53991;
  wire _53993 = _52129 ^ _10312;
  wire _53994 = _53993 ^ _51529;
  wire _53995 = _51530 ^ _52405;
  wire _53996 = _53994 ^ _53995;
  wire _53997 = _51845 ^ _33536;
  wire _53998 = _50070 ^ _46219;
  wire _53999 = _53997 ^ _53998;
  wire _54000 = _53996 ^ _53999;
  wire _54001 = _30123 ^ _3361;
  wire _54002 = _50076 ^ _1835;
  wire _54003 = _54001 ^ _54002;
  wire _54004 = _9796 ^ _51854;
  wire _54005 = _54003 ^ _54004;
  wire _54006 = _13646 ^ _16177;
  wire _54007 = _49710 ^ _54006;
  wire _54008 = _2629 ^ _1054;
  wire _54009 = _54008 ^ _52151;
  wire _54010 = _54007 ^ _54009;
  wire _54011 = _54005 ^ _54010;
  wire _54012 = _54000 ^ _54011;
  wire _54013 = uncoded_block[431] ^ uncoded_block[441];
  wire _54014 = _54013 ^ _21974;
  wire _54015 = _54014 ^ _46239;
  wire _54016 = _9280 ^ _13662;
  wire _54017 = _54016 ^ _9284;
  wire _54018 = _54015 ^ _54017;
  wire _54019 = _24721 ^ _51559;
  wire _54020 = _54019 ^ _51561;
  wire _54021 = _27769 ^ _4905;
  wire _54022 = _10375 ^ _3437;
  wire _54023 = _54021 ^ _54022;
  wire _54024 = _54020 ^ _54023;
  wire _54025 = _54018 ^ _54024;
  wire _54026 = _13148 ^ _4208;
  wire _54027 = _54026 ^ _8709;
  wire _54028 = _1905 ^ _3451;
  wire _54029 = _30173 ^ _54028;
  wire _54030 = _54027 ^ _54029;
  wire _54031 = _244 ^ _5628;
  wire _54032 = _45658 ^ _54031;
  wire _54033 = _6940 ^ _24745;
  wire _54034 = _31044 ^ _54033;
  wire _54035 = _54032 ^ _54034;
  wire _54036 = _54030 ^ _54035;
  wire _54037 = _54025 ^ _54036;
  wire _54038 = _54012 ^ _54037;
  wire _54039 = _53992 ^ _54038;
  wire _54040 = _33602 ^ _51233;
  wire _54041 = _46269 ^ _54040;
  wire _54042 = _18227 ^ _279;
  wire _54043 = _2719 ^ _1156;
  wire _54044 = _46274 ^ _54043;
  wire _54045 = _54042 ^ _54044;
  wire _54046 = _54041 ^ _54045;
  wire _54047 = _6330 ^ _4249;
  wire _54048 = _54047 ^ _12077;
  wire _54049 = _46280 ^ _46282;
  wire _54050 = _54048 ^ _54049;
  wire _54051 = _46283 ^ _17251;
  wire _54052 = _1971 ^ _52469;
  wire _54053 = _54052 ^ _51600;
  wire _54054 = _54051 ^ _54053;
  wire _54055 = _54050 ^ _54054;
  wire _54056 = _54046 ^ _54055;
  wire _54057 = _51257 ^ _53172;
  wire _54058 = _53174 ^ _12104;
  wire _54059 = _54057 ^ _54058;
  wire _54060 = _43417 ^ _30659;
  wire _54061 = _49788 ^ _54060;
  wire _54062 = _53452 ^ _54061;
  wire _54063 = _54059 ^ _54062;
  wire _54064 = _3568 ^ _51274;
  wire _54065 = _7621 ^ _54064;
  wire _54066 = _31551 ^ _34062;
  wire _54067 = _376 ^ _54066;
  wire _54068 = _54065 ^ _54067;
  wire _54069 = _53460 ^ _50903;
  wire _54070 = uncoded_block[823] ^ uncoded_block[835];
  wire _54071 = _54070 ^ _12138;
  wire _54072 = _54071 ^ _47095;
  wire _54073 = _54069 ^ _54072;
  wire _54074 = _54068 ^ _54073;
  wire _54075 = _54063 ^ _54074;
  wire _54076 = _54056 ^ _54075;
  wire _54077 = _52506 ^ _2828;
  wire _54078 = _54077 ^ _51943;
  wire _54079 = _51632 ^ _54078;
  wire _54080 = _4351 ^ _14821;
  wire _54081 = _54080 ^ _50917;
  wire _54082 = _5085 ^ _1278;
  wire _54083 = _54082 ^ _52515;
  wire _54084 = _54081 ^ _54083;
  wire _54085 = _54079 ^ _54084;
  wire _54086 = _37717 ^ _53204;
  wire _54087 = _3631 ^ _33684;
  wire _54088 = _54087 ^ _49341;
  wire _54089 = _54086 ^ _54088;
  wire _54090 = _52234 ^ _4383;
  wire _54091 = _12726 ^ _1308;
  wire _54092 = _54091 ^ _51646;
  wire _54093 = _54090 ^ _54092;
  wire _54094 = _54089 ^ _54093;
  wire _54095 = _54085 ^ _54094;
  wire _54096 = _13271 ^ _52532;
  wire _54097 = _23939 ^ _28985;
  wire _54098 = _51654 ^ _54097;
  wire _54099 = _54096 ^ _54098;
  wire _54100 = _23945 ^ _2114;
  wire _54101 = _54100 ^ _48251;
  wire _54102 = _54101 ^ _51968;
  wire _54103 = _54099 ^ _54102;
  wire _54104 = _30306 ^ _511;
  wire _54105 = _2910 ^ _42039;
  wire _54106 = _54104 ^ _54105;
  wire _54107 = _54106 ^ _52250;
  wire _54108 = _49010 ^ _18822;
  wire _54109 = _52251 ^ _54108;
  wire _54110 = _54107 ^ _54109;
  wire _54111 = _54103 ^ _54110;
  wire _54112 = _54095 ^ _54111;
  wire _54113 = _54076 ^ _54112;
  wire _54114 = _54039 ^ _54113;
  wire _54115 = _1380 ^ _8910;
  wire _54116 = _34943 ^ _51674;
  wire _54117 = _54115 ^ _54116;
  wire _54118 = _45019 ^ _30329;
  wire _54119 = _49380 ^ _54118;
  wire _54120 = _54117 ^ _54119;
  wire _54121 = _52264 ^ _46392;
  wire _54122 = _17392 ^ _5872;
  wire _54123 = _51997 ^ _54122;
  wire _54124 = _54121 ^ _54123;
  wire _54125 = _54120 ^ _54124;
  wire _54126 = _29891 ^ _49883;
  wire _54127 = _52001 ^ _54126;
  wire _54128 = _40166 ^ _31231;
  wire _54129 = _49399 ^ _54128;
  wire _54130 = _51698 ^ _54129;
  wire _54131 = _54127 ^ _54130;
  wire _54132 = _54125 ^ _54131;
  wire _54133 = _48303 ^ _30359;
  wire _54134 = _34564 ^ _51707;
  wire _54135 = _54133 ^ _54134;
  wire _54136 = _51712 ^ _53516;
  wire _54137 = _15459 ^ _14941;
  wire _54138 = _54136 ^ _54137;
  wire _54139 = _54135 ^ _54138;
  wire _54140 = _9552 ^ _12287;
  wire _54141 = _40190 ^ _1494;
  wire _54142 = _54140 ^ _54141;
  wire _54143 = _14440 ^ _17938;
  wire _54144 = _37817 ^ _54143;
  wire _54145 = _54142 ^ _54144;
  wire _54146 = _21303 ^ _5940;
  wire _54147 = _54146 ^ _53293;
  wire _54148 = _2283 ^ _6594;
  wire _54149 = _54148 ^ _52605;
  wire _54150 = _54147 ^ _54149;
  wire _54151 = _54145 ^ _54150;
  wire _54152 = _54139 ^ _54151;
  wire _54153 = _54132 ^ _54152;
  wire _54154 = _6596 ^ _1513;
  wire _54155 = _54154 ^ _5953;
  wire _54156 = _13938 ^ _4572;
  wire _54157 = _54156 ^ _29501;
  wire _54158 = _54155 ^ _54157;
  wire _54159 = _701 ^ _5961;
  wire _54160 = _33374 ^ _16463;
  wire _54161 = _54159 ^ _54160;
  wire _54162 = _21783 ^ _3857;
  wire _54163 = _52614 ^ _54162;
  wire _54164 = _54161 ^ _54163;
  wire _54165 = _54158 ^ _54164;
  wire _54166 = _18913 ^ _4592;
  wire _54167 = _717 ^ _42512;
  wire _54168 = _2329 ^ _726;
  wire _54169 = _54167 ^ _54168;
  wire _54170 = _54166 ^ _54169;
  wire _54171 = _7247 ^ _23179;
  wire _54172 = _47599 ^ _54171;
  wire _54173 = uncoded_block[1489] ^ uncoded_block[1495];
  wire _54174 = _54173 ^ _743;
  wire _54175 = _51748 ^ _54174;
  wire _54176 = _54172 ^ _54175;
  wire _54177 = _54170 ^ _54176;
  wire _54178 = _54165 ^ _54177;
  wire _54179 = _4617 ^ _9055;
  wire _54180 = _6643 ^ _15004;
  wire _54181 = _54179 ^ _54180;
  wire _54182 = _53542 ^ _54181;
  wire _54183 = _29122 ^ _5345;
  wire _54184 = _46475 ^ _13988;
  wire _54185 = _54183 ^ _54184;
  wire _54186 = _54182 ^ _54185;
  wire _54187 = _13472 ^ _5358;
  wire _54188 = _54187 ^ _49958;
  wire _54189 = _2376 ^ _16020;
  wire _54190 = _54189 ^ _46486;
  wire _54191 = _54188 ^ _54190;
  wire _54192 = _53549 ^ _46490;
  wire _54193 = _5373 ^ _9088;
  wire _54194 = _54193 ^ _52077;
  wire _54195 = _54192 ^ _54194;
  wire _54196 = _54191 ^ _54195;
  wire _54197 = _54186 ^ _54196;
  wire _54198 = _54178 ^ _54197;
  wire _54199 = _54153 ^ _54198;
  wire _54200 = uncoded_block[1622] ^ uncoded_block[1630];
  wire _54201 = _54200 ^ _5388;
  wire _54202 = _29145 ^ _54201;
  wire _54203 = _18965 ^ _7309;
  wire _54204 = _4673 ^ _6691;
  wire _54205 = _54203 ^ _54204;
  wire _54206 = _54202 ^ _54205;
  wire _54207 = _19463 ^ _10762;
  wire _54208 = _33012 ^ _19475;
  wire _54209 = _52089 ^ _54208;
  wire _54210 = _54207 ^ _54209;
  wire _54211 = _54206 ^ _54210;
  wire _54212 = _837 ^ _9115;
  wire _54213 = _54212 ^ _52094;
  wire _54214 = _35477 ^ _10214;
  wire _54215 = uncoded_block[1710] ^ uncoded_block[1714];
  wire _54216 = uncoded_block[1715] ^ uncoded_block[1718];
  wire _54217 = _54215 ^ _54216;
  wire _54218 = _54214 ^ _54217;
  wire _54219 = _54213 ^ _54218;
  wire _54220 = _54219 ^ _861;
  wire _54221 = _54211 ^ _54220;
  wire _54222 = _54199 ^ _54221;
  wire _54223 = _54114 ^ _54222;
  wire _54224 = _4712 ^ _2454;
  wire _54225 = _3998 ^ _13537;
  wire _54226 = _54224 ^ _54225;
  wire _54227 = _24606 ^ _19501;
  wire _54228 = _3221 ^ _54227;
  wire _54229 = _54226 ^ _54228;
  wire _54230 = uncoded_block[38] ^ uncoded_block[50];
  wire _54231 = _54230 ^ _886;
  wire _54232 = uncoded_block[57] ^ uncoded_block[64];
  wire _54233 = _10238 ^ _54232;
  wire _54234 = _54231 ^ _54233;
  wire _54235 = _4728 ^ _39;
  wire _54236 = _10246 ^ _18077;
  wire _54237 = _54235 ^ _54236;
  wire _54238 = _54234 ^ _54237;
  wire _54239 = _54229 ^ _54238;
  wire _54240 = _4745 ^ _19025;
  wire _54241 = _17081 ^ _54240;
  wire _54242 = _50 ^ _15103;
  wire _54243 = _54242 ^ _28445;
  wire _54244 = _54241 ^ _54243;
  wire _54245 = _6128 ^ _20961;
  wire _54246 = _54245 ^ _36318;
  wire _54247 = _11918 ^ _11381;
  wire _54248 = _47691 ^ _54247;
  wire _54249 = _54246 ^ _54248;
  wire _54250 = _54244 ^ _54249;
  wire _54251 = _54239 ^ _54250;
  wire _54252 = _42602 ^ _21905;
  wire _54253 = _54252 ^ _25532;
  wire _54254 = _4054 ^ _7399;
  wire _54255 = _10841 ^ _85;
  wire _54256 = _54254 ^ _54255;
  wire _54257 = _54253 ^ _54256;
  wire _54258 = _8009 ^ _15631;
  wire _54259 = _54258 ^ _21453;
  wire _54260 = _94 ^ _8018;
  wire _54261 = _28796 ^ _102;
  wire _54262 = _54260 ^ _54261;
  wire _54263 = _54259 ^ _54262;
  wire _54264 = _54257 ^ _54263;
  wire _54265 = _4791 ^ _18123;
  wire _54266 = _106 ^ _54265;
  wire _54267 = _9211 ^ _1781;
  wire _54268 = _30090 ^ _54267;
  wire _54269 = _54266 ^ _54268;
  wire _54270 = _11954 ^ _9761;
  wire _54271 = _54270 ^ _6828;
  wire _54272 = uncoded_block[264] ^ uncoded_block[271];
  wire _54273 = _54272 ^ _5512;
  wire _54274 = _10303 ^ _7446;
  wire _54275 = _54273 ^ _54274;
  wire _54276 = _54271 ^ _54275;
  wire _54277 = _54269 ^ _54276;
  wire _54278 = _54264 ^ _54277;
  wire _54279 = _54251 ^ _54278;
  wire _54280 = _31842 ^ _4820;
  wire _54281 = _21016 ^ _6845;
  wire _54282 = _54280 ^ _54281;
  wire _54283 = _6846 ^ _16149;
  wire _54284 = _1008 ^ _3347;
  wire _54285 = _54283 ^ _54284;
  wire _54286 = _54282 ^ _54285;
  wire _54287 = _6853 ^ _5536;
  wire _54288 = _54287 ^ _6215;
  wire _54289 = _3355 ^ _1023;
  wire _54290 = _11454 ^ _3361;
  wire _54291 = _54289 ^ _54290;
  wire _54292 = _54288 ^ _54291;
  wire _54293 = _54286 ^ _54292;
  wire _54294 = uncoded_block[363] ^ uncoded_block[369];
  wire _54295 = _6864 ^ _54294;
  wire _54296 = uncoded_block[370] ^ uncoded_block[377];
  wire _54297 = _54296 ^ _10899;
  wire _54298 = _54295 ^ _54297;
  wire _54299 = _9801 ^ _6240;
  wire _54300 = _54298 ^ _54299;
  wire _54301 = _1849 ^ _4865;
  wire _54302 = _26924 ^ _54301;
  wire _54303 = _49231 ^ _8091;
  wire _54304 = uncoded_block[417] ^ uncoded_block[423];
  wire _54305 = _2630 ^ _54304;
  wire _54306 = _54303 ^ _54305;
  wire _54307 = _54302 ^ _54306;
  wire _54308 = _54300 ^ _54307;
  wire _54309 = _54293 ^ _54308;
  wire _54310 = _1857 ^ _9820;
  wire _54311 = _51863 ^ _54310;
  wire _54312 = _5577 ^ _21974;
  wire _54313 = _54312 ^ _35581;
  wire _54314 = _54311 ^ _54313;
  wire _54315 = _2652 ^ _26942;
  wire _54316 = _21059 ^ _1082;
  wire _54317 = _54316 ^ _27356;
  wire _54318 = _54315 ^ _54317;
  wire _54319 = _54314 ^ _54318;
  wire _54320 = _5598 ^ _7515;
  wire _54321 = _7516 ^ _27769;
  wire _54322 = _54320 ^ _54321;
  wire _54323 = uncoded_block[500] ^ uncoded_block[506];
  wire _54324 = _4905 ^ _54323;
  wire _54325 = _9294 ^ _8705;
  wire _54326 = _54324 ^ _54325;
  wire _54327 = _54322 ^ _54326;
  wire _54328 = _4918 ^ _1898;
  wire _54329 = _4921 ^ _1111;
  wire _54330 = _54328 ^ _54329;
  wire _54331 = _6292 ^ _24279;
  wire _54332 = _54331 ^ _38818;
  wire _54333 = _54330 ^ _54332;
  wire _54334 = _54327 ^ _54333;
  wire _54335 = _54319 ^ _54334;
  wire _54336 = _54309 ^ _54335;
  wire _54337 = _54279 ^ _54336;
  wire _54338 = _1123 ^ _1125;
  wire _54339 = _3460 ^ _54338;
  wire _54340 = _5635 ^ _20615;
  wire _54341 = _54340 ^ _16723;
  wire _54342 = _54339 ^ _54341;
  wire _54343 = _16225 ^ _42668;
  wire _54344 = _4953 ^ _5646;
  wire _54345 = _22466 ^ _54344;
  wire _54346 = _54343 ^ _54345;
  wire _54347 = _54342 ^ _54346;
  wire _54348 = _9870 ^ _2713;
  wire _54349 = _8744 ^ _22024;
  wire _54350 = _54348 ^ _54349;
  wire _54351 = _8159 ^ _289;
  wire _54352 = _27395 ^ _2727;
  wire _54353 = _54351 ^ _54352;
  wire _54354 = _54350 ^ _54353;
  wire _54355 = _4256 ^ _15766;
  wire _54356 = _54355 ^ _40796;
  wire _54357 = _1173 ^ _28158;
  wire _54358 = _15769 ^ _54357;
  wire _54359 = _54356 ^ _54358;
  wire _54360 = _54354 ^ _54359;
  wire _54361 = _54347 ^ _54360;
  wire _54362 = uncoded_block[674] ^ uncoded_block[682];
  wire _54363 = _54362 ^ _15281;
  wire _54364 = _1974 ^ _4272;
  wire _54365 = _54363 ^ _54364;
  wire _54366 = _8186 ^ _14766;
  wire _54367 = _6361 ^ _23863;
  wire _54368 = _54366 ^ _54367;
  wire _54369 = _54365 ^ _54368;
  wire _54370 = _5690 ^ _3544;
  wire _54371 = _44939 ^ _54370;
  wire _54372 = _13205 ^ _47436;
  wire _54373 = _54371 ^ _54372;
  wire _54374 = _54369 ^ _54373;
  wire _54375 = _5010 ^ _5702;
  wire _54376 = _1999 ^ _357;
  wire _54377 = _54375 ^ _54376;
  wire _54378 = _13213 ^ _2783;
  wire _54379 = uncoded_block[772] ^ uncoded_block[782];
  wire _54380 = _7617 ^ _54379;
  wire _54381 = _54378 ^ _54380;
  wire _54382 = _54377 ^ _54381;
  wire _54383 = _4309 ^ _8215;
  wire _54384 = _10475 ^ _6391;
  wire _54385 = _54383 ^ _54384;
  wire _54386 = _43803 ^ _20178;
  wire _54387 = _54385 ^ _54386;
  wire _54388 = _54382 ^ _54387;
  wire _54389 = _54374 ^ _54388;
  wire _54390 = _54361 ^ _54389;
  wire _54391 = _12131 ^ _1246;
  wire _54392 = _51930 ^ _54391;
  wire _54393 = uncoded_block[827] ^ uncoded_block[835];
  wire _54394 = _54393 ^ _2814;
  wire _54395 = _5737 ^ _1257;
  wire _54396 = _54394 ^ _54395;
  wire _54397 = _54392 ^ _54396;
  wire _54398 = uncoded_block[848] ^ uncoded_block[853];
  wire _54399 = _54398 ^ _3600;
  wire _54400 = _6410 ^ _49330;
  wire _54401 = _54399 ^ _54400;
  wire _54402 = uncoded_block[877] ^ uncoded_block[884];
  wire _54403 = _30260 ^ _54402;
  wire _54404 = _11059 ^ _3614;
  wire _54405 = _54403 ^ _54404;
  wire _54406 = _54401 ^ _54405;
  wire _54407 = _54397 ^ _54406;
  wire _54408 = uncoded_block[902] ^ uncoded_block[909];
  wire _54409 = _54408 ^ _19252;
  wire _54410 = _13802 ^ _54409;
  wire _54411 = _1287 ^ _23917;
  wire _54412 = _29379 ^ _7075;
  wire _54413 = _54411 ^ _54412;
  wire _54414 = _54410 ^ _54413;
  wire _54415 = _25736 ^ _9971;
  wire _54416 = _54415 ^ _52523;
  wire _54417 = _5777 ^ _8842;
  wire _54418 = _461 ^ _45753;
  wire _54419 = _54417 ^ _54418;
  wire _54420 = _54416 ^ _54419;
  wire _54421 = _54414 ^ _54420;
  wire _54422 = _54407 ^ _54421;
  wire _54423 = _5785 ^ _1314;
  wire _54424 = _4390 ^ _8853;
  wire _54425 = _54423 ^ _54424;
  wire _54426 = uncoded_block[989] ^ uncoded_block[993];
  wire _54427 = _54426 ^ _479;
  wire _54428 = _35310 ^ _54427;
  wire _54429 = _54425 ^ _54428;
  wire _54430 = _32431 ^ _484;
  wire _54431 = _54430 ^ _13284;
  wire _54432 = _47133 ^ _5806;
  wire _54433 = _42033 ^ _54432;
  wire _54434 = _54431 ^ _54433;
  wire _54435 = _54429 ^ _54434;
  wire _54436 = _9464 ^ _1359;
  wire _54437 = _8883 ^ _54436;
  wire _54438 = _7117 ^ _2140;
  wire _54439 = _54438 ^ _24880;
  wire _54440 = _54437 ^ _54439;
  wire _54441 = _9479 ^ _51976;
  wire _54442 = _15401 ^ _12774;
  wire _54443 = _5840 ^ _11139;
  wire _54444 = _54442 ^ _54443;
  wire _54445 = _54441 ^ _54444;
  wire _54446 = _54440 ^ _54445;
  wire _54447 = _54435 ^ _54446;
  wire _54448 = _54422 ^ _54447;
  wire _54449 = _54390 ^ _54448;
  wire _54450 = _54337 ^ _54449;
  wire _54451 = _12224 ^ _9484;
  wire _54452 = _4450 ^ _46066;
  wire _54453 = _54451 ^ _54452;
  wire _54454 = _2942 ^ _5854;
  wire _54455 = _6499 ^ _6501;
  wire _54456 = _54454 ^ _54455;
  wire _54457 = _54453 ^ _54456;
  wire _54458 = _41288 ^ _5184;
  wire _54459 = _2185 ^ _8354;
  wire _54460 = _54458 ^ _54459;
  wire _54461 = _30756 ^ _1408;
  wire _54462 = _5191 ^ _54461;
  wire _54463 = _54460 ^ _54462;
  wire _54464 = _54457 ^ _54463;
  wire _54465 = _32064 ^ _3742;
  wire _54466 = _43510 ^ _11721;
  wire _54467 = _54465 ^ _54466;
  wire _54468 = _2217 ^ _26694;
  wire _54469 = _4492 ^ _54468;
  wire _54470 = _54467 ^ _54469;
  wire _54471 = uncoded_block[1213] ^ uncoded_block[1219];
  wire _54472 = _54471 ^ _608;
  wire _54473 = _11177 ^ _13357;
  wire _54474 = _54472 ^ _54473;
  wire _54475 = _31228 ^ _15927;
  wire _54476 = _5221 ^ _31231;
  wire _54477 = _54475 ^ _54476;
  wire _54478 = _54474 ^ _54477;
  wire _54479 = _54470 ^ _54478;
  wire _54480 = _54464 ^ _54479;
  wire _54481 = _7780 ^ _2238;
  wire _54482 = _6550 ^ _46419;
  wire _54483 = _54481 ^ _54482;
  wire _54484 = _54133 ^ _54483;
  wire _54485 = _49897 ^ _3793;
  wire _54486 = _54485 ^ _53279;
  wire _54487 = _35379 ^ _9548;
  wire _54488 = _54486 ^ _54487;
  wire _54489 = _54484 ^ _54488;
  wire _54490 = _17435 ^ _5919;
  wire _54491 = _49054 ^ _54490;
  wire _54492 = _1487 ^ _34581;
  wire _54493 = _660 ^ _9563;
  wire _54494 = _54492 ^ _54493;
  wire _54495 = _54491 ^ _54494;
  wire _54496 = _4553 ^ _11215;
  wire _54497 = uncoded_block[1346] ^ uncoded_block[1353];
  wire _54498 = uncoded_block[1355] ^ uncoded_block[1363];
  wire _54499 = _54497 ^ _54498;
  wire _54500 = _54496 ^ _54499;
  wire _54501 = uncoded_block[1381] ^ uncoded_block[1385];
  wire _54502 = _10669 ^ _54501;
  wire _54503 = _8422 ^ _54502;
  wire _54504 = _54500 ^ _54503;
  wire _54505 = _54495 ^ _54504;
  wire _54506 = _54489 ^ _54505;
  wire _54507 = _54480 ^ _54506;
  wire _54508 = _1513 ^ _23157;
  wire _54509 = _54508 ^ _28689;
  wire _54510 = uncoded_block[1403] ^ uncoded_block[1410];
  wire _54511 = uncoded_block[1412] ^ uncoded_block[1417];
  wire _54512 = _54510 ^ _54511;
  wire _54513 = _5964 ^ _1527;
  wire _54514 = _54512 ^ _54513;
  wire _54515 = _54509 ^ _54514;
  wire _54516 = _3075 ^ _5299;
  wire _54517 = _54516 ^ _30832;
  wire _54518 = uncoded_block[1441] ^ uncoded_block[1446];
  wire _54519 = _54518 ^ _11246;
  wire _54520 = _13437 ^ _726;
  wire _54521 = _54519 ^ _54520;
  wire _54522 = _54517 ^ _54521;
  wire _54523 = _54515 ^ _54522;
  wire _54524 = _8455 ^ _5314;
  wire _54525 = _1551 ^ _42807;
  wire _54526 = _54524 ^ _54525;
  wire _54527 = _740 ^ _5329;
  wire _54528 = _16979 ^ _54527;
  wire _54529 = _54526 ^ _54528;
  wire _54530 = _2352 ^ _1571;
  wire _54531 = _11813 ^ _5333;
  wire _54532 = _54530 ^ _54531;
  wire _54533 = _1575 ^ _751;
  wire _54534 = _54533 ^ _51757;
  wire _54535 = _54532 ^ _54534;
  wire _54536 = _54529 ^ _54535;
  wire _54537 = _54523 ^ _54536;
  wire _54538 = _9059 ^ _9626;
  wire _54539 = _54538 ^ _18488;
  wire _54540 = _5347 ^ _15009;
  wire _54541 = _43967 ^ _7277;
  wire _54542 = _54540 ^ _54541;
  wire _54543 = _54539 ^ _54542;
  wire _54544 = _769 ^ _3914;
  wire _54545 = _54544 ^ _45887;
  wire _54546 = _14506 ^ _3924;
  wire _54547 = _25008 ^ _792;
  wire _54548 = _54546 ^ _54547;
  wire _54549 = _54545 ^ _54548;
  wire _54550 = _54543 ^ _54549;
  wire _54551 = uncoded_block[1605] ^ uncoded_block[1613];
  wire _54552 = _54551 ^ _29997;
  wire _54553 = _12376 ^ _3941;
  wire _54554 = _54552 ^ _54553;
  wire _54555 = _5388 ^ _14009;
  wire _54556 = _32173 ^ _54555;
  wire _54557 = _54554 ^ _54556;
  wire _54558 = _3169 ^ _7312;
  wire _54559 = _12387 ^ _10760;
  wire _54560 = _54558 ^ _54559;
  wire _54561 = _4681 ^ _38677;
  wire _54562 = _54560 ^ _54561;
  wire _54563 = _54557 ^ _54562;
  wire _54564 = _54550 ^ _54563;
  wire _54565 = _54537 ^ _54564;
  wire _54566 = _54507 ^ _54565;
  wire _54567 = _8521 ^ _33012;
  wire _54568 = _13517 ^ _3187;
  wire _54569 = _54567 ^ _54568;
  wire _54570 = _23232 ^ _32189;
  wire _54571 = _54570 ^ _51473;
  wire _54572 = _54569 ^ _54571;
  wire _54573 = _9127 ^ _3202;
  wire _54574 = _54573 ^ uncoded_block[1721];
  wire _54575 = _54572 ^ _54574;
  wire _54576 = _54566 ^ _54575;
  wire _54577 = _54450 ^ _54576;
  wire _54578 = _3212 ^ _33031;
  wire _54579 = _3211 ^ _54578;
  wire _54580 = _54579 ^ _53577;
  wire _54581 = _2462 ^ _14571;
  wire _54582 = _54581 ^ _26387;
  wire _54583 = _13547 ^ _12429;
  wire _54584 = _23256 ^ _2472;
  wire _54585 = _54583 ^ _54584;
  wire _54586 = _54582 ^ _54585;
  wire _54587 = _54580 ^ _54586;
  wire _54588 = uncoded_block[62] ^ uncoded_block[66];
  wire _54589 = _54588 ^ _25950;
  wire _54590 = _34689 ^ _19019;
  wire _54591 = _54589 ^ _54590;
  wire _54592 = _11364 ^ _9713;
  wire _54593 = _21429 ^ _7986;
  wire _54594 = _54592 ^ _54593;
  wire _54595 = _54591 ^ _54594;
  wire _54596 = uncoded_block[112] ^ uncoded_block[116];
  wire _54597 = _54596 ^ _2497;
  wire _54598 = _24627 ^ _54597;
  wire _54599 = _1735 ^ _926;
  wire _54600 = _8577 ^ _54599;
  wire _54601 = _54598 ^ _54600;
  wire _54602 = _54595 ^ _54601;
  wire _54603 = _54587 ^ _54602;
  wire _54604 = uncoded_block[139] ^ uncoded_block[145];
  wire _54605 = _2510 ^ _54604;
  wire _54606 = _4046 ^ _18100;
  wire _54607 = _54605 ^ _54606;
  wire _54608 = _44446 ^ _25532;
  wire _54609 = _54607 ^ _54608;
  wire _54610 = uncoded_block[169] ^ uncoded_block[172];
  wire _54611 = _53604 ^ _54610;
  wire _54612 = _54611 ^ _15630;
  wire _54613 = _18110 ^ _2528;
  wire _54614 = _18111 ^ _6798;
  wire _54615 = _54613 ^ _54614;
  wire _54616 = _54612 ^ _54615;
  wire _54617 = _54609 ^ _54616;
  wire _54618 = _89 ^ _41068;
  wire _54619 = _4070 ^ _11405;
  wire _54620 = _54618 ^ _54619;
  wire _54621 = _50414 ^ _4076;
  wire _54622 = _54621 ^ _37564;
  wire _54623 = _54620 ^ _54622;
  wire _54624 = _1775 ^ _6822;
  wire _54625 = _54624 ^ _17125;
  wire _54626 = _4797 ^ _5505;
  wire _54627 = _39154 ^ _14117;
  wire _54628 = _54626 ^ _54627;
  wire _54629 = _54625 ^ _54628;
  wire _54630 = _54623 ^ _54629;
  wire _54631 = _54617 ^ _54630;
  wire _54632 = _54603 ^ _54631;
  wire _54633 = _33510 ^ _119;
  wire _54634 = _54633 ^ _42909;
  wire _54635 = _11421 ^ _5512;
  wire _54636 = _54635 ^ _53632;
  wire _54637 = _54634 ^ _54636;
  wire _54638 = _19072 ^ _134;
  wire _54639 = _54638 ^ _8047;
  wire _54640 = _999 ^ _1002;
  wire _54641 = _16644 ^ _54640;
  wire _54642 = _54639 ^ _54641;
  wire _54643 = _54637 ^ _54642;
  wire _54644 = _13619 ^ _3340;
  wire _54645 = uncoded_block[320] ^ uncoded_block[324];
  wire _54646 = _4830 ^ _54645;
  wire _54647 = _54644 ^ _54646;
  wire _54648 = _1819 ^ _13629;
  wire _54649 = _53647 ^ _3359;
  wire _54650 = _54648 ^ _54649;
  wire _54651 = _54647 ^ _54650;
  wire _54652 = _36782 ^ _3362;
  wire _54653 = uncoded_block[359] ^ uncoded_block[364];
  wire _54654 = _54653 ^ _7470;
  wire _54655 = _54652 ^ _54654;
  wire _54656 = _13093 ^ _6873;
  wire _54657 = _27334 ^ _2609;
  wire _54658 = _54656 ^ _54657;
  wire _54659 = _54655 ^ _54658;
  wire _54660 = _54651 ^ _54659;
  wire _54661 = _54643 ^ _54660;
  wire _54662 = _2612 ^ _3380;
  wire _54663 = _23779 ^ _6879;
  wire _54664 = _54662 ^ _54663;
  wire _54665 = _31870 ^ _5559;
  wire _54666 = _7487 ^ _12545;
  wire _54667 = _54665 ^ _54666;
  wire _54668 = _54664 ^ _54667;
  wire _54669 = _2629 ^ _19612;
  wire _54670 = _13112 ^ _194;
  wire _54671 = _54669 ^ _54670;
  wire _54672 = _197 ^ _6894;
  wire _54673 = _13117 ^ _21049;
  wire _54674 = _54672 ^ _54673;
  wire _54675 = _54671 ^ _54674;
  wire _54676 = _54668 ^ _54675;
  wire _54677 = _2650 ^ _13127;
  wire _54678 = _17183 ^ _54677;
  wire _54679 = _1878 ^ _16692;
  wire _54680 = _20579 ^ _54679;
  wire _54681 = _54678 ^ _54680;
  wire _54682 = uncoded_block[486] ^ uncoded_block[490];
  wire _54683 = _4897 ^ _54682;
  wire _54684 = _3422 ^ _54683;
  wire _54685 = _30167 ^ _19135;
  wire _54686 = _54685 ^ _10377;
  wire _54687 = _54684 ^ _54686;
  wire _54688 = _54681 ^ _54687;
  wire _54689 = _54676 ^ _54688;
  wire _54690 = _54661 ^ _54689;
  wire _54691 = _54632 ^ _54690;
  wire _54692 = _8705 ^ _32722;
  wire _54693 = _18206 ^ _13684;
  wire _54694 = _54692 ^ _54693;
  wire _54695 = _6929 ^ _20603;
  wire _54696 = _16215 ^ _14719;
  wire _54697 = _54695 ^ _54696;
  wire _54698 = _54694 ^ _54697;
  wire _54699 = _39608 ^ _38410;
  wire _54700 = _17217 ^ _46650;
  wire _54701 = _54699 ^ _54700;
  wire _54702 = _54698 ^ _54701;
  wire _54703 = _20110 ^ _8727;
  wire _54704 = _54703 ^ _23831;
  wire _54705 = _263 ^ _14214;
  wire _54706 = _38826 ^ _15247;
  wire _54707 = _54705 ^ _54706;
  wire _54708 = _54704 ^ _54707;
  wire _54709 = _28520 ^ _24297;
  wire _54710 = _280 ^ _6959;
  wire _54711 = _6960 ^ _31924;
  wire _54712 = _54710 ^ _54711;
  wire _54713 = _54709 ^ _54712;
  wire _54714 = _54708 ^ _54713;
  wire _54715 = _54702 ^ _54714;
  wire _54716 = _14745 ^ _3501;
  wire _54717 = _1160 ^ _5665;
  wire _54718 = _54716 ^ _54717;
  wire _54719 = _6336 ^ _6338;
  wire _54720 = _54719 ^ _40424;
  wire _54721 = _54718 ^ _54720;
  wire _54722 = _3513 ^ _5670;
  wire _54723 = _17742 ^ _1177;
  wire _54724 = _54722 ^ _54723;
  wire _54725 = _15775 ^ _10434;
  wire _54726 = uncoded_block[679] ^ uncoded_block[685];
  wire _54727 = _13731 ^ _54726;
  wire _54728 = _54725 ^ _54727;
  wire _54729 = _54724 ^ _54728;
  wire _54730 = _54721 ^ _54729;
  wire _54731 = _31076 ^ _6985;
  wire _54732 = _3529 ^ _45691;
  wire _54733 = _54731 ^ _54732;
  wire _54734 = _1191 ^ _3535;
  wire _54735 = _54734 ^ _31526;
  wire _54736 = _54733 ^ _54735;
  wire _54737 = _341 ^ _7603;
  wire _54738 = _54737 ^ _53726;
  wire _54739 = _42361 ^ _16774;
  wire _54740 = _54738 ^ _54739;
  wire _54741 = _54736 ^ _54740;
  wire _54742 = _54730 ^ _54741;
  wire _54743 = _54715 ^ _54742;
  wire _54744 = _2778 ^ _359;
  wire _54745 = _38457 ^ _54744;
  wire _54746 = _36466 ^ _6382;
  wire _54747 = _41204 ^ _54746;
  wire _54748 = _54745 ^ _54747;
  wire _54749 = _13216 ^ _20165;
  wire _54750 = _54749 ^ _18278;
  wire _54751 = _7622 ^ _11024;
  wire _54752 = uncoded_block[799] ^ uncoded_block[805];
  wire _54753 = _382 ^ _54752;
  wire _54754 = _54751 ^ _54753;
  wire _54755 = _54750 ^ _54754;
  wire _54756 = _54748 ^ _54755;
  wire _54757 = _1238 ^ _5042;
  wire _54758 = _54757 ^ _31114;
  wire _54759 = _40071 ^ _2812;
  wire _54760 = _50903 ^ _54759;
  wire _54761 = _54758 ^ _54760;
  wire _54762 = uncoded_block[837] ^ uncoded_block[845];
  wire _54763 = _26160 ^ _54762;
  wire _54764 = _54763 ^ _14298;
  wire _54765 = _6406 ^ _14300;
  wire _54766 = _11614 ^ _14302;
  wire _54767 = _54765 ^ _54766;
  wire _54768 = _54764 ^ _54767;
  wire _54769 = _54761 ^ _54768;
  wire _54770 = _54756 ^ _54769;
  wire _54771 = _22540 ^ _9953;
  wire _54772 = _31131 ^ _14821;
  wire _54773 = _54771 ^ _54772;
  wire _54774 = _9416 ^ _19735;
  wire _54775 = _2844 ^ _18311;
  wire _54776 = _54774 ^ _54775;
  wire _54777 = _54773 ^ _54776;
  wire _54778 = _44607 ^ _5093;
  wire _54779 = _3631 ^ _40484;
  wire _54780 = _9968 ^ _24837;
  wire _54781 = _54779 ^ _54780;
  wire _54782 = _54778 ^ _54781;
  wire _54783 = _54777 ^ _54782;
  wire _54784 = _4377 ^ _9433;
  wire _54785 = _13266 ^ _34496;
  wire _54786 = _54784 ^ _54785;
  wire _54787 = _34095 ^ _51646;
  wire _54788 = _54786 ^ _54787;
  wire _54789 = _50206 ^ _35305;
  wire _54790 = _21660 ^ _8855;
  wire _54791 = _11098 ^ _2882;
  wire _54792 = _54790 ^ _54791;
  wire _54793 = _54789 ^ _54792;
  wire _54794 = _54788 ^ _54793;
  wire _54795 = _54783 ^ _54794;
  wire _54796 = _54770 ^ _54795;
  wire _54797 = _54743 ^ _54796;
  wire _54798 = _54691 ^ _54797;
  wire _54799 = _22122 ^ _3666;
  wire _54800 = _22118 ^ _54799;
  wire _54801 = _7703 ^ _8299;
  wire _54802 = _22589 ^ _54801;
  wire _54803 = _54800 ^ _54802;
  wire _54804 = _8875 ^ _2127;
  wire _54805 = uncoded_block[1043] ^ uncoded_block[1049];
  wire _54806 = _502 ^ _54805;
  wire _54807 = _54804 ^ _54806;
  wire _54808 = _23966 ^ _1363;
  wire _54809 = _29412 ^ _54808;
  wire _54810 = _54807 ^ _54809;
  wire _54811 = _54803 ^ _54810;
  wire _54812 = _8889 ^ _1366;
  wire _54813 = _23502 ^ _54812;
  wire _54814 = _5158 ^ _9478;
  wire _54815 = _54814 ^ _12773;
  wire _54816 = _54813 ^ _54815;
  wire _54817 = _17363 ^ _2149;
  wire _54818 = _4440 ^ _11137;
  wire _54819 = _54817 ^ _54818;
  wire _54820 = _53810 ^ _2164;
  wire _54821 = _19309 ^ _54820;
  wire _54822 = _54819 ^ _54821;
  wire _54823 = _54816 ^ _54822;
  wire _54824 = _54811 ^ _54823;
  wire _54825 = _2165 ^ _12782;
  wire _54826 = _11147 ^ _7736;
  wire _54827 = _54825 ^ _54826;
  wire _54828 = _3718 ^ _5854;
  wire _54829 = _15894 ^ _13866;
  wire _54830 = _54828 ^ _54829;
  wire _54831 = _54827 ^ _54830;
  wire _54832 = _27528 ^ _2953;
  wire _54833 = _12794 ^ _54832;
  wire _54834 = _577 ^ _8354;
  wire _54835 = _4467 ^ _54834;
  wire _54836 = _54833 ^ _54835;
  wire _54837 = _54831 ^ _54836;
  wire _54838 = _10043 ^ _22627;
  wire _54839 = _17390 ^ _5870;
  wire _54840 = _54838 ^ _54839;
  wire _54841 = _13339 ^ _589;
  wire _54842 = _16393 ^ _35354;
  wire _54843 = _54841 ^ _54842;
  wire _54844 = _54840 ^ _54843;
  wire _54845 = _22179 ^ _7758;
  wire _54846 = _27547 ^ _54845;
  wire _54847 = _29042 ^ _23103;
  wire _54848 = _54846 ^ _54847;
  wire _54849 = _54844 ^ _54848;
  wire _54850 = _54837 ^ _54849;
  wire _54851 = _54824 ^ _54850;
  wire _54852 = _11726 ^ _3765;
  wire _54853 = uncoded_block[1223] ^ uncoded_block[1227];
  wire _54854 = _54853 ^ _13357;
  wire _54855 = _54852 ^ _54854;
  wire _54856 = _5219 ^ _1443;
  wire _54857 = _17910 ^ _2995;
  wire _54858 = _54856 ^ _54857;
  wire _54859 = _54855 ^ _54858;
  wire _54860 = _2232 ^ _24010;
  wire _54861 = _39766 ^ _19834;
  wire _54862 = _54860 ^ _54861;
  wire _54863 = _16419 ^ _3011;
  wire _54864 = _642 ^ _4531;
  wire _54865 = _54863 ^ _54864;
  wire _54866 = _54862 ^ _54865;
  wire _54867 = _54859 ^ _54866;
  wire _54868 = _10082 ^ _34177;
  wire _54869 = _21293 ^ _654;
  wire _54870 = _54869 ^ _7810;
  wire _54871 = _54868 ^ _54870;
  wire _54872 = _53861 ^ _5261;
  wire _54873 = _54872 ^ _53863;
  wire _54874 = uncoded_block[1349] ^ uncoded_block[1354];
  wire _54875 = _54874 ^ _12857;
  wire _54876 = _54875 ^ _36616;
  wire _54877 = _54873 ^ _54876;
  wire _54878 = _54871 ^ _54877;
  wire _54879 = _54867 ^ _54878;
  wire _54880 = uncoded_block[1368] ^ uncoded_block[1372];
  wire _54881 = _21306 ^ _54880;
  wire _54882 = _15966 ^ _3058;
  wire _54883 = _54881 ^ _54882;
  wire _54884 = _27590 ^ _692;
  wire _54885 = _54884 ^ _4573;
  wire _54886 = _54883 ^ _54885;
  wire _54887 = _12315 ^ _9585;
  wire _54888 = _20347 ^ _12322;
  wire _54889 = _54887 ^ _54888;
  wire _54890 = uncoded_block[1420] ^ uncoded_block[1424];
  wire _54891 = _54890 ^ _2308;
  wire _54892 = _54891 ^ _27172;
  wire _54893 = _54889 ^ _54892;
  wire _54894 = _54886 ^ _54893;
  wire _54895 = _7237 ^ _3083;
  wire _54896 = _54895 ^ _9034;
  wire _54897 = _23174 ^ _3870;
  wire _54898 = _22250 ^ _54897;
  wire _54899 = _54896 ^ _54898;
  wire _54900 = _42519 ^ _17484;
  wire _54901 = _17980 ^ _25426;
  wire _54902 = _53891 ^ _54901;
  wire _54903 = _54900 ^ _54902;
  wire _54904 = _54899 ^ _54903;
  wire _54905 = _54894 ^ _54904;
  wire _54906 = _54879 ^ _54905;
  wire _54907 = _54851 ^ _54906;
  wire _54908 = _12344 ^ _53894;
  wire _54909 = _47225 ^ _54908;
  wire _54910 = _750 ^ _19429;
  wire _54911 = _9621 ^ _7265;
  wire _54912 = _54910 ^ _54911;
  wire _54913 = _54909 ^ _54912;
  wire _54914 = _7269 ^ _3118;
  wire _54915 = _54914 ^ _53902;
  wire _54916 = uncoded_block[1541] ^ uncoded_block[1548];
  wire _54917 = _4632 ^ _54916;
  wire _54918 = _54917 ^ _24556;
  wire _54919 = _54915 ^ _54918;
  wire _54920 = _54913 ^ _54919;
  wire _54921 = _4638 ^ _3139;
  wire _54922 = _6019 ^ _1606;
  wire _54923 = _54921 ^ _54922;
  wire _54924 = _2379 ^ _4648;
  wire _54925 = _6029 ^ _15537;
  wire _54926 = _54924 ^ _54925;
  wire _54927 = _54923 ^ _54926;
  wire _54928 = _16515 ^ _45502;
  wire _54929 = _797 ^ _3151;
  wire _54930 = _54928 ^ _54929;
  wire _54931 = uncoded_block[1606] ^ uncoded_block[1611];
  wire _54932 = _54931 ^ _7908;
  wire _54933 = _6679 ^ _7911;
  wire _54934 = _54932 ^ _54933;
  wire _54935 = _54930 ^ _54934;
  wire _54936 = _54927 ^ _54935;
  wire _54937 = _54920 ^ _54936;
  wire _54938 = _20899 ^ _5389;
  wire _54939 = _1642 ^ _10755;
  wire _54940 = _54939 ^ _53933;
  wire _54941 = _54938 ^ _54940;
  wire _54942 = _12960 ^ _15566;
  wire _54943 = _41406 ^ _54942;
  wire _54944 = _8521 ^ _832;
  wire _54945 = _54944 ^ _38681;
  wire _54946 = _54943 ^ _54945;
  wire _54947 = _54941 ^ _54946;
  wire _54948 = _14543 ^ _837;
  wire _54949 = _7331 ^ _2430;
  wire _54950 = _54948 ^ _54949;
  wire _54951 = _24137 ^ _3976;
  wire _54952 = _44408 ^ _852;
  wire _54953 = _54951 ^ _54952;
  wire _54954 = _54950 ^ _54953;
  wire _54955 = _7944 ^ _7946;
  wire _54956 = _54955 ^ uncoded_block[1722];
  wire _54957 = _54954 ^ _54956;
  wire _54958 = _54947 ^ _54957;
  wire _54959 = _54937 ^ _54958;
  wire _54960 = _54907 ^ _54959;
  wire _54961 = _54798 ^ _54960;
  wire _54962 = _41 ^ _17077;
  wire _54963 = _54962 ^ _51809;
  wire _54964 = _54963 ^ _51811;
  wire _54965 = _11918 ^ _33909;
  wire _54966 = _23272 ^ _54965;
  wire _54967 = _53067 ^ _54966;
  wire _54968 = _54964 ^ _54967;
  wire _54969 = _53371 ^ _54968;
  wire _54970 = _52371 ^ _24182;
  wire _54971 = _54970 ^ _16108;
  wire _54972 = _52120 ^ _52379;
  wire _54973 = _54971 ^ _54972;
  wire _54974 = _51509 ^ _51512;
  wire _54975 = _17613 ^ _104;
  wire _54976 = _53083 ^ _54975;
  wire _54977 = _54974 ^ _54976;
  wire _54978 = _54973 ^ _54977;
  wire _54979 = uncoded_block[236] ^ uncoded_block[242];
  wire _54980 = _968 ^ _54979;
  wire _54981 = _51516 ^ _54980;
  wire _54982 = _50768 ^ _13607;
  wire _54983 = _54981 ^ _54982;
  wire _54984 = _54983 ^ _51840;
  wire _54985 = _54978 ^ _54984;
  wire _54986 = _54969 ^ _54985;
  wire _54987 = _33536 ^ _50070;
  wire _54988 = _46219 ^ _54001;
  wire _54989 = _54987 ^ _54988;
  wire _54990 = _53398 ^ _54989;
  wire _54991 = _52419 ^ _27747;
  wire _54992 = _52151 ^ _48126;
  wire _54993 = _54991 ^ _54992;
  wire _54994 = _53405 ^ _54993;
  wire _54995 = _54990 ^ _54994;
  wire _54996 = _49241 ^ _52157;
  wire _54997 = _13662 ^ _9283;
  wire _54998 = _54997 ^ _51556;
  wire _54999 = _54996 ^ _54998;
  wire _55000 = _54021 ^ _51881;
  wire _55001 = _51562 ^ _55000;
  wire _55002 = _54999 ^ _55001;
  wire _55003 = _52446 ^ _46261;
  wire _55004 = _46259 ^ _55003;
  wire _55005 = _51570 ^ _55004;
  wire _55006 = _55002 ^ _55005;
  wire _55007 = _54995 ^ _55006;
  wire _55008 = _54986 ^ _55007;
  wire _55009 = _42668 ^ _3481;
  wire _55010 = _46269 ^ _55009;
  wire _55011 = _46272 ^ _14219;
  wire _55012 = _51900 ^ _51904;
  wire _55013 = _55011 ^ _55012;
  wire _55014 = _55010 ^ _55013;
  wire _55015 = _1163 ^ _4972;
  wire _55016 = _51905 ^ _55015;
  wire _55017 = _298 ^ _52190;
  wire _55018 = _55016 ^ _55017;
  wire _55019 = _1971 ^ _322;
  wire _55020 = _55019 ^ _15283;
  wire _55021 = _54051 ^ _55020;
  wire _55022 = _55018 ^ _55021;
  wire _55023 = _55014 ^ _55022;
  wire _55024 = _52477 ^ _25672;
  wire _55025 = _4999 ^ _6367;
  wire _55026 = _6999 ^ _46300;
  wire _55027 = _55025 ^ _55026;
  wire _55028 = _55024 ^ _55027;
  wire _55029 = _46302 ^ _18736;
  wire _55030 = _46306 ^ _46308;
  wire _55031 = _55029 ^ _55030;
  wire _55032 = _55028 ^ _55031;
  wire _55033 = _46309 ^ _52210;
  wire _55034 = _51615 ^ _1234;
  wire _55035 = _55033 ^ _55034;
  wire _55036 = _2022 ^ _34062;
  wire _55037 = _55036 ^ _53460;
  wire _55038 = _55037 ^ _53462;
  wire _55039 = _55035 ^ _55038;
  wire _55040 = _55032 ^ _55039;
  wire _55041 = _55023 ^ _55040;
  wire _55042 = uncoded_block[882] ^ uncoded_block[886];
  wire _55043 = _3608 ^ _55042;
  wire _55044 = _52223 ^ _55043;
  wire _55045 = _50917 ^ _30690;
  wire _55046 = _55044 ^ _55045;
  wire _55047 = _53469 ^ _55046;
  wire _55048 = _25728 ^ _52231;
  wire _55049 = _3629 ^ _8259;
  wire _55050 = _55049 ^ _51954;
  wire _55051 = _55048 ^ _55050;
  wire _55052 = _55051 ^ _53480;
  wire _55053 = _55047 ^ _55052;
  wire _55054 = _53486 ^ _54102;
  wire _55055 = _51333 ^ _7117;
  wire _55056 = _53230 ^ _55055;
  wire _55057 = _34932 ^ _46370;
  wire _55058 = _55056 ^ _55057;
  wire _55059 = _46371 ^ _25777;
  wire _55060 = _48266 ^ _46377;
  wire _55061 = _55059 ^ _55060;
  wire _55062 = _55058 ^ _55061;
  wire _55063 = _55054 ^ _55062;
  wire _55064 = _55053 ^ _55063;
  wire _55065 = _55041 ^ _55064;
  wire _55066 = _55008 ^ _55065;
  wire _55067 = _46378 ^ _51988;
  wire _55068 = _30329 ^ _46389;
  wire _55069 = _48272 ^ _55068;
  wire _55070 = _55067 ^ _55069;
  wire _55071 = _2185 ^ _46391;
  wire _55072 = _55071 ^ _3735;
  wire _55073 = _51996 ^ _32064;
  wire _55074 = _55073 ^ _46398;
  wire _55075 = _55072 ^ _55074;
  wire _55076 = _55070 ^ _55075;
  wire _55077 = _9508 ^ _10612;
  wire _55078 = _2203 ^ _2206;
  wire _55079 = _55077 ^ _55078;
  wire _55080 = _51694 ^ _28298;
  wire _55081 = _55079 ^ _55080;
  wire _55082 = _2220 ^ _19347;
  wire _55083 = _55082 ^ _46409;
  wire _55084 = _17911 ^ _8385;
  wire _55085 = _52010 ^ _55084;
  wire _55086 = _55083 ^ _55085;
  wire _55087 = _55081 ^ _55086;
  wire _55088 = _55076 ^ _55087;
  wire _55089 = _5232 ^ _34564;
  wire _55090 = _55089 ^ _52285;
  wire _55091 = _55090 ^ _53518;
  wire _55092 = _2283 ^ _3054;
  wire _55093 = _55092 ^ _52033;
  wire _55094 = _55093 ^ _52040;
  wire _55095 = _53522 ^ _55094;
  wire _55096 = _55091 ^ _55095;
  wire _55097 = _55088 ^ _55096;
  wire _55098 = _4572 ^ _2299;
  wire _55099 = _55098 ^ _48340;
  wire _55100 = _3075 ^ _1531;
  wire _55101 = _53529 ^ _55100;
  wire _55102 = _55099 ^ _55101;
  wire _55103 = _49443 ^ _52309;
  wire _55104 = _55102 ^ _55103;
  wire _55105 = _40603 ^ _3100;
  wire _55106 = _47599 ^ _55105;
  wire _55107 = _19888 ^ _39039;
  wire _55108 = _55106 ^ _55107;
  wire _55109 = _55108 ^ _53545;
  wire _55110 = _55104 ^ _55109;
  wire _55111 = _10720 ^ _32972;
  wire _55112 = _55111 ^ _52322;
  wire _55113 = _52639 ^ _46480;
  wire _55114 = _24102 ^ _10163;
  wire _55115 = _55114 ^ _50688;
  wire _55116 = _55113 ^ _55115;
  wire _55117 = _55112 ^ _55116;
  wire _55118 = _52326 ^ _52329;
  wire _55119 = _52080 ^ _13501;
  wire _55120 = _52330 ^ _55119;
  wire _55121 = _55118 ^ _55120;
  wire _55122 = _55117 ^ _55121;
  wire _55123 = _55110 ^ _55122;
  wire _55124 = _55097 ^ _55123;
  wire _55125 = _17029 ^ _25024;
  wire _55126 = _10761 ^ _52088;
  wire _55127 = _19939 ^ _33012;
  wire _55128 = _55126 ^ _55127;
  wire _55129 = _55125 ^ _55128;
  wire _55130 = _19476 ^ _32190;
  wire _55131 = _6068 ^ _1672;
  wire _55132 = _851 ^ _854;
  wire _55133 = _55131 ^ _55132;
  wire _55134 = _55130 ^ _55133;
  wire _55135 = _55129 ^ _55134;
  wire _55136 = _55135 ^ _21402;
  wire _55137 = _55124 ^ _55136;
  wire _55138 = _55066 ^ _55137;
  wire _55139 = _6724 ^ _2454;
  wire _55140 = _49148 ^ _55139;
  wire _55141 = _46150 ^ _11343;
  wire _55142 = _11344 ^ _6732;
  wire _55143 = _55141 ^ _55142;
  wire _55144 = _55140 ^ _55143;
  wire _55145 = _39103 ^ _51486;
  wire _55146 = _6742 ^ _9705;
  wire _55147 = uncoded_block[77] ^ uncoded_block[81];
  wire _55148 = _10244 ^ _55147;
  wire _55149 = _55146 ^ _55148;
  wire _55150 = _55145 ^ _55149;
  wire _55151 = _55144 ^ _55150;
  wire _55152 = uncoded_block[88] ^ uncoded_block[95];
  wire _55153 = _55152 ^ _15101;
  wire _55154 = _54962 ^ _55153;
  wire _55155 = _6120 ^ _9720;
  wire _55156 = _46171 ^ _13016;
  wire _55157 = _55155 ^ _55156;
  wire _55158 = _55154 ^ _55157;
  wire _55159 = _23720 ^ _4043;
  wire _55160 = _49174 ^ _55159;
  wire _55161 = _12460 ^ _2514;
  wire _55162 = _6785 ^ _46182;
  wire _55163 = _55161 ^ _55162;
  wire _55164 = _55160 ^ _55163;
  wire _55165 = _55158 ^ _55164;
  wire _55166 = _55151 ^ _55165;
  wire _55167 = _2521 ^ _940;
  wire _55168 = _11395 ^ _22368;
  wire _55169 = _55167 ^ _55168;
  wire _55170 = _51509 ^ _46188;
  wire _55171 = _55169 ^ _55170;
  wire _55172 = _28043 ^ _46189;
  wire _55173 = _23296 ^ _5497;
  wire _55174 = _55172 ^ _55173;
  wire _55175 = _2545 ^ _18123;
  wire _55176 = _55175 ^ _51831;
  wire _55177 = _55174 ^ _55176;
  wire _55178 = _55171 ^ _55177;
  wire _55179 = _49197 ^ _6828;
  wire _55180 = _6187 ^ _7440;
  wire _55181 = _55180 ^ _53986;
  wire _55182 = _55179 ^ _55181;
  wire _55183 = _11967 ^ _49687;
  wire _55184 = _55183 ^ _42917;
  wire _55185 = _8636 ^ _14652;
  wire _55186 = _6845 ^ _22866;
  wire _55187 = _55185 ^ _55186;
  wire _55188 = _55184 ^ _55187;
  wire _55189 = _55182 ^ _55188;
  wire _55190 = _55178 ^ _55189;
  wire _55191 = _55166 ^ _55190;
  wire _55192 = uncoded_block[319] ^ uncoded_block[325];
  wire _55193 = _15671 ^ _55192;
  wire _55194 = _55193 ^ _10320;
  wire _55195 = _15172 ^ _6857;
  wire _55196 = _55195 ^ _51175;
  wire _55197 = _55194 ^ _55196;
  wire _55198 = _8652 ^ _21028;
  wire _55199 = _2602 ^ _35170;
  wire _55200 = _55198 ^ _55199;
  wire _55201 = _31862 ^ _4858;
  wire _55202 = _46987 ^ _55201;
  wire _55203 = _55200 ^ _55202;
  wire _55204 = _55197 ^ _55203;
  wire _55205 = _51855 ^ _52419;
  wire _55206 = _1051 ^ _2629;
  wire _55207 = _55206 ^ _21044;
  wire _55208 = _55205 ^ _55207;
  wire _55209 = _2633 ^ _14163;
  wire _55210 = _6254 ^ _205;
  wire _55211 = _55209 ^ _55210;
  wire _55212 = _24716 ^ _208;
  wire _55213 = _6261 ^ _4181;
  wire _55214 = _55212 ^ _55213;
  wire _55215 = _55211 ^ _55214;
  wire _55216 = _55208 ^ _55215;
  wire _55217 = _55204 ^ _55216;
  wire _55218 = _26944 ^ _11494;
  wire _55219 = _51871 ^ _55218;
  wire _55220 = _2659 ^ _12577;
  wire _55221 = _55220 ^ _54021;
  wire _55222 = _55219 ^ _55221;
  wire _55223 = _11508 ^ _4208;
  wire _55224 = _51881 ^ _55223;
  wire _55225 = _3446 ^ _46254;
  wire _55226 = _55224 ^ _55225;
  wire _55227 = _55222 ^ _55226;
  wire _55228 = uncoded_block[546] ^ uncoded_block[550];
  wire _55229 = _55228 ^ _3459;
  wire _55230 = _6304 ^ _6940;
  wire _55231 = _55229 ^ _55230;
  wire _55232 = _52170 ^ _55231;
  wire _55233 = _51571 ^ _51578;
  wire _55234 = _13170 ^ _33602;
  wire _55235 = _55233 ^ _55234;
  wire _55236 = _55232 ^ _55235;
  wire _55237 = _55227 ^ _55236;
  wire _55238 = _55217 ^ _55237;
  wire _55239 = _55191 ^ _55238;
  wire _55240 = _4953 ^ _11535;
  wire _55241 = _55240 ^ _19165;
  wire _55242 = _5652 ^ _16238;
  wire _55243 = _12618 ^ _1156;
  wire _55244 = _55242 ^ _55243;
  wire _55245 = _55241 ^ _55244;
  wire _55246 = _17735 ^ _55015;
  wire _55247 = _41172 ^ _32755;
  wire _55248 = _55246 ^ _55247;
  wire _55249 = _55245 ^ _55248;
  wire _55250 = _3515 ^ _50507;
  wire _55251 = _8180 ^ _322;
  wire _55252 = _49772 ^ _55251;
  wire _55253 = _55250 ^ _55252;
  wire _55254 = _1186 ^ _18719;
  wire _55255 = _55254 ^ _52477;
  wire _55256 = _12647 ^ _6367;
  wire _55257 = _3537 ^ _55256;
  wire _55258 = _55255 ^ _55257;
  wire _55259 = _55253 ^ _55258;
  wire _55260 = _55249 ^ _55259;
  wire _55261 = _6999 ^ _7603;
  wire _55262 = _55261 ^ _38862;
  wire _55263 = _2774 ^ _12107;
  wire _55264 = _2002 ^ _5017;
  wire _55265 = _55263 ^ _55264;
  wire _55266 = _55262 ^ _55265;
  wire _55267 = _5019 ^ _2783;
  wire _55268 = _55267 ^ _49307;
  wire _55269 = _55268 ^ _49311;
  wire _55270 = _55266 ^ _55269;
  wire _55271 = _374 ^ _8223;
  wire _55272 = _26589 ^ _34062;
  wire _55273 = _55271 ^ _55272;
  wire _55274 = uncoded_block[818] ^ uncoded_block[823];
  wire _55275 = _5046 ^ _55274;
  wire _55276 = _5730 ^ _55275;
  wire _55277 = _55273 ^ _55276;
  wire _55278 = _14291 ^ _27846;
  wire _55279 = _12138 ^ _7043;
  wire _55280 = _55278 ^ _55279;
  wire _55281 = _5058 ^ _11609;
  wire _55282 = _12141 ^ _7644;
  wire _55283 = _55281 ^ _55282;
  wire _55284 = _55280 ^ _55283;
  wire _55285 = _55277 ^ _55284;
  wire _55286 = _55270 ^ _55285;
  wire _55287 = _55260 ^ _55286;
  wire _55288 = _30680 ^ _6410;
  wire _55289 = _55288 ^ _22087;
  wire _55290 = _2828 ^ _5752;
  wire _55291 = _11621 ^ _3613;
  wire _55292 = _55290 ^ _55291;
  wire _55293 = _55289 ^ _55292;
  wire _55294 = _14827 ^ _5085;
  wire _55295 = _1278 ^ _429;
  wire _55296 = _55294 ^ _55295;
  wire _55297 = _1282 ^ _52231;
  wire _55298 = _55296 ^ _55297;
  wire _55299 = _55293 ^ _55298;
  wire _55300 = _24832 ^ _2076;
  wire _55301 = _2857 ^ _4377;
  wire _55302 = _55300 ^ _55301;
  wire _55303 = _55302 ^ _54090;
  wire _55304 = _11646 ^ _467;
  wire _55305 = _46348 ^ _55304;
  wire _55306 = _468 ^ _13821;
  wire _55307 = _55306 ^ _7686;
  wire _55308 = _55305 ^ _55307;
  wire _55309 = _55303 ^ _55308;
  wire _55310 = _55299 ^ _55309;
  wire _55311 = _7689 ^ _24853;
  wire _55312 = _16338 ^ _8293;
  wire _55313 = _55311 ^ _55312;
  wire _55314 = _55313 ^ _52539;
  wire _55315 = uncoded_block[1017] ^ uncoded_block[1022];
  wire _55316 = _9996 ^ _55315;
  wire _55317 = _9455 ^ _3675;
  wire _55318 = _55316 ^ _55317;
  wire _55319 = _4418 ^ _3678;
  wire _55320 = _2910 ^ _45005;
  wire _55321 = _55319 ^ _55320;
  wire _55322 = _55318 ^ _55321;
  wire _55323 = _55314 ^ _55322;
  wire _55324 = _3684 ^ _14357;
  wire _55325 = _21681 ^ _55324;
  wire _55326 = _3689 ^ _12217;
  wire _55327 = _5832 ^ _5163;
  wire _55328 = _55326 ^ _55327;
  wire _55329 = _55325 ^ _55328;
  wire _55330 = _49369 ^ _20759;
  wire _55331 = _3707 ^ _550;
  wire _55332 = _8911 ^ _55331;
  wire _55333 = _55330 ^ _55332;
  wire _55334 = _55329 ^ _55333;
  wire _55335 = _55323 ^ _55334;
  wire _55336 = _55310 ^ _55335;
  wire _55337 = _55287 ^ _55336;
  wire _55338 = _55239 ^ _55337;
  wire _55339 = _19313 ^ _8339;
  wire _55340 = uncoded_block[1126] ^ uncoded_block[1138];
  wire _55341 = _14376 ^ _55340;
  wire _55342 = _55339 ^ _55341;
  wire _55343 = uncoded_block[1140] ^ uncoded_block[1149];
  wire _55344 = _55343 ^ _2185;
  wire _55345 = _55344 ^ _46392;
  wire _55346 = _55342 ^ _55345;
  wire _55347 = _3734 ^ _21248;
  wire _55348 = _2192 ^ _5872;
  wire _55349 = _55347 ^ _55348;
  wire _55350 = _27539 ^ _592;
  wire _55351 = _2196 ^ _13346;
  wire _55352 = _55350 ^ _55351;
  wire _55353 = _55349 ^ _55352;
  wire _55354 = _55346 ^ _55353;
  wire _55355 = _24910 ^ _8951;
  wire _55356 = _55355 ^ _52003;
  wire _55357 = _2218 ^ _28298;
  wire _55358 = _55356 ^ _55357;
  wire _55359 = _30352 ^ _5891;
  wire _55360 = uncoded_block[1233] ^ uncoded_block[1239];
  wire _55361 = _3769 ^ _55360;
  wire _55362 = _55359 ^ _55361;
  wire _55363 = _53270 ^ _13367;
  wire _55364 = _55362 ^ _55363;
  wire _55365 = _55358 ^ _55364;
  wire _55366 = _55354 ^ _55365;
  wire _55367 = _32082 ^ _1456;
  wire _55368 = _3786 ^ _39379;
  wire _55369 = _55367 ^ _55368;
  wire _55370 = uncoded_block[1292] ^ uncoded_block[1299];
  wire _55371 = _13380 ^ _55370;
  wire _55372 = _53279 ^ _55371;
  wire _55373 = _55369 ^ _55372;
  wire _55374 = _3018 ^ _649;
  wire _55375 = uncoded_block[1313] ^ uncoded_block[1317];
  wire _55376 = _8407 ^ _55375;
  wire _55377 = _55374 ^ _55376;
  wire _55378 = _12287 ^ _1487;
  wire _55379 = _55378 ^ _17935;
  wire _55380 = _55377 ^ _55379;
  wire _55381 = _55373 ^ _55380;
  wire _55382 = uncoded_block[1343] ^ uncoded_block[1351];
  wire _55383 = _14440 ^ _55382;
  wire _55384 = _37817 ^ _55383;
  wire _55385 = _55384 ^ _46439;
  wire _55386 = uncoded_block[1367] ^ uncoded_block[1374];
  wire _55387 = _55386 ^ _49071;
  wire _55388 = _55387 ^ _46446;
  wire _55389 = _27164 ^ _32940;
  wire _55390 = _55388 ^ _55389;
  wire _55391 = _55385 ^ _55390;
  wire _55392 = _55381 ^ _55391;
  wire _55393 = _55366 ^ _55392;
  wire _55394 = _5961 ^ _21780;
  wire _55395 = _55394 ^ _55100;
  wire _55396 = _10124 ^ _17470;
  wire _55397 = _55396 ^ _51042;
  wire _55398 = _55395 ^ _55397;
  wire _55399 = _5309 ^ _726;
  wire _55400 = _54167 ^ _55399;
  wire _55401 = _35423 ^ _23179;
  wire _55402 = _47599 ^ _55401;
  wire _55403 = _55400 ^ _55402;
  wire _55404 = _55398 ^ _55403;
  wire _55405 = uncoded_block[1489] ^ uncoded_block[1496];
  wire _55406 = _55405 ^ _2352;
  wire _55407 = _51748 ^ _55406;
  wire _55408 = _15516 ^ _32142;
  wire _55409 = _55407 ^ _55408;
  wire _55410 = _6642 ^ _11267;
  wire _55411 = _55410 ^ _24993;
  wire _55412 = _55411 ^ _55111;
  wire _55413 = _55409 ^ _55412;
  wire _55414 = _55404 ^ _55413;
  wire _55415 = _51759 ^ _2368;
  wire _55416 = uncoded_block[1559] ^ uncoded_block[1564];
  wire _55417 = _3914 ^ _55416;
  wire _55418 = _54187 ^ _55417;
  wire _55419 = _55415 ^ _55418;
  wire _55420 = uncoded_block[1581] ^ uncoded_block[1593];
  wire _55421 = _2380 ^ _55420;
  wire _55422 = _46481 ^ _55421;
  wire _55423 = _55422 ^ _52075;
  wire _55424 = _55419 ^ _55423;
  wire _55425 = _3154 ^ _3157;
  wire _55426 = _55425 ^ _52653;
  wire _55427 = _14006 ^ _1639;
  wire _55428 = _55427 ^ _52080;
  wire _55429 = _55426 ^ _55428;
  wire _55430 = _2408 ^ _7921;
  wire _55431 = _55430 ^ _17029;
  wire _55432 = _25024 ^ _41411;
  wire _55433 = _55431 ^ _55432;
  wire _55434 = _55429 ^ _55433;
  wire _55435 = _55424 ^ _55434;
  wire _55436 = _55414 ^ _55435;
  wire _55437 = _55393 ^ _55436;
  wire _55438 = _3186 ^ _23671;
  wire _55439 = _49985 ^ _55438;
  wire _55440 = _3191 ^ _52667;
  wire _55441 = _55439 ^ _55440;
  wire _55442 = _54215 ^ _855;
  wire _55443 = _15064 ^ _55442;
  wire _55444 = _55443 ^ _861;
  wire _55445 = _55441 ^ _55444;
  wire _55446 = _55437 ^ _55445;
  wire _55447 = _55338 ^ _55446;
  wire _55448 = _3209 ^ _4712;
  wire _55449 = _14560 ^ _5423;
  wire _55450 = _55448 ^ _55449;
  wire _55451 = _53574 ^ _10791;
  wire _55452 = _22790 ^ _21412;
  wire _55453 = _55451 ^ _55452;
  wire _55454 = _55450 ^ _55453;
  wire _55455 = uncoded_block[33] ^ uncoded_block[39];
  wire _55456 = uncoded_block[45] ^ uncoded_block[50];
  wire _55457 = _55455 ^ _55456;
  wire _55458 = _25948 ^ _9156;
  wire _55459 = _55457 ^ _55458;
  wire _55460 = _6745 ^ _5443;
  wire _55461 = _55460 ^ _41041;
  wire _55462 = _55459 ^ _55461;
  wire _55463 = _55454 ^ _55462;
  wire _55464 = _11364 ^ _18077;
  wire _55465 = _15603 ^ _21429;
  wire _55466 = _55464 ^ _55465;
  wire _55467 = _17084 ^ _36311;
  wire _55468 = _55466 ^ _55467;
  wire _55469 = _33056 ^ _2498;
  wire _55470 = _10821 ^ _1730;
  wire _55471 = _55469 ^ _55470;
  wire _55472 = _25075 ^ _30945;
  wire _55473 = _11376 ^ _55472;
  wire _55474 = _55471 ^ _55473;
  wire _55475 = _55468 ^ _55474;
  wire _55476 = _55463 ^ _55475;
  wire _55477 = uncoded_block[149] ^ uncoded_block[152];
  wire _55478 = _6780 ^ _55477;
  wire _55479 = _4048 ^ _15118;
  wire _55480 = _55478 ^ _55479;
  wire _55481 = _74 ^ _3276;
  wire _55482 = _1752 ^ _10270;
  wire _55483 = _55481 ^ _55482;
  wire _55484 = _55480 ^ _55483;
  wire _55485 = _7408 ^ _18111;
  wire _55486 = _8010 ^ _55485;
  wire _55487 = _6158 ^ _8600;
  wire _55488 = _54618 ^ _55487;
  wire _55489 = _55486 ^ _55488;
  wire _55490 = _55484 ^ _55489;
  wire _55491 = uncoded_block[218] ^ uncoded_block[223];
  wire _55492 = _956 ^ _55491;
  wire _55493 = _8608 ^ _4791;
  wire _55494 = _55492 ^ _55493;
  wire _55495 = _53390 ^ _44060;
  wire _55496 = _55494 ^ _55495;
  wire _55497 = _20996 ^ _11955;
  wire _55498 = _38753 ^ _6186;
  wire _55499 = _55497 ^ _55498;
  wire _55500 = _55496 ^ _55499;
  wire _55501 = _55490 ^ _55500;
  wire _55502 = _55476 ^ _55501;
  wire _55503 = _21472 ^ _5512;
  wire _55504 = _6189 ^ _55503;
  wire _55505 = _4103 ^ _5515;
  wire _55506 = _55505 ^ _54638;
  wire _55507 = _55504 ^ _55506;
  wire _55508 = _992 ^ _42916;
  wire _55509 = _8051 ^ _143;
  wire _55510 = _55508 ^ _55509;
  wire _55511 = _3341 ^ _6850;
  wire _55512 = _24218 ^ _55511;
  wire _55513 = _55510 ^ _55512;
  wire _55514 = _55507 ^ _55513;
  wire _55515 = _21947 ^ _2584;
  wire _55516 = _2586 ^ _5536;
  wire _55517 = _55515 ^ _55516;
  wire _55518 = uncoded_block[340] ^ uncoded_block[343];
  wire _55519 = _55518 ^ _4131;
  wire _55520 = _6215 ^ _55519;
  wire _55521 = _55517 ^ _55520;
  wire _55522 = _161 ^ _36782;
  wire _55523 = _3362 ^ _35170;
  wire _55524 = _55522 ^ _55523;
  wire _55525 = _42282 ^ _28838;
  wire _55526 = _45618 ^ _55525;
  wire _55527 = _55524 ^ _55526;
  wire _55528 = _55521 ^ _55527;
  wire _55529 = _55514 ^ _55528;
  wire _55530 = uncoded_block[378] ^ uncoded_block[381];
  wire _55531 = _55530 ^ _4858;
  wire _55532 = _4149 ^ _6879;
  wire _55533 = _55531 ^ _55532;
  wire _55534 = _46613 ^ _9808;
  wire _55535 = _55533 ^ _55534;
  wire _55536 = _12545 ^ _4867;
  wire _55537 = _1055 ^ _13112;
  wire _55538 = _55536 ^ _55537;
  wire _55539 = _4165 ^ _9817;
  wire _55540 = _55538 ^ _55539;
  wire _55541 = _55535 ^ _55540;
  wire _55542 = _4169 ^ _19115;
  wire _55543 = _23792 ^ _55542;
  wire _55544 = _9275 ^ _6259;
  wire _55545 = _19621 ^ _1076;
  wire _55546 = _55544 ^ _55545;
  wire _55547 = _55543 ^ _55546;
  wire _55548 = _4181 ^ _2654;
  wire _55549 = _6906 ^ _11494;
  wire _55550 = _55548 ^ _55549;
  wire _55551 = _3423 ^ _54682;
  wire _55552 = _3422 ^ _55551;
  wire _55553 = _55550 ^ _55552;
  wire _55554 = _55547 ^ _55553;
  wire _55555 = _55541 ^ _55554;
  wire _55556 = _55529 ^ _55555;
  wire _55557 = _55502 ^ _55556;
  wire _55558 = _42965 ^ _19135;
  wire _55559 = _55558 ^ _18201;
  wire _55560 = _32722 ^ _19638;
  wire _55561 = _4206 ^ _55560;
  wire _55562 = _55559 ^ _55561;
  wire _55563 = _10947 ^ _13684;
  wire _55564 = _55563 ^ _16214;
  wire _55565 = _24278 ^ _14199;
  wire _55566 = _55564 ^ _55565;
  wire _55567 = _55562 ^ _55566;
  wire _55568 = uncoded_block[547] ^ uncoded_block[557];
  wire _55569 = _55568 ^ _5633;
  wire _55570 = _1910 ^ _55569;
  wire _55571 = _3465 ^ _8727;
  wire _55572 = uncoded_block[577] ^ uncoded_block[581];
  wire _55573 = _1931 ^ _55572;
  wire _55574 = _55571 ^ _55573;
  wire _55575 = _55570 ^ _55574;
  wire _55576 = _2696 ^ _270;
  wire _55577 = _55576 ^ _15248;
  wire _55578 = uncoded_block[598] ^ uncoded_block[604];
  wire _55579 = _55578 ^ _6323;
  wire _55580 = _21098 ^ _281;
  wire _55581 = _55579 ^ _55580;
  wire _55582 = _55577 ^ _55581;
  wire _55583 = _55575 ^ _55582;
  wire _55584 = _55567 ^ _55583;
  wire _55585 = _1946 ^ _4964;
  wire _55586 = _55585 ^ _33182;
  wire _55587 = uncoded_block[634] ^ uncoded_block[637];
  wire _55588 = _55587 ^ _6336;
  wire _55589 = uncoded_block[644] ^ uncoded_block[648];
  wire _55590 = _55589 ^ _10427;
  wire _55591 = _55588 ^ _55590;
  wire _55592 = _55586 ^ _55591;
  wire _55593 = _3513 ^ _7582;
  wire _55594 = _311 ^ _10434;
  wire _55595 = _55593 ^ _55594;
  wire _55596 = _12089 ^ _13735;
  wire _55597 = _33622 ^ _55596;
  wire _55598 = _55595 ^ _55597;
  wire _55599 = _55592 ^ _55598;
  wire _55600 = uncoded_block[700] ^ uncoded_block[705];
  wire _55601 = _19195 ^ _55600;
  wire _55602 = _19685 ^ _55601;
  wire _55603 = _33205 ^ _17266;
  wire _55604 = _340 ^ _8198;
  wire _55605 = _55603 ^ _55604;
  wire _55606 = _55602 ^ _55605;
  wire _55607 = _14774 ^ _349;
  wire _55608 = _350 ^ _5699;
  wire _55609 = _55607 ^ _55608;
  wire _55610 = _5703 ^ _38457;
  wire _55611 = _55609 ^ _55610;
  wire _55612 = _55606 ^ _55611;
  wire _55613 = _55599 ^ _55612;
  wire _55614 = _55584 ^ _55613;
  wire _55615 = _43792 ^ _10470;
  wire _55616 = _14781 ^ _55615;
  wire _55617 = _11587 ^ _5714;
  wire _55618 = _55616 ^ _55617;
  wire _55619 = uncoded_block[785] ^ uncoded_block[793];
  wire _55620 = _12669 ^ _55619;
  wire _55621 = _14282 ^ _2801;
  wire _55622 = _55620 ^ _55621;
  wire _55623 = _20178 ^ _14801;
  wire _55624 = _55622 ^ _55623;
  wire _55625 = _55618 ^ _55624;
  wire _55626 = _2029 ^ _40071;
  wire _55627 = _44958 ^ _55626;
  wire _55628 = _5734 ^ _400;
  wire _55629 = uncoded_block[838] ^ uncoded_block[843];
  wire _55630 = _13781 ^ _55629;
  wire _55631 = _55628 ^ _55630;
  wire _55632 = _55627 ^ _55631;
  wire _55633 = _9943 ^ _11048;
  wire _55634 = _14300 ^ _4344;
  wire _55635 = _55633 ^ _55634;
  wire _55636 = _4346 ^ _16303;
  wire _55637 = _8820 ^ _7660;
  wire _55638 = _55636 ^ _55637;
  wire _55639 = _55635 ^ _55638;
  wire _55640 = _55632 ^ _55639;
  wire _55641 = _55625 ^ _55640;
  wire _55642 = _4356 ^ _5760;
  wire _55643 = _18311 ^ _12708;
  wire _55644 = _55643 ^ _54411;
  wire _55645 = _55642 ^ _55644;
  wire _55646 = _2076 ^ _2857;
  wire _55647 = _1294 ^ _55646;
  wire _55648 = uncoded_block[930] ^ uncoded_block[934];
  wire _55649 = _55648 ^ _7080;
  wire _55650 = _453 ^ _2865;
  wire _55651 = _55649 ^ _55650;
  wire _55652 = _55647 ^ _55651;
  wire _55653 = _55645 ^ _55652;
  wire _55654 = _54785 ^ _34095;
  wire _55655 = uncoded_block[971] ^ uncoded_block[981];
  wire _55656 = _11087 ^ _55655;
  wire _55657 = _50203 ^ _55656;
  wire _55658 = _55654 ^ _55657;
  wire _55659 = _50567 ^ _2105;
  wire _55660 = _17340 ^ _28241;
  wire _55661 = _55659 ^ _55660;
  wire _55662 = _4404 ^ _6459;
  wire _55663 = _13283 ^ _19763;
  wire _55664 = _55662 ^ _55663;
  wire _55665 = _55661 ^ _55664;
  wire _55666 = _55658 ^ _55665;
  wire _55667 = _55653 ^ _55666;
  wire _55668 = _55641 ^ _55667;
  wire _55669 = _55614 ^ _55668;
  wire _55670 = _55557 ^ _55669;
  wire _55671 = _12750 ^ _5138;
  wire _55672 = _55671 ^ _20232;
  wire _55673 = _2129 ^ _1356;
  wire _55674 = _43098 ^ _55673;
  wire _55675 = _55672 ^ _55674;
  wire _55676 = _1359 ^ _1363;
  wire _55677 = _17355 ^ _55676;
  wire _55678 = _33294 ^ _18355;
  wire _55679 = _55677 ^ _55678;
  wire _55680 = _55675 ^ _55679;
  wire _55681 = _17362 ^ _10575;
  wire _55682 = _8323 ^ _55681;
  wire _55683 = _3696 ^ _536;
  wire _55684 = _55683 ^ _19309;
  wire _55685 = _55682 ^ _55684;
  wire _55686 = _3711 ^ _552;
  wire _55687 = _21690 ^ _55686;
  wire _55688 = _553 ^ _7736;
  wire _55689 = _55688 ^ _21701;
  wire _55690 = _55687 ^ _55689;
  wire _55691 = _55685 ^ _55690;
  wire _55692 = _55680 ^ _55691;
  wire _55693 = _18832 ^ _13866;
  wire _55694 = _5856 ^ _31201;
  wire _55695 = _55693 ^ _55694;
  wire _55696 = _40893 ^ _19806;
  wire _55697 = _55695 ^ _55696;
  wire _55698 = _17392 ^ _1411;
  wire _55699 = _27545 ^ _19815;
  wire _55700 = _55698 ^ _55699;
  wire _55701 = _25341 ^ _55700;
  wire _55702 = _55697 ^ _55701;
  wire _55703 = _40904 ^ _1427;
  wire _55704 = _42457 ^ _55703;
  wire _55705 = _7168 ^ _13357;
  wire _55706 = _30353 ^ _55705;
  wire _55707 = _55704 ^ _55706;
  wire _55708 = _5221 ^ _17910;
  wire _55709 = _43519 ^ _55708;
  wire _55710 = _2995 ^ _2232;
  wire _55711 = _5902 ^ _2238;
  wire _55712 = _55710 ^ _55711;
  wire _55713 = _55709 ^ _55712;
  wire _55714 = _55707 ^ _55713;
  wire _55715 = _55702 ^ _55714;
  wire _55716 = _55692 ^ _55715;
  wire _55717 = _1458 ^ _11746;
  wire _55718 = _1463 ^ _16924;
  wire _55719 = _55717 ^ _55718;
  wire _55720 = _40925 ^ _10646;
  wire _55721 = _38993 ^ _18870;
  wire _55722 = _55720 ^ _55721;
  wire _55723 = _55719 ^ _55722;
  wire _55724 = _3805 ^ _649;
  wire _55725 = _3808 ^ _5919;
  wire _55726 = _55724 ^ _55725;
  wire _55727 = _1489 ^ _1494;
  wire _55728 = _54869 ^ _55727;
  wire _55729 = _55726 ^ _55728;
  wire _55730 = _55723 ^ _55729;
  wire _55731 = _4551 ^ _5261;
  wire _55732 = _5266 ^ _10659;
  wire _55733 = _55731 ^ _55732;
  wire _55734 = _23581 ^ _12300;
  wire _55735 = _41730 ^ _55734;
  wire _55736 = _55733 ^ _55735;
  wire _55737 = _21762 ^ _1509;
  wire _55738 = _55737 ^ _54882;
  wire _55739 = _54501 ^ _12867;
  wire _55740 = uncoded_block[1398] ^ uncoded_block[1403];
  wire _55741 = _20340 ^ _55740;
  wire _55742 = _55739 ^ _55741;
  wire _55743 = _55738 ^ _55742;
  wire _55744 = _55736 ^ _55743;
  wire _55745 = _55730 ^ _55744;
  wire _55746 = uncoded_block[1415] ^ uncoded_block[1420];
  wire _55747 = _20347 ^ _55746;
  wire _55748 = _34197 ^ _55747;
  wire _55749 = _10683 ^ _14466;
  wire _55750 = _5968 ^ _4586;
  wire _55751 = _55749 ^ _55750;
  wire _55752 = _55748 ^ _55751;
  wire _55753 = _14978 ^ _4590;
  wire _55754 = _55753 ^ _6614;
  wire _55755 = _26763 ^ _20852;
  wire _55756 = _8452 ^ _3094;
  wire _55757 = _55755 ^ _55756;
  wire _55758 = _55754 ^ _55757;
  wire _55759 = _55752 ^ _55758;
  wire _55760 = uncoded_block[1467] ^ uncoded_block[1471];
  wire _55761 = _55760 ^ _3097;
  wire _55762 = _41757 ^ _17980;
  wire _55763 = _55761 ^ _55762;
  wire _55764 = _5329 ^ _2352;
  wire _55765 = _49097 ^ _6637;
  wire _55766 = _55764 ^ _55765;
  wire _55767 = _55763 ^ _55766;
  wire _55768 = _17494 ^ _54911;
  wire _55769 = _7269 ^ _2359;
  wire _55770 = _3123 ^ _6002;
  wire _55771 = _55769 ^ _55770;
  wire _55772 = _55768 ^ _55771;
  wire _55773 = _55767 ^ _55772;
  wire _55774 = _55759 ^ _55773;
  wire _55775 = _55745 ^ _55774;
  wire _55776 = _55716 ^ _55775;
  wire _55777 = _5347 ^ _3908;
  wire _55778 = _55777 ^ _36659;
  wire _55779 = _8482 ^ _767;
  wire _55780 = _55779 ^ _39833;
  wire _55781 = _55778 ^ _55780;
  wire _55782 = _28386 ^ _20392;
  wire _55783 = uncoded_block[1568] ^ uncoded_block[1574];
  wire _55784 = _55783 ^ _4648;
  wire _55785 = _55782 ^ _55784;
  wire _55786 = _6663 ^ _1609;
  wire _55787 = _15537 ^ _789;
  wire _55788 = _55786 ^ _55787;
  wire _55789 = _55785 ^ _55788;
  wire _55790 = _55781 ^ _55789;
  wire _55791 = _11847 ^ _6039;
  wire _55792 = _28396 ^ _55791;
  wire _55793 = _42166 ^ _12940;
  wire _55794 = _7297 ^ _7911;
  wire _55795 = _55793 ^ _55794;
  wire _55796 = _55792 ^ _55795;
  wire _55797 = _11308 ^ _28405;
  wire _55798 = _14530 ^ _820;
  wire _55799 = _18028 ^ _55798;
  wire _55800 = _55797 ^ _55799;
  wire _55801 = _55796 ^ _55800;
  wire _55802 = _55790 ^ _55801;
  wire _55803 = _2420 ^ _6059;
  wire _55804 = _4681 ^ _55803;
  wire _55805 = _832 ^ _9113;
  wire _55806 = _18982 ^ _24130;
  wire _55807 = _55805 ^ _55806;
  wire _55808 = _55804 ^ _55807;
  wire _55809 = _7331 ^ _6710;
  wire _55810 = _22772 ^ _20920;
  wire _55811 = _55809 ^ _55810;
  wire _55812 = uncoded_block[1705] ^ uncoded_block[1709];
  wire _55813 = uncoded_block[1711] ^ uncoded_block[1715];
  wire _55814 = _55812 ^ _55813;
  wire _55815 = _55814 ^ _39873;
  wire _55816 = _55811 ^ _55815;
  wire _55817 = _55808 ^ _55816;
  wire _55818 = _55802 ^ _55817;
  wire _55819 = _55776 ^ _55818;
  wire _55820 = _55670 ^ _55819;
  wire _55821 = uncoded_block[11] ^ uncoded_block[15];
  wire _55822 = _3212 ^ _55821;
  wire _55823 = _3211 ^ _55822;
  wire _55824 = _871 ^ _19963;
  wire _55825 = _4001 ^ _7959;
  wire _55826 = _55824 ^ _55825;
  wire _55827 = _55823 ^ _55826;
  wire _55828 = _9144 ^ _880;
  wire _55829 = _55828 ^ _18066;
  wire _55830 = _13548 ^ _25506;
  wire _55831 = _55829 ^ _55830;
  wire _55832 = _55827 ^ _55831;
  wire _55833 = _34 ^ _37127;
  wire _55834 = _55833 ^ _30932;
  wire _55835 = _9713 ^ _21429;
  wire _55836 = _9166 ^ _2491;
  wire _55837 = _55835 ^ _55836;
  wire _55838 = _55834 ^ _55837;
  wire _55839 = _9721 ^ _10821;
  wire _55840 = _52699 ^ _55839;
  wire _55841 = uncoded_block[125] ^ uncoded_block[131];
  wire _55842 = _55841 ^ _20963;
  wire _55843 = _8581 ^ _64;
  wire _55844 = _55842 ^ _55843;
  wire _55845 = _55840 ^ _55844;
  wire _55846 = _55838 ^ _55845;
  wire _55847 = _55832 ^ _55846;
  wire _55848 = _5469 ^ _14085;
  wire _55849 = _54606 ^ _55848;
  wire _55850 = _54610 ^ _82;
  wire _55851 = _53605 ^ _55850;
  wire _55852 = _55849 ^ _55851;
  wire _55853 = _85 ^ _18110;
  wire _55854 = _55853 ^ _44826;
  wire _55855 = _6798 ^ _3284;
  wire _55856 = uncoded_block[198] ^ uncoded_block[204];
  wire _55857 = _55856 ^ _6806;
  wire _55858 = _55855 ^ _55857;
  wire _55859 = _55854 ^ _55858;
  wire _55860 = _55852 ^ _55859;
  wire _55861 = uncoded_block[211] ^ uncoded_block[218];
  wire _55862 = _97 ^ _55861;
  wire _55863 = _35136 ^ _6168;
  wire _55864 = _55862 ^ _55863;
  wire _55865 = _45192 ^ _7424;
  wire _55866 = _55864 ^ _55865;
  wire _55867 = _5500 ^ _5503;
  wire _55868 = _55867 ^ _54626;
  wire _55869 = _39154 ^ _11419;
  wire _55870 = _55869 ^ _17132;
  wire _55871 = _55868 ^ _55870;
  wire _55872 = _55866 ^ _55871;
  wire _55873 = _55860 ^ _55872;
  wire _55874 = _55847 ^ _55873;
  wire _55875 = _119 ^ _25108;
  wire _55876 = uncoded_block[266] ^ uncoded_block[275];
  wire _55877 = _977 ^ _55876;
  wire _55878 = _55875 ^ _55877;
  wire _55879 = _53632 ^ _9773;
  wire _55880 = _55878 ^ _55879;
  wire _55881 = _10312 ^ _999;
  wire _55882 = _35546 ^ _55881;
  wire _55883 = _20536 ^ _145;
  wire _55884 = _55883 ^ _4831;
  wire _55885 = _55882 ^ _55884;
  wire _55886 = _55880 ^ _55885;
  wire _55887 = uncoded_block[320] ^ uncoded_block[326];
  wire _55888 = _55887 ^ _9782;
  wire _55889 = _55888 ^ _29669;
  wire _55890 = uncoded_block[343] ^ uncoded_block[348];
  wire _55891 = _55890 ^ _2599;
  wire _55892 = _55891 ^ _53650;
  wire _55893 = _55889 ^ _55892;
  wire _55894 = _30127 ^ _28836;
  wire _55895 = _28838 ^ _7476;
  wire _55896 = _55895 ^ _54662;
  wire _55897 = _55894 ^ _55896;
  wire _55898 = _55893 ^ _55897;
  wire _55899 = _55886 ^ _55898;
  wire _55900 = _23779 ^ _53657;
  wire _55901 = _4155 ^ _2625;
  wire _55902 = _55900 ^ _55901;
  wire _55903 = _6244 ^ _37205;
  wire _55904 = _9266 ^ _13112;
  wire _55905 = _55903 ^ _55904;
  wire _55906 = _55902 ^ _55905;
  wire _55907 = _53666 ^ _8097;
  wire _55908 = _25601 ^ _4174;
  wire _55909 = _6259 ^ _19621;
  wire _55910 = _55908 ^ _55909;
  wire _55911 = _55907 ^ _55910;
  wire _55912 = _55906 ^ _55911;
  wire _55913 = _1076 ^ _4181;
  wire _55914 = uncoded_block[463] ^ uncoded_block[469];
  wire _55915 = _55914 ^ _16692;
  wire _55916 = _55913 ^ _55915;
  wire _55917 = _1090 ^ _9832;
  wire _55918 = _3422 ^ _55917;
  wire _55919 = _55916 ^ _55918;
  wire _55920 = _27769 ^ _12033;
  wire _55921 = uncoded_block[502] ^ uncoded_block[505];
  wire _55922 = _55921 ^ _1892;
  wire _55923 = _55920 ^ _55922;
  wire _55924 = _10376 ^ _8705;
  wire _55925 = _55924 ^ _23371;
  wire _55926 = _55923 ^ _55925;
  wire _55927 = _55919 ^ _55926;
  wire _55928 = _55912 ^ _55927;
  wire _55929 = _55899 ^ _55928;
  wire _55930 = _55874 ^ _55929;
  wire _55931 = _1898 ^ _4921;
  wire _55932 = _55931 ^ _54695;
  wire _55933 = _20605 ^ _49739;
  wire _55934 = _55932 ^ _55933;
  wire _55935 = _5628 ^ _2687;
  wire _55936 = _52786 ^ _6940;
  wire _55937 = _55935 ^ _55936;
  wire _55938 = _7550 ^ _13698;
  wire _55939 = _9321 ^ _55938;
  wire _55940 = _55937 ^ _55939;
  wire _55941 = _55934 ^ _55940;
  wire _55942 = _1931 ^ _17718;
  wire _55943 = _270 ^ _9330;
  wire _55944 = _55942 ^ _55943;
  wire _55945 = _15247 ^ _2706;
  wire _55946 = _55945 ^ _34017;
  wire _55947 = _55944 ^ _55946;
  wire _55948 = _12609 ^ _13713;
  wire _55949 = _55948 ^ _25646;
  wire _55950 = _4964 ^ _7576;
  wire _55951 = _7577 ^ _11543;
  wire _55952 = _55950 ^ _55951;
  wire _55953 = _55949 ^ _55952;
  wire _55954 = _55947 ^ _55953;
  wire _55955 = _55941 ^ _55954;
  wire _55956 = _15766 ^ _10427;
  wire _55957 = _46666 ^ _55956;
  wire _55958 = _1963 ^ _311;
  wire _55959 = _3515 ^ _55958;
  wire _55960 = _55957 ^ _55959;
  wire _55961 = _40427 ^ _10434;
  wire _55962 = _55961 ^ _54727;
  wire _55963 = _31076 ^ _4272;
  wire _55964 = _55963 ^ _5682;
  wire _55965 = _55962 ^ _55964;
  wire _55966 = _55960 ^ _55965;
  wire _55967 = _45691 ^ _6364;
  wire _55968 = _8190 ^ _40044;
  wire _55969 = _55967 ^ _55968;
  wire _55970 = uncoded_block[721] ^ uncoded_block[726];
  wire _55971 = _55970 ^ _7603;
  wire _55972 = _13745 ^ _55971;
  wire _55973 = _55969 ^ _55972;
  wire _55974 = _53726 ^ _38868;
  wire _55975 = _5014 ^ _38457;
  wire _55976 = _55974 ^ _55975;
  wire _55977 = _55973 ^ _55976;
  wire _55978 = _55966 ^ _55977;
  wire _55979 = _55955 ^ _55978;
  wire _55980 = _8781 ^ _4301;
  wire _55981 = _54744 ^ _55980;
  wire _55982 = _3562 ^ _19217;
  wire _55983 = _16276 ^ _55982;
  wire _55984 = _55981 ^ _55983;
  wire _55985 = _2794 ^ _2018;
  wire _55986 = _55985 ^ _45327;
  wire _55987 = _54753 ^ _54757;
  wire _55988 = _55986 ^ _55987;
  wire _55989 = _55984 ^ _55988;
  wire _55990 = _31114 ^ _50903;
  wire _55991 = uncoded_block[823] ^ uncoded_block[828];
  wire _55992 = _55991 ^ _7039;
  wire _55993 = _45336 ^ _1257;
  wire _55994 = _55992 ^ _55993;
  wire _55995 = _55990 ^ _55994;
  wire _55996 = _14300 ^ _29800;
  wire _55997 = _6407 ^ _55996;
  wire _55998 = _31131 ^ _1272;
  wire _55999 = _54771 ^ _55998;
  wire _56000 = _55997 ^ _55999;
  wire _56001 = _55995 ^ _56000;
  wire _56002 = _55989 ^ _56001;
  wire _56003 = _9416 ^ _4355;
  wire _56004 = _37714 ^ _9960;
  wire _56005 = _56003 ^ _56004;
  wire _56006 = _3625 ^ _2852;
  wire _56007 = _433 ^ _56006;
  wire _56008 = _56005 ^ _56007;
  wire _56009 = _29379 ^ _55648;
  wire _56010 = _3633 ^ _56009;
  wire _56011 = _12725 ^ _4381;
  wire _56012 = _11077 ^ _56011;
  wire _56013 = _56010 ^ _56012;
  wire _56014 = _56008 ^ _56013;
  wire _56015 = _2091 ^ _16840;
  wire _56016 = _56015 ^ _54789;
  wire _56017 = _476 ^ _43844;
  wire _56018 = _56017 ^ _32017;
  wire _56019 = _2111 ^ _484;
  wire _56020 = _56019 ^ _5132;
  wire _56021 = _56018 ^ _56020;
  wire _56022 = _56016 ^ _56021;
  wire _56023 = _56014 ^ _56022;
  wire _56024 = _56002 ^ _56023;
  wire _56025 = _55979 ^ _56024;
  wire _56026 = _55930 ^ _56025;
  wire _56027 = _12750 ^ _8875;
  wire _56028 = _4417 ^ _2127;
  wire _56029 = _56027 ^ _56028;
  wire _56030 = _54806 ^ _29412;
  wire _56031 = _56029 ^ _56030;
  wire _56032 = _25768 ^ _521;
  wire _56033 = _56032 ^ _23502;
  wire _56034 = _8889 ^ _3691;
  wire _56035 = _56034 ^ _16871;
  wire _56036 = _56033 ^ _56035;
  wire _56037 = _56031 ^ _56036;
  wire _56038 = _3695 ^ _530;
  wire _56039 = _10575 ^ _3696;
  wire _56040 = _56038 ^ _56039;
  wire _56041 = _1374 ^ _536;
  wire _56042 = _537 ^ _5843;
  wire _56043 = _56041 ^ _56042;
  wire _56044 = _56040 ^ _56043;
  wire _56045 = _5169 ^ _53810;
  wire _56046 = _56045 ^ _2166;
  wire _56047 = _14375 ^ _15412;
  wire _56048 = _56046 ^ _56047;
  wire _56049 = _56044 ^ _56048;
  wire _56050 = _56037 ^ _56049;
  wire _56051 = _13866 ^ _6501;
  wire _56052 = _32462 ^ _56051;
  wire _56053 = _54832 ^ _4467;
  wire _56054 = _56052 ^ _56053;
  wire _56055 = _54834 ^ _54838;
  wire _56056 = _17390 ^ _11160;
  wire _56057 = _52928 ^ _3740;
  wire _56058 = _56056 ^ _56057;
  wire _56059 = _56055 ^ _56058;
  wire _56060 = _56054 ^ _56059;
  wire _56061 = _4488 ^ _22179;
  wire _56062 = _54842 ^ _56061;
  wire _56063 = _27549 ^ _7163;
  wire _56064 = _56063 ^ _23103;
  wire _56065 = _56062 ^ _56064;
  wire _56066 = _1433 ^ _1436;
  wire _56067 = _36984 ^ _56066;
  wire _56068 = _7169 ^ _2226;
  wire _56069 = _56068 ^ _20296;
  wire _56070 = _56067 ^ _56069;
  wire _56071 = _56065 ^ _56070;
  wire _56072 = _56060 ^ _56071;
  wire _56073 = _56050 ^ _56072;
  wire _56074 = _2235 ^ _24471;
  wire _56075 = _53843 ^ _56074;
  wire _56076 = _30361 ^ _7179;
  wire _56077 = uncoded_block[1275] ^ uncoded_block[1279];
  wire _56078 = _26718 ^ _56077;
  wire _56079 = _56076 ^ _56078;
  wire _56080 = _56075 ^ _56079;
  wire _56081 = _16924 ^ _642;
  wire _56082 = _56081 ^ _16928;
  wire _56083 = _10081 ^ _3807;
  wire _56084 = _1480 ^ _7197;
  wire _56085 = _56083 ^ _56084;
  wire _56086 = _56082 ^ _56085;
  wire _56087 = _56080 ^ _56086;
  wire _56088 = _1489 ^ _53861;
  wire _56089 = _6577 ^ _56088;
  wire _56090 = _10659 ^ _33363;
  wire _56091 = _29076 ^ _56090;
  wire _56092 = _56089 ^ _56091;
  wire _56093 = _12300 ^ _21762;
  wire _56094 = _42493 ^ _56093;
  wire _56095 = _1509 ^ _15966;
  wire _56096 = _3058 ^ _3061;
  wire _56097 = _56095 ^ _56096;
  wire _56098 = _56094 ^ _56097;
  wire _56099 = _56092 ^ _56098;
  wire _56100 = _56087 ^ _56099;
  wire _56101 = _12867 ^ _5952;
  wire _56102 = _56101 ^ _4573;
  wire _56103 = _12315 ^ _16954;
  wire _56104 = uncoded_block[1408] ^ uncoded_block[1413];
  wire _56105 = _56104 ^ _13422;
  wire _56106 = _56103 ^ _56105;
  wire _56107 = _56102 ^ _56106;
  wire _56108 = _11792 ^ _9022;
  wire _56109 = _2308 ^ _10684;
  wire _56110 = _56108 ^ _56109;
  wire _56111 = _23168 ^ _13432;
  wire _56112 = _56111 ^ _52620;
  wire _56113 = _56110 ^ _56112;
  wire _56114 = _56107 ^ _56113;
  wire _56115 = _26763 ^ _2326;
  wire _56116 = _2328 ^ _23174;
  wire _56117 = _56115 ^ _56116;
  wire _56118 = _2338 ^ _9608;
  wire _56119 = _13441 ^ _56118;
  wire _56120 = _56117 ^ _56119;
  wire _56121 = _4603 ^ _3884;
  wire _56122 = _56121 ^ _54901;
  wire _56123 = _56122 ^ _54909;
  wire _56124 = _56120 ^ _56123;
  wire _56125 = _56114 ^ _56124;
  wire _56126 = _56100 ^ _56125;
  wire _56127 = _56073 ^ _56126;
  wire _56128 = _7875 ^ _9055;
  wire _56129 = _5337 ^ _3898;
  wire _56130 = _56128 ^ _56129;
  wire _56131 = _5343 ^ _53901;
  wire _56132 = _22265 ^ _56131;
  wire _56133 = _56130 ^ _56132;
  wire _56134 = _4638 ^ _4640;
  wire _56135 = _5361 ^ _11284;
  wire _56136 = _56134 ^ _56135;
  wire _56137 = _54918 ^ _56136;
  wire _56138 = _56133 ^ _56137;
  wire _56139 = _7891 ^ _781;
  wire _56140 = _782 ^ _3924;
  wire _56141 = _56139 ^ _56140;
  wire _56142 = _2386 ^ _4653;
  wire _56143 = _56142 ^ _15036;
  wire _56144 = _56141 ^ _56143;
  wire _56145 = _801 ^ _6679;
  wire _56146 = _18505 ^ _56145;
  wire _56147 = _6680 ^ _3160;
  wire _56148 = _9656 ^ _5388;
  wire _56149 = _56147 ^ _56148;
  wire _56150 = _56146 ^ _56149;
  wire _56151 = _56144 ^ _56150;
  wire _56152 = _56138 ^ _56151;
  wire _56153 = _10755 ^ _2412;
  wire _56154 = _1643 ^ _56153;
  wire _56155 = _10757 ^ _820;
  wire _56156 = _56155 ^ _4681;
  wire _56157 = _56154 ^ _56156;
  wire _56158 = _22761 ^ _19939;
  wire _56159 = _30014 ^ _832;
  wire _56160 = _56158 ^ _56159;
  wire _56161 = _38681 ^ _49492;
  wire _56162 = _56160 ^ _56161;
  wire _56163 = _56157 ^ _56162;
  wire _56164 = _16060 ^ _5409;
  wire _56165 = _56164 ^ _54951;
  wire _56166 = _44408 ^ _7944;
  wire _56167 = _56166 ^ _7947;
  wire _56168 = _56165 ^ _56167;
  wire _56169 = _56163 ^ _56168;
  wire _56170 = _56152 ^ _56169;
  wire _56171 = _56127 ^ _56170;
  wire _56172 = _56026 ^ _56171;
  wire _56173 = _35096 ^ _49152;
  wire _56174 = _19501 ^ _21871;
  wire _56175 = _56173 ^ _56174;
  wire _56176 = _51482 ^ _56175;
  wire _56177 = _20457 ^ _19972;
  wire _56178 = _56177 ^ _49159;
  wire _56179 = _32 ^ _51804;
  wire _56180 = _56179 ^ _51488;
  wire _56181 = _56178 ^ _56180;
  wire _56182 = _56176 ^ _56181;
  wire _56183 = uncoded_block[88] ^ uncoded_block[94];
  wire _56184 = _56183 ^ _6758;
  wire _56185 = _31377 ^ _56184;
  wire _56186 = _56185 ^ _51495;
  wire _56187 = _46176 ^ _54970;
  wire _56188 = _52113 ^ _56187;
  wire _56189 = _56186 ^ _56188;
  wire _56190 = _56182 ^ _56189;
  wire _56191 = _53974 ^ _46185;
  wire _56192 = _52121 ^ _56191;
  wire _56193 = _46188 ^ _51826;
  wire _56194 = _104 ^ _20990;
  wire _56195 = _56194 ^ _11948;
  wire _56196 = _56193 ^ _56195;
  wire _56197 = _56192 ^ _56196;
  wire _56198 = _7423 ^ _10860;
  wire _56199 = _35145 ^ _39154;
  wire _56200 = _56198 ^ _56199;
  wire _56201 = _4095 ^ _26000;
  wire _56202 = _33934 ^ _56201;
  wire _56203 = _56200 ^ _56202;
  wire _56204 = _51838 ^ _46206;
  wire _56205 = _52128 ^ _56204;
  wire _56206 = _56203 ^ _56205;
  wire _56207 = _56197 ^ _56206;
  wire _56208 = _56190 ^ _56207;
  wire _56209 = _53995 ^ _53997;
  wire _56210 = _21029 ^ _51542;
  wire _56211 = _53998 ^ _56210;
  wire _56212 = _56209 ^ _56211;
  wire _56213 = _1838 ^ _48114;
  wire _56214 = _4858 ^ _10907;
  wire _56215 = _56213 ^ _56214;
  wire _56216 = _7487 ^ _1051;
  wire _56217 = _49230 ^ _56216;
  wire _56218 = _56215 ^ _56217;
  wire _56219 = _2629 ^ _51861;
  wire _56220 = _48870 ^ _14163;
  wire _56221 = _56219 ^ _56220;
  wire _56222 = _56221 ^ _52153;
  wire _56223 = _56218 ^ _56222;
  wire _56224 = _56212 ^ _56223;
  wire _56225 = _55213 ^ _51871;
  wire _56226 = _55218 ^ _51874;
  wire _56227 = _56225 ^ _56226;
  wire _56228 = _12577 ^ _27769;
  wire _56229 = _56228 ^ _52162;
  wire _56230 = _15220 ^ _4208;
  wire _56231 = _53421 ^ _56230;
  wire _56232 = _56229 ^ _56231;
  wire _56233 = _56227 ^ _56232;
  wire _56234 = _51884 ^ _48150;
  wire _56235 = _53138 ^ _55230;
  wire _56236 = _46261 ^ _46268;
  wire _56237 = _56235 ^ _56236;
  wire _56238 = _56234 ^ _56237;
  wire _56239 = _56233 ^ _56238;
  wire _56240 = _56224 ^ _56239;
  wire _56241 = _56208 ^ _56240;
  wire _56242 = _41939 ^ _42668;
  wire _56243 = _8148 ^ _4953;
  wire _56244 = _56243 ^ _47041;
  wire _56245 = _56242 ^ _56244;
  wire _56246 = _53157 ^ _50497;
  wire _56247 = _53440 ^ _56246;
  wire _56248 = _56245 ^ _56247;
  wire _56249 = _294 ^ _2729;
  wire _56250 = _56249 ^ _39633;
  wire _56251 = _3514 ^ _1173;
  wire _56252 = _36021 ^ _56251;
  wire _56253 = _56250 ^ _56252;
  wire _56254 = _1971 ^ _15281;
  wire _56255 = _17251 ^ _56254;
  wire _56256 = _1974 ^ _11556;
  wire _56257 = _56256 ^ _52477;
  wire _56258 = _56255 ^ _56257;
  wire _56259 = _56253 ^ _56258;
  wire _56260 = _56248 ^ _56259;
  wire _56261 = _25672 ^ _55025;
  wire _56262 = _55026 ^ _46302;
  wire _56263 = _56261 ^ _56262;
  wire _56264 = _353 ^ _1210;
  wire _56265 = _5017 ^ _5019;
  wire _56266 = _56264 ^ _56265;
  wire _56267 = _49307 ^ _7621;
  wire _56268 = _56266 ^ _56267;
  wire _56269 = _56263 ^ _56268;
  wire _56270 = _2019 ^ _12676;
  wire _56271 = _49310 ^ _56270;
  wire _56272 = _8223 ^ _7629;
  wire _56273 = _15814 ^ _51929;
  wire _56274 = _56272 ^ _56273;
  wire _56275 = _56271 ^ _56274;
  wire _56276 = _3587 ^ _27846;
  wire _56277 = _50903 ^ _56276;
  wire _56278 = _55279 ^ _55281;
  wire _56279 = _56277 ^ _56278;
  wire _56280 = _56275 ^ _56279;
  wire _56281 = _56269 ^ _56280;
  wire _56282 = _56260 ^ _56281;
  wire _56283 = _53468 ^ _55292;
  wire _56284 = _47103 ^ _9959;
  wire _56285 = _56284 ^ _55048;
  wire _56286 = _56283 ^ _56285;
  wire _56287 = _29379 ^ _7670;
  wire _56288 = _55049 ^ _56287;
  wire _56289 = _56288 ^ _51644;
  wire _56290 = _52528 ^ _16840;
  wire _56291 = uncoded_block[965] ^ uncoded_block[970];
  wire _56292 = _56291 ^ _468;
  wire _56293 = _56292 ^ _46351;
  wire _56294 = _56290 ^ _56293;
  wire _56295 = _56289 ^ _56294;
  wire _56296 = _56286 ^ _56295;
  wire _56297 = _24853 ^ _18333;
  wire _56298 = _10538 ^ _56297;
  wire _56299 = _56298 ^ _52539;
  wire _56300 = _8872 ^ _27496;
  wire _56301 = _26211 ^ _56300;
  wire _56302 = _3678 ^ _2910;
  wire _56303 = _56302 ^ _21681;
  wire _56304 = _56301 ^ _56303;
  wire _56305 = _56299 ^ _56304;
  wire _56306 = _8893 ^ _20251;
  wire _56307 = _56306 ^ _49010;
  wire _56308 = _49849 ^ _56307;
  wire _56309 = _18822 ^ _22612;
  wire _56310 = _19794 ^ _550;
  wire _56311 = _56310 ^ _55339;
  wire _56312 = _56309 ^ _56311;
  wire _56313 = _56308 ^ _56312;
  wire _56314 = _56305 ^ _56313;
  wire _56315 = _56296 ^ _56314;
  wire _56316 = _56282 ^ _56315;
  wire _56317 = _56241 ^ _56316;
  wire _56318 = _3718 ^ _33312;
  wire _56319 = _43121 ^ _27532;
  wire _56320 = _56318 ^ _56319;
  wire _56321 = _577 ^ _11711;
  wire _56322 = _56321 ^ _52268;
  wire _56323 = _56320 ^ _56322;
  wire _56324 = _52269 ^ _52000;
  wire _56325 = _49392 ^ _14909;
  wire _56326 = _56324 ^ _56325;
  wire _56327 = _56323 ^ _56326;
  wire _56328 = _4504 ^ _14919;
  wire _56329 = _55082 ^ _56328;
  wire _56330 = _55080 ^ _56329;
  wire _56331 = _52583 ^ _9528;
  wire _56332 = _1456 ^ _627;
  wire _56333 = _16413 ^ _56332;
  wire _56334 = _56331 ^ _56333;
  wire _56335 = _56330 ^ _56334;
  wire _56336 = _56327 ^ _56335;
  wire _56337 = _46419 ^ _29468;
  wire _56338 = _16924 ^ _24482;
  wire _56339 = _56337 ^ _56338;
  wire _56340 = _45826 ^ _4532;
  wire _56341 = _56340 ^ _48316;
  wire _56342 = _56339 ^ _56341;
  wire _56343 = _8407 ^ _21293;
  wire _56344 = _9555 ^ _19375;
  wire _56345 = _56343 ^ _56344;
  wire _56346 = _56345 ^ _53520;
  wire _56347 = _56342 ^ _56346;
  wire _56348 = _2283 ^ _55386;
  wire _56349 = _7824 ^ _6596;
  wire _56350 = _56348 ^ _56349;
  wire _56351 = _53521 ^ _56350;
  wire _56352 = _14968 ^ _3849;
  wire _56353 = _55098 ^ _56352;
  wire _56354 = _52040 ^ _56353;
  wire _56355 = _56351 ^ _56354;
  wire _56356 = _56347 ^ _56355;
  wire _56357 = _56336 ^ _56356;
  wire _56358 = _5968 ^ _21783;
  wire _56359 = _52044 ^ _56358;
  wire _56360 = _3857 ^ _13432;
  wire _56361 = _45085 ^ _9033;
  wire _56362 = _56360 ^ _56361;
  wire _56363 = _56359 ^ _56362;
  wire _56364 = _1550 ^ _23179;
  wire _56365 = _56364 ^ _51748;
  wire _56366 = _51745 ^ _56365;
  wire _56367 = _56363 ^ _56366;
  wire _56368 = _15996 ^ _3890;
  wire _56369 = _56368 ^ _28707;
  wire _56370 = _36227 ^ _51754;
  wire _56371 = _56369 ^ _56370;
  wire _56372 = _3900 ^ _9626;
  wire _56373 = _51757 ^ _56372;
  wire _56374 = _56373 ^ _46476;
  wire _56375 = _56371 ^ _56374;
  wire _56376 = _56367 ^ _56375;
  wire _56377 = _13988 ^ _16502;
  wire _56378 = _56377 ^ _53334;
  wire _56379 = _13478 ^ _3921;
  wire _56380 = _32567 ^ _3145;
  wire _56381 = _56379 ^ _56380;
  wire _56382 = _56381 ^ _46492;
  wire _56383 = _56378 ^ _56382;
  wire _56384 = _19929 ^ _12949;
  wire _56385 = _53555 ^ _56384;
  wire _56386 = _53553 ^ _56385;
  wire _56387 = _46506 ^ _17029;
  wire _56388 = _10761 ^ _1654;
  wire _56389 = _25024 ^ _56388;
  wire _56390 = _56387 ^ _56389;
  wire _56391 = _56386 ^ _56390;
  wire _56392 = _56383 ^ _56391;
  wire _56393 = _56376 ^ _56392;
  wire _56394 = _56357 ^ _56393;
  wire _56395 = _3186 ^ _19475;
  wire _56396 = _49985 ^ _56395;
  wire _56397 = _837 ^ _9675;
  wire _56398 = _56397 ^ _52667;
  wire _56399 = _56396 ^ _56398;
  wire _56400 = _52670 ^ uncoded_block[1721];
  wire _56401 = _56399 ^ _56400;
  wire _56402 = _56394 ^ _56401;
  wire _56403 = _56317 ^ _56402;
  wire _56404 = uncoded_block[0] ^ uncoded_block[9];
  wire _56405 = _56404 ^ _25498;
  wire _56406 = _1691 ^ _18;
  wire _56407 = _56405 ^ _56406;
  wire _56408 = uncoded_block[39] ^ uncoded_block[44];
  wire _56409 = uncoded_block[51] ^ uncoded_block[59];
  wire _56410 = _56408 ^ _56409;
  wire _56411 = uncoded_block[65] ^ uncoded_block[75];
  wire _56412 = uncoded_block[79] ^ uncoded_block[85];
  wire _56413 = _56411 ^ _56412;
  wire _56414 = _56410 ^ _56413;
  wire _56415 = _56407 ^ _56414;
  wire _56416 = uncoded_block[124] ^ uncoded_block[133];
  wire _56417 = _33056 ^ _56416;
  wire _56418 = _43642 ^ _56417;
  wire _56419 = uncoded_block[142] ^ uncoded_block[150];
  wire _56420 = _56419 ^ _1745;
  wire _56421 = _29623 ^ _54610;
  wire _56422 = _56420 ^ _56421;
  wire _56423 = _56418 ^ _56422;
  wire _56424 = _56415 ^ _56423;
  wire _56425 = _5477 ^ _41473;
  wire _56426 = uncoded_block[200] ^ uncoded_block[208];
  wire _56427 = _89 ^ _56426;
  wire _56428 = _56425 ^ _56427;
  wire _56429 = uncoded_block[212] ^ uncoded_block[219];
  wire _56430 = _56429 ^ _3299;
  wire _56431 = uncoded_block[232] ^ uncoded_block[249];
  wire _56432 = uncoded_block[251] ^ uncoded_block[259];
  wire _56433 = _56431 ^ _56432;
  wire _56434 = _56430 ^ _56433;
  wire _56435 = _56428 ^ _56434;
  wire _56436 = uncoded_block[267] ^ uncoded_block[273];
  wire _56437 = _53628 ^ _56436;
  wire _56438 = uncoded_block[274] ^ uncoded_block[280];
  wire _56439 = uncoded_block[287] ^ uncoded_block[292];
  wire _56440 = _56438 ^ _56439;
  wire _56441 = _56437 ^ _56440;
  wire _56442 = uncoded_block[316] ^ uncoded_block[324];
  wire _56443 = _995 ^ _56442;
  wire _56444 = uncoded_block[333] ^ uncoded_block[342];
  wire _56445 = _52740 ^ _56444;
  wire _56446 = _56443 ^ _56445;
  wire _56447 = _56441 ^ _56446;
  wire _56448 = _56435 ^ _56447;
  wire _56449 = _56424 ^ _56448;
  wire _56450 = uncoded_block[363] ^ uncoded_block[370];
  wire _56451 = _10329 ^ _56450;
  wire _56452 = uncoded_block[388] ^ uncoded_block[396];
  wire _56453 = _13101 ^ _56452;
  wire _56454 = _56451 ^ _56453;
  wire _56455 = uncoded_block[419] ^ uncoded_block[428];
  wire _56456 = _16177 ^ _56455;
  wire _56457 = uncoded_block[433] ^ uncoded_block[440];
  wire _56458 = _4167 ^ _56457;
  wire _56459 = _56456 ^ _56458;
  wire _56460 = _56454 ^ _56459;
  wire _56461 = uncoded_block[441] ^ uncoded_block[446];
  wire _56462 = uncoded_block[456] ^ uncoded_block[463];
  wire _56463 = _56461 ^ _56462;
  wire _56464 = uncoded_block[464] ^ uncoded_block[477];
  wire _56465 = _56464 ^ _42654;
  wire _56466 = _56463 ^ _56465;
  wire _56467 = _225 ^ _2667;
  wire _56468 = uncoded_block[530] ^ uncoded_block[536];
  wire _56469 = _25167 ^ _56468;
  wire _56470 = _56467 ^ _56469;
  wire _56471 = _56466 ^ _56470;
  wire _56472 = _56460 ^ _56471;
  wire _56473 = uncoded_block[543] ^ uncoded_block[553];
  wire _56474 = _24279 ^ _56473;
  wire _56475 = _1916 ^ _8139;
  wire _56476 = _56474 ^ _56475;
  wire _56477 = _52447 ^ _26096;
  wire _56478 = uncoded_block[595] ^ uncoded_block[602];
  wire _56479 = _20618 ^ _56478;
  wire _56480 = _56477 ^ _56479;
  wire _56481 = _56476 ^ _56480;
  wire _56482 = uncoded_block[616] ^ uncoded_block[624];
  wire _56483 = _14218 ^ _56482;
  wire _56484 = uncoded_block[627] ^ uncoded_block[631];
  wire _56485 = _56484 ^ _4249;
  wire _56486 = _56483 ^ _56485;
  wire _56487 = _4255 ^ _22954;
  wire _56488 = uncoded_block[649] ^ uncoded_block[655];
  wire _56489 = _56488 ^ _15270;
  wire _56490 = _56487 ^ _56489;
  wire _56491 = _56486 ^ _56490;
  wire _56492 = _56481 ^ _56491;
  wire _56493 = _56472 ^ _56492;
  wire _56494 = _56449 ^ _56493;
  wire _56495 = uncoded_block[669] ^ uncoded_block[689];
  wire _56496 = _56495 ^ _11556;
  wire _56497 = _22499 ^ _38450;
  wire _56498 = _56496 ^ _56497;
  wire _56499 = _2768 ^ _1206;
  wire _56500 = uncoded_block[741] ^ uncoded_block[747];
  wire _56501 = _56500 ^ _4293;
  wire _56502 = _56499 ^ _56501;
  wire _56503 = _56498 ^ _56502;
  wire _56504 = _12109 ^ _17776;
  wire _56505 = uncoded_block[771] ^ uncoded_block[779];
  wire _56506 = uncoded_block[784] ^ uncoded_block[793];
  wire _56507 = _56505 ^ _56506;
  wire _56508 = _56504 ^ _56507;
  wire _56509 = uncoded_block[801] ^ uncoded_block[811];
  wire _56510 = _56509 ^ _10486;
  wire _56511 = _56510 ^ _402;
  wire _56512 = _56508 ^ _56511;
  wire _56513 = _56503 ^ _56512;
  wire _56514 = uncoded_block[838] ^ uncoded_block[847];
  wire _56515 = uncoded_block[862] ^ uncoded_block[869];
  wire _56516 = _56514 ^ _56515;
  wire _56517 = uncoded_block[870] ^ uncoded_block[876];
  wire _56518 = uncoded_block[881] ^ uncoded_block[889];
  wire _56519 = _56517 ^ _56518;
  wire _56520 = _56516 ^ _56519;
  wire _56521 = uncoded_block[920] ^ uncoded_block[933];
  wire _56522 = _16312 ^ _56521;
  wire _56523 = _27049 ^ _56522;
  wire _56524 = _56520 ^ _56523;
  wire _56525 = uncoded_block[946] ^ uncoded_block[954];
  wire _56526 = _2083 ^ _56525;
  wire _56527 = uncoded_block[956] ^ uncoded_block[963];
  wire _56528 = uncoded_block[964] ^ uncoded_block[970];
  wire _56529 = _56527 ^ _56528;
  wire _56530 = _56526 ^ _56529;
  wire _56531 = _3657 ^ _32427;
  wire _56532 = uncoded_block[988] ^ uncoded_block[999];
  wire _56533 = _56532 ^ _1326;
  wire _56534 = _56531 ^ _56533;
  wire _56535 = _56530 ^ _56534;
  wire _56536 = _56524 ^ _56535;
  wire _56537 = _56513 ^ _56536;
  wire _56538 = _5129 ^ _6462;
  wire _56539 = uncoded_block[1020] ^ uncoded_block[1033];
  wire _56540 = uncoded_block[1034] ^ uncoded_block[1043];
  wire _56541 = _56539 ^ _56540;
  wire _56542 = _56538 ^ _56541;
  wire _56543 = uncoded_block[1051] ^ uncoded_block[1062];
  wire _56544 = _1356 ^ _56543;
  wire _56545 = uncoded_block[1068] ^ uncoded_block[1074];
  wire _56546 = _56545 ^ _2924;
  wire _56547 = _56544 ^ _56546;
  wire _56548 = _56542 ^ _56547;
  wire _56549 = uncoded_block[1090] ^ uncoded_block[1096];
  wire _56550 = _2925 ^ _56549;
  wire _56551 = _44259 ^ _34943;
  wire _56552 = _56550 ^ _56551;
  wire _56553 = uncoded_block[1108] ^ uncoded_block[1119];
  wire _56554 = _56553 ^ _2172;
  wire _56555 = uncoded_block[1136] ^ uncoded_block[1145];
  wire _56556 = _56555 ^ _5184;
  wire _56557 = _56554 ^ _56556;
  wire _56558 = _56552 ^ _56557;
  wire _56559 = _56548 ^ _56558;
  wire _56560 = _14894 ^ _22627;
  wire _56561 = _7151 ^ _10602;
  wire _56562 = _56560 ^ _56561;
  wire _56563 = uncoded_block[1176] ^ uncoded_block[1187];
  wire _56564 = _56563 ^ _5882;
  wire _56565 = _1425 ^ _36581;
  wire _56566 = _56564 ^ _56565;
  wire _56567 = _56562 ^ _56566;
  wire _56568 = uncoded_block[1224] ^ uncoded_block[1229];
  wire _56569 = uncoded_block[1231] ^ uncoded_block[1239];
  wire _56570 = _56568 ^ _56569;
  wire _56571 = _5228 ^ _7778;
  wire _56572 = _56570 ^ _56571;
  wire _56573 = uncoded_block[1257] ^ uncoded_block[1261];
  wire _56574 = uncoded_block[1263] ^ uncoded_block[1274];
  wire _56575 = _56573 ^ _56574;
  wire _56576 = _3011 ^ _3014;
  wire _56577 = _56575 ^ _56576;
  wire _56578 = _56572 ^ _56577;
  wire _56579 = _56567 ^ _56578;
  wire _56580 = _56559 ^ _56579;
  wire _56581 = _56537 ^ _56580;
  wire _56582 = _56494 ^ _56581;
  wire _56583 = _4532 ^ _4536;
  wire _56584 = uncoded_block[1312] ^ uncoded_block[1324];
  wire _56585 = uncoded_block[1330] ^ uncoded_block[1338];
  wire _56586 = _56584 ^ _56585;
  wire _56587 = _56583 ^ _56586;
  wire _56588 = uncoded_block[1341] ^ uncoded_block[1350];
  wire _56589 = _56588 ^ _5272;
  wire _56590 = uncoded_block[1360] ^ uncoded_block[1368];
  wire _56591 = _56590 ^ _3832;
  wire _56592 = _56589 ^ _56591;
  wire _56593 = _56587 ^ _56592;
  wire _56594 = uncoded_block[1377] ^ uncoded_block[1391];
  wire _56595 = _56594 ^ _2297;
  wire _56596 = uncoded_block[1406] ^ uncoded_block[1414];
  wire _56597 = _56596 ^ _5968;
  wire _56598 = _56595 ^ _56597;
  wire _56599 = uncoded_block[1439] ^ uncoded_block[1447];
  wire _56600 = _29508 ^ _56599;
  wire _56601 = _3865 ^ _2328;
  wire _56602 = _56600 ^ _56601;
  wire _56603 = _56598 ^ _56602;
  wire _56604 = _56593 ^ _56603;
  wire _56605 = _22252 ^ _4601;
  wire _56606 = _56605 ^ _22709;
  wire _56607 = _8461 ^ _1566;
  wire _56608 = _19421 ^ _13975;
  wire _56609 = _56607 ^ _56608;
  wire _56610 = _56606 ^ _56609;
  wire _56611 = _22723 ^ _1582;
  wire _56612 = _24994 ^ _5347;
  wire _56613 = _56611 ^ _56612;
  wire _56614 = uncoded_block[1566] ^ uncoded_block[1571];
  wire _56615 = _56614 ^ _18949;
  wire _56616 = _785 ^ _21827;
  wire _56617 = _56615 ^ _56616;
  wire _56618 = _56613 ^ _56617;
  wire _56619 = _56610 ^ _56618;
  wire _56620 = _56604 ^ _56619;
  wire _56621 = uncoded_block[1603] ^ uncoded_block[1612];
  wire _56622 = _29550 ^ _56621;
  wire _56623 = _47634 ^ _14006;
  wire _56624 = _56622 ^ _56623;
  wire _56625 = uncoded_block[1633] ^ uncoded_block[1643];
  wire _56626 = uncoded_block[1652] ^ uncoded_block[1663];
  wire _56627 = _56625 ^ _56626;
  wire _56628 = uncoded_block[1665] ^ uncoded_block[1679];
  wire _56629 = _56628 ^ _3967;
  wire _56630 = _56627 ^ _56629;
  wire _56631 = _56624 ^ _56630;
  wire _56632 = _1671 ^ uncoded_block[1714];
  wire _56633 = _56631 ^ _56632;
  wire _56634 = _56620 ^ _56633;
  wire _56635 = _56582 ^ _56634;
  wire _56636 = _4712 ^ _3995;
  wire _56637 = _4713 ^ _44790;
  wire _56638 = _56636 ^ _56637;
  wire _56639 = _3219 ^ _3224;
  wire _56640 = _11 ^ _10796;
  wire _56641 = _56639 ^ _56640;
  wire _56642 = _56638 ^ _56641;
  wire _56643 = _12425 ^ _34682;
  wire _56644 = _56643 ^ _19012;
  wire _56645 = _35 ^ _19511;
  wire _56646 = _56645 ^ _45160;
  wire _56647 = _56644 ^ _56646;
  wire _56648 = _56642 ^ _56647;
  wire _56649 = uncoded_block[85] ^ uncoded_block[90];
  wire _56650 = _11364 ^ _56649;
  wire _56651 = _6758 ^ _7377;
  wire _56652 = _56650 ^ _56651;
  wire _56653 = uncoded_block[104] ^ uncoded_block[108];
  wire _56654 = _56653 ^ _37537;
  wire _56655 = uncoded_block[114] ^ uncoded_block[121];
  wire _56656 = _56655 ^ _7386;
  wire _56657 = _56654 ^ _56656;
  wire _56658 = _56652 ^ _56657;
  wire _56659 = uncoded_block[142] ^ uncoded_block[149];
  wire _56660 = _4760 ^ _56659;
  wire _56661 = _36318 ^ _56660;
  wire _56662 = _41850 ^ _21906;
  wire _56663 = _28788 ^ _8591;
  wire _56664 = _56662 ^ _56663;
  wire _56665 = _56661 ^ _56664;
  wire _56666 = _56658 ^ _56665;
  wire _56667 = _56648 ^ _56666;
  wire _56668 = uncoded_block[179] ^ uncoded_block[186];
  wire _56669 = _938 ^ _56668;
  wire _56670 = _18111 ^ _5483;
  wire _56671 = _56669 ^ _56670;
  wire _56672 = _1763 ^ _6801;
  wire _56673 = _6158 ^ _21459;
  wire _56674 = _56672 ^ _56673;
  wire _56675 = _56671 ^ _56674;
  wire _56676 = uncoded_block[218] ^ uncoded_block[226];
  wire _56677 = _3296 ^ _56676;
  wire _56678 = _109 ^ _5500;
  wire _56679 = _56677 ^ _56678;
  wire _56680 = _2557 ^ _13055;
  wire _56681 = _35146 ^ _56680;
  wire _56682 = _56679 ^ _56681;
  wire _56683 = _56675 ^ _56682;
  wire _56684 = _4099 ^ _19566;
  wire _56685 = _20527 ^ _11967;
  wire _56686 = _56684 ^ _56685;
  wire _56687 = uncoded_block[288] ^ uncoded_block[293];
  wire _56688 = _19072 ^ _56687;
  wire _56689 = _21483 ^ _4824;
  wire _56690 = _56688 ^ _56689;
  wire _56691 = _56686 ^ _56690;
  wire _56692 = _4830 ^ _6209;
  wire _56693 = _45214 ^ _56692;
  wire _56694 = _1014 ^ _9240;
  wire _56695 = _56694 ^ _50070;
  wire _56696 = _56693 ^ _56695;
  wire _56697 = _56691 ^ _56696;
  wire _56698 = _56683 ^ _56697;
  wire _56699 = _56667 ^ _56698;
  wire _56700 = uncoded_block[347] ^ uncoded_block[353];
  wire _56701 = _4131 ^ _56700;
  wire _56702 = _1029 ^ _13093;
  wire _56703 = _56701 ^ _56702;
  wire _56704 = _21502 ^ _48117;
  wire _56705 = _29677 ^ _56704;
  wire _56706 = _56703 ^ _56705;
  wire _56707 = uncoded_block[406] ^ uncoded_block[413];
  wire _56708 = _5559 ^ _56707;
  wire _56709 = _41520 ^ _56708;
  wire _56710 = uncoded_block[421] ^ uncoded_block[424];
  wire _56711 = _56710 ^ _8672;
  wire _56712 = _34771 ^ _14690;
  wire _56713 = _56711 ^ _56712;
  wire _56714 = _56709 ^ _56713;
  wire _56715 = _56706 ^ _56714;
  wire _56716 = uncoded_block[454] ^ uncoded_block[463];
  wire _56717 = _208 ^ _56716;
  wire _56718 = _22431 ^ _56717;
  wire _56719 = _7507 ^ _21523;
  wire _56720 = _14176 ^ _16693;
  wire _56721 = _56719 ^ _56720;
  wire _56722 = _56718 ^ _56721;
  wire _56723 = _10934 ^ _7516;
  wire _56724 = _5603 ^ _21536;
  wire _56725 = _56723 ^ _56724;
  wire _56726 = uncoded_block[514] ^ uncoded_block[521];
  wire _56727 = _3439 ^ _56726;
  wire _56728 = _21538 ^ _56727;
  wire _56729 = _56725 ^ _56728;
  wire _56730 = _56722 ^ _56729;
  wire _56731 = _56715 ^ _56730;
  wire _56732 = uncoded_block[526] ^ uncoded_block[532];
  wire _56733 = _56732 ^ _40400;
  wire _56734 = _6298 ^ _24282;
  wire _56735 = _56733 ^ _56734;
  wire _56736 = uncoded_block[567] ^ uncoded_block[572];
  wire _56737 = _56736 ^ _10399;
  wire _56738 = _8726 ^ _56737;
  wire _56739 = _56735 ^ _56738;
  wire _56740 = uncoded_block[585] ^ uncoded_block[590];
  wire _56741 = _56740 ^ _2700;
  wire _56742 = _9860 ^ _56741;
  wire _56743 = _14737 ^ _14218;
  wire _56744 = _1942 ^ _17232;
  wire _56745 = _56743 ^ _56744;
  wire _56746 = _56742 ^ _56745;
  wire _56747 = _56739 ^ _56746;
  wire _56748 = _5652 ^ _7567;
  wire _56749 = uncoded_block[622] ^ uncoded_block[627];
  wire _56750 = _1946 ^ _56749;
  wire _56751 = _56748 ^ _56750;
  wire _56752 = _24760 ^ _22953;
  wire _56753 = _56751 ^ _56752;
  wire _56754 = uncoded_block[640] ^ uncoded_block[647];
  wire _56755 = uncoded_block[648] ^ uncoded_block[663];
  wire _56756 = _56754 ^ _56755;
  wire _56757 = _51249 ^ _17745;
  wire _56758 = _56756 ^ _56757;
  wire _56759 = uncoded_block[676] ^ uncoded_block[685];
  wire _56760 = _56759 ^ _11556;
  wire _56761 = _6990 ^ _4989;
  wire _56762 = _56760 ^ _56761;
  wire _56763 = _56758 ^ _56762;
  wire _56764 = _56753 ^ _56763;
  wire _56765 = _56747 ^ _56764;
  wire _56766 = _56731 ^ _56765;
  wire _56767 = _56699 ^ _56766;
  wire _56768 = _6992 ^ _6364;
  wire _56769 = _1192 ^ _10452;
  wire _56770 = _56768 ^ _56769;
  wire _56771 = uncoded_block[715] ^ uncoded_block[720];
  wire _56772 = _56771 ^ _4283;
  wire _56773 = _50518 ^ _7605;
  wire _56774 = _56772 ^ _56773;
  wire _56775 = _56770 ^ _56774;
  wire _56776 = _4289 ^ _5704;
  wire _56777 = _21605 ^ _1215;
  wire _56778 = _56776 ^ _56777;
  wire _56779 = _3559 ^ _2783;
  wire _56780 = uncoded_block[773] ^ uncoded_block[779];
  wire _56781 = _17776 ^ _56780;
  wire _56782 = _56779 ^ _56781;
  wire _56783 = _56778 ^ _56782;
  wire _56784 = _56775 ^ _56783;
  wire _56785 = _2018 ^ _12675;
  wire _56786 = _21614 ^ _386;
  wire _56787 = _56785 ^ _56786;
  wire _56788 = uncoded_block[808] ^ uncoded_block[814];
  wire _56789 = _12127 ^ _56788;
  wire _56790 = _5046 ^ _1242;
  wire _56791 = _56789 ^ _56790;
  wire _56792 = _56787 ^ _56791;
  wire _56793 = uncoded_block[824] ^ uncoded_block[832];
  wire _56794 = _56793 ^ _5057;
  wire _56795 = _11046 ^ _12141;
  wire _56796 = _56794 ^ _56795;
  wire _56797 = _8237 ^ _5066;
  wire _56798 = _4344 ^ _2828;
  wire _56799 = _56797 ^ _56798;
  wire _56800 = _56796 ^ _56799;
  wire _56801 = _56792 ^ _56800;
  wire _56802 = _56784 ^ _56801;
  wire _56803 = uncoded_block[872] ^ uncoded_block[877];
  wire _56804 = _6415 ^ _56803;
  wire _56805 = _29803 ^ _1272;
  wire _56806 = _56804 ^ _56805;
  wire _56807 = uncoded_block[892] ^ uncoded_block[897];
  wire _56808 = _15342 ^ _56807;
  wire _56809 = _56808 ^ _48610;
  wire _56810 = _56806 ^ _56809;
  wire _56811 = _432 ^ _7665;
  wire _56812 = _56811 ^ _48613;
  wire _56813 = _4368 ^ _1296;
  wire _56814 = _53771 ^ _2863;
  wire _56815 = _56813 ^ _56814;
  wire _56816 = _56812 ^ _56815;
  wire _56817 = _56810 ^ _56816;
  wire _56818 = uncoded_block[956] ^ uncoded_block[960];
  wire _56819 = _56818 ^ _12180;
  wire _56820 = _40098 ^ _56819;
  wire _56821 = _22113 ^ _5114;
  wire _56822 = uncoded_block[990] ^ uncoded_block[1001];
  wire _56823 = _11094 ^ _56822;
  wire _56824 = _56821 ^ _56823;
  wire _56825 = _56820 ^ _56824;
  wire _56826 = _4404 ^ _48991;
  wire _56827 = _492 ^ _495;
  wire _56828 = _56826 ^ _56827;
  wire _56829 = _6474 ^ _11677;
  wire _56830 = _7714 ^ _9465;
  wire _56831 = _56829 ^ _56830;
  wire _56832 = _56828 ^ _56831;
  wire _56833 = _56825 ^ _56832;
  wire _56834 = _56817 ^ _56833;
  wire _56835 = _56802 ^ _56834;
  wire _56836 = _10013 ^ _8889;
  wire _56837 = _5156 ^ _20251;
  wire _56838 = _56836 ^ _56837;
  wire _56839 = _534 ^ _13857;
  wire _56840 = _537 ^ _3704;
  wire _56841 = _56839 ^ _56840;
  wire _56842 = _56838 ^ _56841;
  wire _56843 = _15405 ^ _32042;
  wire _56844 = uncoded_block[1111] ^ uncoded_block[1117];
  wire _56845 = uncoded_block[1120] ^ uncoded_block[1127];
  wire _56846 = _56844 ^ _56845;
  wire _56847 = _56843 ^ _56846;
  wire _56848 = _8343 ^ _10593;
  wire _56849 = _20269 ^ _5862;
  wire _56850 = _56848 ^ _56849;
  wire _56851 = _56847 ^ _56850;
  wire _56852 = _56842 ^ _56851;
  wire _56853 = _2956 ^ _29439;
  wire _56854 = _3733 ^ _7749;
  wire _56855 = _56853 ^ _56854;
  wire _56856 = _2965 ^ _2195;
  wire _56857 = _44670 ^ _3749;
  wire _56858 = _56856 ^ _56857;
  wire _56859 = _56855 ^ _56858;
  wire _56860 = _51369 ^ _18389;
  wire _56861 = _1425 ^ _12813;
  wire _56862 = _56860 ^ _56861;
  wire _56863 = uncoded_block[1222] ^ uncoded_block[1227];
  wire _56864 = _15921 ^ _56863;
  wire _56865 = _56864 ^ _10066;
  wire _56866 = _56862 ^ _56865;
  wire _56867 = _56859 ^ _56866;
  wire _56868 = _56852 ^ _56867;
  wire _56869 = _3772 ^ _31231;
  wire _56870 = _6543 ^ _5231;
  wire _56871 = _56869 ^ _56870;
  wire _56872 = uncoded_block[1255] ^ uncoded_block[1260];
  wire _56873 = _56872 ^ _7178;
  wire _56874 = _9532 ^ _10075;
  wire _56875 = _56873 ^ _56874;
  wire _56876 = _56871 ^ _56875;
  wire _56877 = _7792 ^ _6560;
  wire _56878 = _24482 ^ _9545;
  wire _56879 = _56877 ^ _56878;
  wire _56880 = _35380 ^ _20812;
  wire _56881 = _56880 ^ _22212;
  wire _56882 = _56879 ^ _56881;
  wire _56883 = _56876 ^ _56882;
  wire _56884 = uncoded_block[1313] ^ uncoded_block[1320];
  wire _56885 = _56884 ^ _3029;
  wire _56886 = _36604 ^ _21753;
  wire _56887 = _56885 ^ _56886;
  wire _56888 = uncoded_block[1345] ^ uncoded_block[1355];
  wire _56889 = _5266 ^ _56888;
  wire _56890 = _56889 ^ _37823;
  wire _56891 = _56887 ^ _56890;
  wire _56892 = _10103 ^ _2290;
  wire _56893 = uncoded_block[1380] ^ uncoded_block[1386];
  wire _56894 = uncoded_block[1387] ^ uncoded_block[1393];
  wire _56895 = _56893 ^ _56894;
  wire _56896 = _56892 ^ _56895;
  wire _56897 = uncoded_block[1397] ^ uncoded_block[1404];
  wire _56898 = _56897 ^ _16954;
  wire _56899 = _56898 ^ _13948;
  wire _56900 = _56896 ^ _56899;
  wire _56901 = _56891 ^ _56900;
  wire _56902 = _56883 ^ _56901;
  wire _56903 = _56868 ^ _56902;
  wire _56904 = _56835 ^ _56903;
  wire _56905 = _56767 ^ _56904;
  wire _56906 = uncoded_block[1425] ^ uncoded_block[1430];
  wire _56907 = _17960 ^ _56906;
  wire _56908 = _56907 ^ _40216;
  wire _56909 = _712 ^ _6613;
  wire _56910 = _2322 ^ _1543;
  wire _56911 = _56909 ^ _56910;
  wire _56912 = _56908 ^ _56911;
  wire _56913 = _721 ^ _38629;
  wire _56914 = uncoded_block[1480] ^ uncoded_block[1486];
  wire _56915 = _56914 ^ _740;
  wire _56916 = _43952 ^ _56915;
  wire _56917 = _56913 ^ _56916;
  wire _56918 = _56912 ^ _56917;
  wire _56919 = _8462 ^ _6634;
  wire _56920 = _56919 ^ _33398;
  wire _56921 = uncoded_block[1524] ^ uncoded_block[1531];
  wire _56922 = uncoded_block[1532] ^ uncoded_block[1541];
  wire _56923 = _56921 ^ _56922;
  wire _56924 = _28371 ^ _56923;
  wire _56925 = _56920 ^ _56924;
  wire _56926 = _1590 ^ _8482;
  wire _56927 = _15020 ^ _9070;
  wire _56928 = _56926 ^ _56927;
  wire _56929 = uncoded_block[1560] ^ uncoded_block[1565];
  wire _56930 = _3914 ^ _56929;
  wire _56931 = _7891 ^ _9080;
  wire _56932 = _56930 ^ _56931;
  wire _56933 = _56928 ^ _56932;
  wire _56934 = _56925 ^ _56933;
  wire _56935 = _56918 ^ _56934;
  wire _56936 = uncoded_block[1576] ^ uncoded_block[1580];
  wire _56937 = _56936 ^ _15537;
  wire _56938 = uncoded_block[1587] ^ uncoded_block[1592];
  wire _56939 = _56938 ^ _29550;
  wire _56940 = _56937 ^ _56939;
  wire _56941 = _11847 ^ _1625;
  wire _56942 = _56941 ^ _48757;
  wire _56943 = _56940 ^ _56942;
  wire _56944 = _37082 ^ _40640;
  wire _56945 = _813 ^ _7309;
  wire _56946 = _56945 ^ _47261;
  wire _56947 = _56944 ^ _56946;
  wire _56948 = _56943 ^ _56947;
  wire _56949 = _13508 ^ _1654;
  wire _56950 = _56949 ^ _52663;
  wire _56951 = _2426 ^ _18982;
  wire _56952 = _11325 ^ _25037;
  wire _56953 = _56951 ^ _56952;
  wire _56954 = _56950 ^ _56953;
  wire _56955 = _852 ^ _855;
  wire _56956 = _9680 ^ _56955;
  wire _56957 = _56956 ^ uncoded_block[1720];
  wire _56958 = _56954 ^ _56957;
  wire _56959 = _56948 ^ _56958;
  wire _56960 = _56935 ^ _56959;
  wire _56961 = _56905 ^ _56960;
  wire _56962 = _4710 ^ _14560;
  wire _56963 = uncoded_block[19] ^ uncoded_block[26];
  wire _56964 = _56963 ^ _1693;
  wire _56965 = _56962 ^ _56964;
  wire _56966 = uncoded_block[34] ^ uncoded_block[40];
  wire _56967 = _56966 ^ _20457;
  wire _56968 = _13552 ^ _23698;
  wire _56969 = _56967 ^ _56968;
  wire _56970 = _56965 ^ _56969;
  wire _56971 = _5440 ^ _21881;
  wire _56972 = _30051 ^ _17578;
  wire _56973 = _56971 ^ _56972;
  wire _56974 = _14068 ^ _17583;
  wire _56975 = uncoded_block[106] ^ uncoded_block[113];
  wire _56976 = _56975 ^ _6769;
  wire _56977 = _56974 ^ _56976;
  wire _56978 = _56973 ^ _56977;
  wire _56979 = _56970 ^ _56978;
  wire _56980 = _4042 ^ _23720;
  wire _56981 = _1731 ^ _56980;
  wire _56982 = uncoded_block[149] ^ uncoded_block[153];
  wire _56983 = _4761 ^ _56982;
  wire _56984 = _10834 ^ _39128;
  wire _56985 = _56983 ^ _56984;
  wire _56986 = _56981 ^ _56985;
  wire _56987 = uncoded_block[173] ^ uncoded_block[179];
  wire _56988 = uncoded_block[180] ^ uncoded_block[185];
  wire _56989 = _56987 ^ _56988;
  wire _56990 = _46183 ^ _56989;
  wire _56991 = _49666 ^ _11402;
  wire _56992 = _10849 ^ _4779;
  wire _56993 = _56991 ^ _56992;
  wire _56994 = _56990 ^ _56993;
  wire _56995 = _56986 ^ _56994;
  wire _56996 = _56979 ^ _56995;
  wire _56997 = uncoded_block[209] ^ uncoded_block[216];
  wire _56998 = _56997 ^ _104;
  wire _56999 = uncoded_block[224] ^ uncoded_block[231];
  wire _57000 = _56999 ^ _25104;
  wire _57001 = _56998 ^ _57000;
  wire _57002 = uncoded_block[243] ^ uncoded_block[249];
  wire _57003 = _57002 ^ _7434;
  wire _57004 = uncoded_block[259] ^ uncoded_block[267];
  wire _57005 = _23746 ^ _57004;
  wire _57006 = _57003 ^ _57005;
  wire _57007 = _57001 ^ _57006;
  wire _57008 = _3320 ^ _26895;
  wire _57009 = _57008 ^ _39546;
  wire _57010 = _5522 ^ _24216;
  wire _57011 = _4824 ^ _12515;
  wire _57012 = _57010 ^ _57011;
  wire _57013 = _57009 ^ _57012;
  wire _57014 = _57007 ^ _57013;
  wire _57015 = _13619 ^ _11439;
  wire _57016 = uncoded_block[318] ^ uncoded_block[325];
  wire _57017 = uncoded_block[326] ^ uncoded_block[333];
  wire _57018 = _57016 ^ _57017;
  wire _57019 = _57015 ^ _57018;
  wire _57020 = _11987 ^ _29670;
  wire _57021 = _6221 ^ _13093;
  wire _57022 = _57020 ^ _57021;
  wire _57023 = _57019 ^ _57022;
  wire _57024 = _4853 ^ _10899;
  wire _57025 = _39961 ^ _2615;
  wire _57026 = _57024 ^ _57025;
  wire _57027 = _1847 ^ _49229;
  wire _57028 = _57027 ^ _56216;
  wire _57029 = _57026 ^ _57028;
  wire _57030 = _57023 ^ _57029;
  wire _57031 = _57014 ^ _57030;
  wire _57032 = _56996 ^ _57031;
  wire _57033 = _191 ^ _11476;
  wire _57034 = _11479 ^ _21974;
  wire _57035 = _57033 ^ _57034;
  wire _57036 = uncoded_block[447] ^ uncoded_block[464];
  wire _57037 = _9275 ^ _57036;
  wire _57038 = _9283 ^ _6266;
  wire _57039 = _57037 ^ _57038;
  wire _57040 = _57035 ^ _57039;
  wire _57041 = _49246 ^ _16200;
  wire _57042 = uncoded_block[496] ^ uncoded_block[505];
  wire _57043 = _10937 ^ _57042;
  wire _57044 = _57041 ^ _57043;
  wire _57045 = uncoded_block[512] ^ uncoded_block[519];
  wire _57046 = _3437 ^ _57045;
  wire _57047 = _1110 ^ _15230;
  wire _57048 = _57046 ^ _57047;
  wire _57049 = _57044 ^ _57048;
  wire _57050 = _57040 ^ _57049;
  wire _57051 = uncoded_block[544] ^ uncoded_block[552];
  wire _57052 = _14719 ^ _57051;
  wire _57053 = _8721 ^ _8724;
  wire _57054 = _57052 ^ _57053;
  wire _57055 = _1916 ^ _17218;
  wire _57056 = _13697 ^ _263;
  wire _57057 = _57055 ^ _57056;
  wire _57058 = _57054 ^ _57057;
  wire _57059 = uncoded_block[581] ^ uncoded_block[590];
  wire _57060 = _57059 ^ _8148;
  wire _57061 = _8738 ^ _277;
  wire _57062 = _57060 ^ _57061;
  wire _57063 = _14743 ^ _287;
  wire _57064 = _41947 ^ _57063;
  wire _57065 = _57062 ^ _57064;
  wire _57066 = _57058 ^ _57065;
  wire _57067 = _57050 ^ _57066;
  wire _57068 = _7576 ^ _13717;
  wire _57069 = _10424 ^ _297;
  wire _57070 = _57068 ^ _57069;
  wire _57071 = uncoded_block[653] ^ uncoded_block[660];
  wire _57072 = _57071 ^ _2742;
  wire _57073 = _38439 ^ _3519;
  wire _57074 = _57072 ^ _57073;
  wire _57075 = _57070 ^ _57074;
  wire _57076 = _22963 ^ _18249;
  wire _57077 = uncoded_block[697] ^ uncoded_block[707];
  wire _57078 = _1186 ^ _57077;
  wire _57079 = _57076 ^ _57078;
  wire _57080 = _10453 ^ _44172;
  wire _57081 = _57079 ^ _57080;
  wire _57082 = _57075 ^ _57081;
  wire _57083 = uncoded_block[726] ^ uncoded_block[735];
  wire _57084 = _57083 ^ _9908;
  wire _57085 = _57084 ^ _32368;
  wire _57086 = _21139 ^ _2005;
  wire _57087 = _11018 ^ _30659;
  wire _57088 = _57086 ^ _57087;
  wire _57089 = _57085 ^ _57088;
  wire _57090 = uncoded_block[773] ^ uncoded_block[778];
  wire _57091 = _57090 ^ _13219;
  wire _57092 = uncoded_block[783] ^ uncoded_block[790];
  wire _57093 = _57092 ^ _14797;
  wire _57094 = _57091 ^ _57093;
  wire _57095 = _31551 ^ _392;
  wire _57096 = _5729 ^ _2028;
  wire _57097 = _57095 ^ _57096;
  wire _57098 = _57094 ^ _57097;
  wire _57099 = _57089 ^ _57098;
  wire _57100 = _57082 ^ _57099;
  wire _57101 = _57067 ^ _57100;
  wire _57102 = _57032 ^ _57101;
  wire _57103 = _4331 ^ _7640;
  wire _57104 = _57103 ^ _37309;
  wire _57105 = uncoded_block[854] ^ uncoded_block[858];
  wire _57106 = _14814 ^ _57105;
  wire _57107 = _25253 ^ _2828;
  wire _57108 = _57106 ^ _57107;
  wire _57109 = _57104 ^ _57108;
  wire _57110 = uncoded_block[876] ^ uncoded_block[884];
  wire _57111 = _12696 ^ _57110;
  wire _57112 = _3613 ^ _8250;
  wire _57113 = _57111 ^ _57112;
  wire _57114 = _19249 ^ _53203;
  wire _57115 = _57113 ^ _57114;
  wire _57116 = _57109 ^ _57115;
  wire _57117 = _438 ^ _4368;
  wire _57118 = _44213 ^ _57117;
  wire _57119 = _2857 ^ _4375;
  wire _57120 = uncoded_block[949] ^ uncoded_block[955];
  wire _57121 = _57120 ^ _7086;
  wire _57122 = _57119 ^ _57121;
  wire _57123 = _57118 ^ _57122;
  wire _57124 = _2092 ^ _7088;
  wire _57125 = _57124 ^ _44987;
  wire _57126 = uncoded_block[976] ^ uncoded_block[984];
  wire _57127 = _57126 ^ _5118;
  wire _57128 = uncoded_block[994] ^ uncoded_block[1003];
  wire _57129 = _23939 ^ _57128;
  wire _57130 = _57127 ^ _57129;
  wire _57131 = _57125 ^ _57130;
  wire _57132 = _57123 ^ _57131;
  wire _57133 = _57116 ^ _57132;
  wire _57134 = _24400 ^ _2890;
  wire _57135 = uncoded_block[1025] ^ uncoded_block[1033];
  wire _57136 = _55315 ^ _57135;
  wire _57137 = _57134 ^ _57136;
  wire _57138 = uncoded_block[1043] ^ uncoded_block[1050];
  wire _57139 = _57138 ^ _4430;
  wire _57140 = _12764 ^ _7717;
  wire _57141 = _57139 ^ _57140;
  wire _57142 = _57137 ^ _57141;
  wire _57143 = uncoded_block[1065] ^ uncoded_block[1074];
  wire _57144 = _57143 ^ _6486;
  wire _57145 = _11126 ^ _20753;
  wire _57146 = _57144 ^ _57145;
  wire _57147 = uncoded_block[1115] ^ uncoded_block[1120];
  wire _57148 = _15405 ^ _57147;
  wire _57149 = _4443 ^ _57148;
  wire _57150 = _57146 ^ _57149;
  wire _57151 = _57142 ^ _57150;
  wire _57152 = uncoded_block[1122] ^ uncoded_block[1127];
  wire _57153 = _57152 ^ _564;
  wire _57154 = _5184 ^ _4469;
  wire _57155 = _57153 ^ _57154;
  wire _57156 = _2188 ^ _13335;
  wire _57157 = _32064 ^ _589;
  wire _57158 = _57156 ^ _57157;
  wire _57159 = _57155 ^ _57158;
  wire _57160 = uncoded_block[1182] ^ uncoded_block[1191];
  wire _57161 = _10608 ^ _57160;
  wire _57162 = _11719 ^ _2206;
  wire _57163 = _57161 ^ _57162;
  wire _57164 = _2209 ^ _5885;
  wire _57165 = _57164 ^ _28643;
  wire _57166 = _57163 ^ _57165;
  wire _57167 = _57159 ^ _57166;
  wire _57168 = _57151 ^ _57167;
  wire _57169 = _57133 ^ _57168;
  wire _57170 = _27555 ^ _46798;
  wire _57171 = uncoded_block[1232] ^ uncoded_block[1244];
  wire _57172 = _57171 ^ _2232;
  wire _57173 = _11737 ^ _3784;
  wire _57174 = _57172 ^ _57173;
  wire _57175 = _57170 ^ _57174;
  wire _57176 = uncoded_block[1266] ^ uncoded_block[1274];
  wire _57177 = _3004 ^ _57176;
  wire _57178 = uncoded_block[1276] ^ uncoded_block[1281];
  wire _57179 = _57178 ^ _24482;
  wire _57180 = _57177 ^ _57179;
  wire _57181 = _45826 ^ _9547;
  wire _57182 = _46091 ^ _1482;
  wire _57183 = _57181 ^ _57182;
  wire _57184 = _57180 ^ _57183;
  wire _57185 = _57175 ^ _57184;
  wire _57186 = _4543 ^ _5932;
  wire _57187 = _32921 ^ _57186;
  wire _57188 = uncoded_block[1350] ^ uncoded_block[1358];
  wire _57189 = _29486 ^ _57188;
  wire _57190 = _57189 ^ _21763;
  wire _57191 = _57187 ^ _57190;
  wire _57192 = uncoded_block[1372] ^ uncoded_block[1378];
  wire _57193 = _57192 ^ _7219;
  wire _57194 = _6596 ^ _9578;
  wire _57195 = _57193 ^ _57194;
  wire _57196 = _5953 ^ _42502;
  wire _57197 = _57195 ^ _57196;
  wire _57198 = _57191 ^ _57197;
  wire _57199 = _57185 ^ _57198;
  wire _57200 = _29095 ^ _5968;
  wire _57201 = _13948 ^ _57200;
  wire _57202 = _17470 ^ _26763;
  wire _57203 = _1544 ^ _10136;
  wire _57204 = _57202 ^ _57203;
  wire _57205 = _57201 ^ _57204;
  wire _57206 = _49091 ^ _15994;
  wire _57207 = _54173 ^ _7864;
  wire _57208 = _57206 ^ _57207;
  wire _57209 = _38636 ^ _7262;
  wire _57210 = _57209 ^ _39049;
  wire _57211 = _57208 ^ _57210;
  wire _57212 = _57205 ^ _57211;
  wire _57213 = _5337 ^ _11270;
  wire _57214 = _57213 ^ _41770;
  wire _57215 = _19903 ^ _32975;
  wire _57216 = uncoded_block[1544] ^ uncoded_block[1549];
  wire _57217 = uncoded_block[1550] ^ uncoded_block[1554];
  wire _57218 = _57216 ^ _57217;
  wire _57219 = _57215 ^ _57218;
  wire _57220 = _57214 ^ _57219;
  wire _57221 = _1596 ^ _5361;
  wire _57222 = _57221 ^ _43221;
  wire _57223 = _3921 ^ _6671;
  wire _57224 = _15538 ^ _11292;
  wire _57225 = _57223 ^ _57224;
  wire _57226 = _57222 ^ _57225;
  wire _57227 = _57220 ^ _57226;
  wire _57228 = _57212 ^ _57227;
  wire _57229 = _57199 ^ _57228;
  wire _57230 = _57169 ^ _57229;
  wire _57231 = _57102 ^ _57230;
  wire _57232 = _51771 ^ _46494;
  wire _57233 = _6680 ^ _38668;
  wire _57234 = uncoded_block[1636] ^ uncoded_block[1644];
  wire _57235 = _1636 ^ _57234;
  wire _57236 = _57233 ^ _57235;
  wire _57237 = _57232 ^ _57236;
  wire _57238 = _9661 ^ _4677;
  wire _57239 = uncoded_block[1653] ^ uncoded_block[1664];
  wire _57240 = _57239 ^ _7319;
  wire _57241 = _57238 ^ _57240;
  wire _57242 = uncoded_block[1672] ^ uncoded_block[1681];
  wire _57243 = _2422 ^ _57242;
  wire _57244 = _33018 ^ _839;
  wire _57245 = _57243 ^ _57244;
  wire _57246 = _57241 ^ _57245;
  wire _57247 = _57237 ^ _57246;
  wire _57248 = _4698 ^ _15063;
  wire _57249 = _2437 ^ _854;
  wire _57250 = _57248 ^ _57249;
  wire _57251 = _57250 ^ _5416;
  wire _57252 = _57247 ^ _57251;
  wire _57253 = _57231 ^ _57252;
  wire _57254 = uncoded_block[10] ^ uncoded_block[16];
  wire _57255 = _24147 ^ _57254;
  wire _57256 = _57255 ^ _9695;
  wire _57257 = _879 ^ _20457;
  wire _57258 = _7966 ^ _3232;
  wire _57259 = _57257 ^ _57258;
  wire _57260 = _57256 ^ _57259;
  wire _57261 = _4014 ^ _15087;
  wire _57262 = _10801 ^ _32;
  wire _57263 = _57261 ^ _57262;
  wire _57264 = _6744 ^ _7367;
  wire _57265 = uncoded_block[74] ^ uncoded_block[78];
  wire _57266 = _57265 ^ _4735;
  wire _57267 = _57264 ^ _57266;
  wire _57268 = _57263 ^ _57267;
  wire _57269 = _57260 ^ _57268;
  wire _57270 = _41 ^ _4738;
  wire _57271 = uncoded_block[90] ^ uncoded_block[96];
  wire _57272 = _57271 ^ _9718;
  wire _57273 = _57270 ^ _57272;
  wire _57274 = _48810 ^ _5453;
  wire _57275 = uncoded_block[112] ^ uncoded_block[117];
  wire _57276 = _57275 ^ _2498;
  wire _57277 = _57274 ^ _57276;
  wire _57278 = _57273 ^ _57277;
  wire _57279 = _33058 ^ _6774;
  wire _57280 = _57279 ^ _31807;
  wire _57281 = _64 ^ _6780;
  wire _57282 = _74 ^ _4054;
  wire _57283 = _57281 ^ _57282;
  wire _57284 = _57280 ^ _57283;
  wire _57285 = _57278 ^ _57284;
  wire _57286 = _57269 ^ _57285;
  wire _57287 = _10271 ^ _39135;
  wire _57288 = _9196 ^ _33077;
  wire _57289 = _9745 ^ _10278;
  wire _57290 = _57288 ^ _57289;
  wire _57291 = _57287 ^ _57290;
  wire _57292 = uncoded_block[220] ^ uncoded_block[229];
  wire _57293 = _27295 ^ _57292;
  wire _57294 = _10281 ^ _57293;
  wire _57295 = _25104 ^ _57002;
  wire _57296 = _4800 ^ _3309;
  wire _57297 = _57295 ^ _57296;
  wire _57298 = _57294 ^ _57297;
  wire _57299 = _57291 ^ _57298;
  wire _57300 = _3311 ^ _7438;
  wire _57301 = _6831 ^ _7441;
  wire _57302 = _57300 ^ _57301;
  wire _57303 = _3321 ^ _7445;
  wire _57304 = _8632 ^ _4820;
  wire _57305 = _57303 ^ _57304;
  wire _57306 = _57302 ^ _57305;
  wire _57307 = _8051 ^ _4826;
  wire _57308 = _57307 ^ _55186;
  wire _57309 = _15671 ^ _2580;
  wire _57310 = _30117 ^ _9235;
  wire _57311 = _57309 ^ _57310;
  wire _57312 = _57308 ^ _57311;
  wire _57313 = _57306 ^ _57312;
  wire _57314 = _57299 ^ _57313;
  wire _57315 = _57286 ^ _57314;
  wire _57316 = _22873 ^ _7463;
  wire _57317 = _32687 ^ _161;
  wire _57318 = _57316 ^ _57317;
  wire _57319 = _23330 ^ _16662;
  wire _57320 = _27735 ^ _57319;
  wire _57321 = _57318 ^ _57320;
  wire _57322 = _1035 ^ _10895;
  wire _57323 = _14671 ^ _4858;
  wire _57324 = _57322 ^ _57323;
  wire _57325 = _12005 ^ _1847;
  wire _57326 = uncoded_block[403] ^ uncoded_block[411];
  wire _57327 = _10341 ^ _57326;
  wire _57328 = _57325 ^ _57327;
  wire _57329 = _57324 ^ _57328;
  wire _57330 = _57321 ^ _57329;
  wire _57331 = _13650 ^ _193;
  wire _57332 = uncoded_block[426] ^ uncoded_block[432];
  wire _57333 = _1059 ^ _57332;
  wire _57334 = _57331 ^ _57333;
  wire _57335 = _9271 ^ _6255;
  wire _57336 = _57335 ^ _50459;
  wire _57337 = _57334 ^ _57336;
  wire _57338 = _39197 ^ _213;
  wire _57339 = _35581 ^ _57338;
  wire _57340 = uncoded_block[460] ^ uncoded_block[468];
  wire _57341 = uncoded_block[469] ^ uncoded_block[473];
  wire _57342 = _57340 ^ _57341;
  wire _57343 = _4189 ^ _20588;
  wire _57344 = _57342 ^ _57343;
  wire _57345 = _57339 ^ _57344;
  wire _57346 = _57337 ^ _57345;
  wire _57347 = _57330 ^ _57346;
  wire _57348 = _49727 ^ _28870;
  wire _57349 = uncoded_block[503] ^ uncoded_block[517];
  wire _57350 = _57349 ^ _3444;
  wire _57351 = _237 ^ _13684;
  wire _57352 = _57350 ^ _57351;
  wire _57353 = _57348 ^ _57352;
  wire _57354 = uncoded_block[526] ^ uncoded_block[531];
  wire _57355 = _57354 ^ _4215;
  wire _57356 = _21079 ^ _25173;
  wire _57357 = _57355 ^ _57356;
  wire _57358 = _10959 ^ _2687;
  wire _57359 = _13159 ^ _12051;
  wire _57360 = _57358 ^ _57359;
  wire _57361 = _57357 ^ _57360;
  wire _57362 = _57353 ^ _57361;
  wire _57363 = _3467 ^ _39617;
  wire _57364 = _57363 ^ _22011;
  wire _57365 = uncoded_block[585] ^ uncoded_block[592];
  wire _57366 = _3475 ^ _57365;
  wire _57367 = uncoded_block[599] ^ uncoded_block[606];
  wire _57368 = _4236 ^ _57367;
  wire _57369 = _57366 ^ _57368;
  wire _57370 = _57364 ^ _57369;
  wire _57371 = _8739 ^ _7564;
  wire _57372 = _57371 ^ _14744;
  wire _57373 = _38046 ^ _10424;
  wire _57374 = _29319 ^ _57373;
  wire _57375 = _57372 ^ _57374;
  wire _57376 = _57370 ^ _57375;
  wire _57377 = _57362 ^ _57376;
  wire _57378 = _57347 ^ _57377;
  wire _57379 = _57315 ^ _57378;
  wire _57380 = _51592 ^ _46671;
  wire _57381 = _308 ^ _10990;
  wire _57382 = _10434 ^ _1968;
  wire _57383 = _57381 ^ _57382;
  wire _57384 = _57380 ^ _57383;
  wire _57385 = _1971 ^ _8180;
  wire _57386 = uncoded_block[690] ^ uncoded_block[695];
  wire _57387 = _322 ^ _57386;
  wire _57388 = _57385 ^ _57387;
  wire _57389 = _3529 ^ _34840;
  wire _57390 = _11565 ^ _2763;
  wire _57391 = _57389 ^ _57390;
  wire _57392 = _57388 ^ _57391;
  wire _57393 = _57384 ^ _57392;
  wire _57394 = uncoded_block[724] ^ uncoded_block[729];
  wire _57395 = _57394 ^ _8201;
  wire _57396 = uncoded_block[736] ^ uncoded_block[740];
  wire _57397 = _57396 ^ _28930;
  wire _57398 = _57395 ^ _57397;
  wire _57399 = _5017 ^ _7614;
  wire _57400 = _13215 ^ _34855;
  wire _57401 = _57399 ^ _57400;
  wire _57402 = _57398 ^ _57401;
  wire _57403 = _3567 ^ _12669;
  wire _57404 = _2015 ^ _43425;
  wire _57405 = _57403 ^ _57404;
  wire _57406 = uncoded_block[796] ^ uncoded_block[803];
  wire _57407 = _57406 ^ _34062;
  wire _57408 = uncoded_block[809] ^ uncoded_block[819];
  wire _57409 = uncoded_block[821] ^ uncoded_block[832];
  wire _57410 = _57408 ^ _57409;
  wire _57411 = _57407 ^ _57410;
  wire _57412 = _57405 ^ _57411;
  wire _57413 = _57402 ^ _57412;
  wire _57414 = _57393 ^ _57413;
  wire _57415 = _1250 ^ _1253;
  wire _57416 = _25710 ^ _2823;
  wire _57417 = _57415 ^ _57416;
  wire _57418 = uncoded_block[864] ^ uncoded_block[870];
  wire _57419 = _57418 ^ _416;
  wire _57420 = uncoded_block[884] ^ uncoded_block[894];
  wire _57421 = _4347 ^ _57420;
  wire _57422 = _57419 ^ _57421;
  wire _57423 = _57417 ^ _57422;
  wire _57424 = _5085 ^ _429;
  wire _57425 = _9960 ^ _2071;
  wire _57426 = _57424 ^ _57425;
  wire _57427 = _21182 ^ _39692;
  wire _57428 = _31995 ^ _18316;
  wire _57429 = _57427 ^ _57428;
  wire _57430 = _57426 ^ _57429;
  wire _57431 = _57423 ^ _57430;
  wire _57432 = _10517 ^ _2083;
  wire _57433 = _57432 ^ _10524;
  wire _57434 = _7680 ^ _10529;
  wire _57435 = _7682 ^ _25283;
  wire _57436 = _57434 ^ _57435;
  wire _57437 = _57433 ^ _57436;
  wire _57438 = uncoded_block[979] ^ uncoded_block[983];
  wire _57439 = _28233 ^ _57438;
  wire _57440 = _5118 ^ _23040;
  wire _57441 = _57439 ^ _57440;
  wire _57442 = _4410 ^ _11663;
  wire _57443 = _43849 ^ _57442;
  wire _57444 = _57441 ^ _57443;
  wire _57445 = _57437 ^ _57444;
  wire _57446 = _57431 ^ _57445;
  wire _57447 = _57414 ^ _57446;
  wire _57448 = _7108 ^ _18801;
  wire _57449 = _499 ^ _50575;
  wire _57450 = _57448 ^ _57449;
  wire _57451 = _6475 ^ _12208;
  wire _57452 = _1357 ^ _38944;
  wire _57453 = _57451 ^ _57452;
  wire _57454 = _57450 ^ _57453;
  wire _57455 = uncoded_block[1062] ^ uncoded_block[1066];
  wire _57456 = _57455 ^ _12213;
  wire _57457 = uncoded_block[1074] ^ uncoded_block[1081];
  wire _57458 = _527 ^ _57457;
  wire _57459 = _57456 ^ _57458;
  wire _57460 = uncoded_block[1086] ^ uncoded_block[1091];
  wire _57461 = _21687 ^ _57460;
  wire _57462 = _5166 ^ _7731;
  wire _57463 = _57461 ^ _57462;
  wire _57464 = _57459 ^ _57463;
  wire _57465 = _57454 ^ _57464;
  wire _57466 = _20761 ^ _14882;
  wire _57467 = _57466 ^ _16884;
  wire _57468 = _7736 ^ _5854;
  wire _57469 = _23523 ^ _8929;
  wire _57470 = _57468 ^ _57469;
  wire _57471 = _57467 ^ _57470;
  wire _57472 = _565 ^ _8932;
  wire _57473 = _29439 ^ _11157;
  wire _57474 = _57472 ^ _57473;
  wire _57475 = _581 ^ _1407;
  wire _57476 = uncoded_block[1169] ^ uncoded_block[1178];
  wire _57477 = _57476 ^ _10608;
  wire _57478 = _57475 ^ _57477;
  wire _57479 = _57474 ^ _57478;
  wire _57480 = _57471 ^ _57479;
  wire _57481 = _57465 ^ _57480;
  wire _57482 = _592 ^ _13883;
  wire _57483 = uncoded_block[1193] ^ uncoded_block[1197];
  wire _57484 = uncoded_block[1199] ^ uncoded_block[1206];
  wire _57485 = _57483 ^ _57484;
  wire _57486 = _57482 ^ _57485;
  wire _57487 = _2216 ^ _10617;
  wire _57488 = _12813 ^ _5215;
  wire _57489 = _57487 ^ _57488;
  wire _57490 = _57486 ^ _57489;
  wire _57491 = _6532 ^ _11177;
  wire _57492 = _8377 ^ _14919;
  wire _57493 = _57491 ^ _57492;
  wire _57494 = _43141 ^ _10067;
  wire _57495 = _57494 ^ _32081;
  wire _57496 = _57493 ^ _57495;
  wire _57497 = _57490 ^ _57496;
  wire _57498 = uncoded_block[1263] ^ uncoded_block[1270];
  wire _57499 = uncoded_block[1274] ^ uncoded_block[1278];
  wire _57500 = _57498 ^ _57499;
  wire _57501 = _55367 ^ _57500;
  wire _57502 = _639 ^ _8980;
  wire _57503 = _13911 ^ _57502;
  wire _57504 = _57501 ^ _57503;
  wire _57505 = _22662 ^ _3808;
  wire _57506 = uncoded_block[1313] ^ uncoded_block[1318];
  wire _57507 = _57506 ^ _37813;
  wire _57508 = _57505 ^ _57507;
  wire _57509 = _7201 ^ _11207;
  wire _57510 = _16437 ^ _1497;
  wire _57511 = _57509 ^ _57510;
  wire _57512 = _57508 ^ _57511;
  wire _57513 = _57504 ^ _57512;
  wire _57514 = _57497 ^ _57513;
  wire _57515 = _57481 ^ _57514;
  wire _57516 = _57447 ^ _57515;
  wire _57517 = _57379 ^ _57516;
  wire _57518 = uncoded_block[1349] ^ uncoded_block[1355];
  wire _57519 = _5268 ^ _57518;
  wire _57520 = _57519 ^ _26286;
  wire _57521 = _12302 ^ _680;
  wire _57522 = _7823 ^ _4564;
  wire _57523 = _57521 ^ _57522;
  wire _57524 = _57520 ^ _57523;
  wire _57525 = _6596 ^ _19864;
  wire _57526 = _57525 ^ _1518;
  wire _57527 = uncoded_block[1409] ^ uncoded_block[1414];
  wire _57528 = _16459 ^ _57527;
  wire _57529 = uncoded_block[1415] ^ uncoded_block[1423];
  wire _57530 = _57529 ^ _9590;
  wire _57531 = _57528 ^ _57530;
  wire _57532 = _57526 ^ _57531;
  wire _57533 = _57524 ^ _57532;
  wire _57534 = _8443 ^ _27175;
  wire _57535 = uncoded_block[1450] ^ uncoded_block[1456];
  wire _57536 = _3864 ^ _57535;
  wire _57537 = _57534 ^ _57536;
  wire _57538 = _4596 ^ _3871;
  wire _57539 = _57538 ^ _49941;
  wire _57540 = _57537 ^ _57539;
  wire _57541 = _5320 ^ _49947;
  wire _57542 = _8458 ^ _57541;
  wire _57543 = _7864 ^ _3891;
  wire _57544 = _57543 ^ _4615;
  wire _57545 = _57542 ^ _57544;
  wire _57546 = _57540 ^ _57545;
  wire _57547 = _57533 ^ _57546;
  wire _57548 = _4616 ^ _3115;
  wire _57549 = _7265 ^ _46860;
  wire _57550 = _57548 ^ _57549;
  wire _57551 = _13459 ^ _8474;
  wire _57552 = _57551 ^ _12916;
  wire _57553 = _57550 ^ _57552;
  wire _57554 = uncoded_block[1558] ^ uncoded_block[1562];
  wire _57555 = _4637 ^ _57554;
  wire _57556 = _44749 ^ _57555;
  wire _57557 = _4644 ^ _7892;
  wire _57558 = _6029 ^ _6031;
  wire _57559 = _57557 ^ _57558;
  wire _57560 = _57556 ^ _57559;
  wire _57561 = _57553 ^ _57560;
  wire _57562 = _1615 ^ _20401;
  wire _57563 = _24565 ^ _3151;
  wire _57564 = _57562 ^ _57563;
  wire _57565 = _16031 ^ _804;
  wire _57566 = _3155 ^ _57565;
  wire _57567 = _57564 ^ _57566;
  wire _57568 = _16529 ^ _12383;
  wire _57569 = _15550 ^ _57568;
  wire _57570 = _1649 ^ _32178;
  wire _57571 = uncoded_block[1659] ^ uncoded_block[1665];
  wire _57572 = _820 ^ _57571;
  wire _57573 = _57570 ^ _57572;
  wire _57574 = _57569 ^ _57573;
  wire _57575 = _57567 ^ _57574;
  wire _57576 = _57561 ^ _57575;
  wire _57577 = _57547 ^ _57576;
  wire _57578 = _9666 ^ _8521;
  wire _57579 = _48774 ^ _45525;
  wire _57580 = _57578 ^ _57579;
  wire _57581 = _13519 ^ _9675;
  wire _57582 = _57581 ^ _26833;
  wire _57583 = _57580 ^ _57582;
  wire _57584 = _8536 ^ _54215;
  wire _57585 = _57584 ^ uncoded_block[1722];
  wire _57586 = _57583 ^ _57585;
  wire _57587 = _57577 ^ _57586;
  wire _57588 = _57517 ^ _57587;
  wire _57589 = uncoded_block[2] ^ uncoded_block[8];
  wire _57590 = uncoded_block[14] ^ uncoded_block[21];
  wire _57591 = _57589 ^ _57590;
  wire _57592 = uncoded_block[25] ^ uncoded_block[34];
  wire _57593 = _57592 ^ _3230;
  wire _57594 = _57591 ^ _57593;
  wire _57595 = uncoded_block[42] ^ uncoded_block[52];
  wire _57596 = uncoded_block[60] ^ uncoded_block[78];
  wire _57597 = _57595 ^ _57596;
  wire _57598 = _25955 ^ _13558;
  wire _57599 = _57597 ^ _57598;
  wire _57600 = _57594 ^ _57599;
  wire _57601 = uncoded_block[97] ^ uncoded_block[113];
  wire _57602 = _14590 ^ _57601;
  wire _57603 = _6128 ^ _40685;
  wire _57604 = _57602 ^ _57603;
  wire _57605 = uncoded_block[133] ^ uncoded_block[139];
  wire _57606 = uncoded_block[149] ^ uncoded_block[159];
  wire _57607 = _57605 ^ _57606;
  wire _57608 = uncoded_block[171] ^ uncoded_block[179];
  wire _57609 = _39128 ^ _57608;
  wire _57610 = _57607 ^ _57609;
  wire _57611 = _57604 ^ _57610;
  wire _57612 = _57600 ^ _57611;
  wire _57613 = _1759 ^ _6798;
  wire _57614 = uncoded_block[193] ^ uncoded_block[200];
  wire _57615 = _57614 ^ _33082;
  wire _57616 = _57613 ^ _57615;
  wire _57617 = uncoded_block[231] ^ uncoded_block[240];
  wire _57618 = _105 ^ _57617;
  wire _57619 = uncoded_block[250] ^ uncoded_block[259];
  wire _57620 = _57619 ^ _21472;
  wire _57621 = _57618 ^ _57620;
  wire _57622 = _57616 ^ _57621;
  wire _57623 = _2568 ^ _11967;
  wire _57624 = uncoded_block[283] ^ uncoded_block[288];
  wire _57625 = _57624 ^ _995;
  wire _57626 = _57623 ^ _57625;
  wire _57627 = uncoded_block[302] ^ uncoded_block[311];
  wire _57628 = _138 ^ _57627;
  wire _57629 = uncoded_block[317] ^ uncoded_block[325];
  wire _57630 = uncoded_block[326] ^ uncoded_block[334];
  wire _57631 = _57629 ^ _57630;
  wire _57632 = _57628 ^ _57631;
  wire _57633 = _57626 ^ _57632;
  wire _57634 = _57622 ^ _57633;
  wire _57635 = _57612 ^ _57634;
  wire _57636 = _11987 ^ _4844;
  wire _57637 = uncoded_block[380] ^ uncoded_block[391];
  wire _57638 = _10899 ^ _57637;
  wire _57639 = _57636 ^ _57638;
  wire _57640 = uncoded_block[396] ^ uncoded_block[407];
  wire _57641 = _1847 ^ _57640;
  wire _57642 = uncoded_block[413] ^ uncoded_block[424];
  wire _57643 = uncoded_block[426] ^ uncoded_block[436];
  wire _57644 = _57642 ^ _57643;
  wire _57645 = _57641 ^ _57644;
  wire _57646 = _57639 ^ _57645;
  wire _57647 = uncoded_block[445] ^ uncoded_block[464];
  wire _57648 = _3405 ^ _57647;
  wire _57649 = uncoded_block[474] ^ uncoded_block[481];
  wire _57650 = _13665 ^ _57649;
  wire _57651 = _57648 ^ _57650;
  wire _57652 = _4194 ^ _21987;
  wire _57653 = _22445 ^ _17694;
  wire _57654 = _57652 ^ _57653;
  wire _57655 = _57651 ^ _57654;
  wire _57656 = _57646 ^ _57655;
  wire _57657 = _3444 ^ _12039;
  wire _57658 = _1117 ^ _1913;
  wire _57659 = _57657 ^ _57658;
  wire _57660 = _28132 ^ _5635;
  wire _57661 = uncoded_block[581] ^ uncoded_block[597];
  wire _57662 = _57661 ^ _14218;
  wire _57663 = _57660 ^ _57662;
  wire _57664 = _57659 ^ _57663;
  wire _57665 = _14223 ^ _5658;
  wire _57666 = uncoded_block[630] ^ uncoded_block[636];
  wire _57667 = _57666 ^ _5665;
  wire _57668 = _57665 ^ _57667;
  wire _57669 = uncoded_block[649] ^ uncoded_block[660];
  wire _57670 = _2730 ^ _57669;
  wire _57671 = _22037 ^ _15775;
  wire _57672 = _57670 ^ _57671;
  wire _57673 = _57668 ^ _57672;
  wire _57674 = _57664 ^ _57673;
  wire _57675 = _57656 ^ _57674;
  wire _57676 = _57635 ^ _57675;
  wire _57677 = uncoded_block[685] ^ uncoded_block[698];
  wire _57678 = _3522 ^ _57677;
  wire _57679 = _23863 ^ _15785;
  wire _57680 = _57678 ^ _57679;
  wire _57681 = _15301 ^ _359;
  wire _57682 = _8205 ^ _57681;
  wire _57683 = _57680 ^ _57682;
  wire _57684 = uncoded_block[779] ^ uncoded_block[790];
  wire _57685 = _57090 ^ _57684;
  wire _57686 = _57087 ^ _57685;
  wire _57687 = _31551 ^ _16791;
  wire _57688 = _5729 ^ _12135;
  wire _57689 = _57687 ^ _57688;
  wire _57690 = _57686 ^ _57689;
  wire _57691 = _57683 ^ _57690;
  wire _57692 = uncoded_block[832] ^ uncoded_block[843];
  wire _57693 = _57692 ^ _11609;
  wire _57694 = uncoded_block[854] ^ uncoded_block[860];
  wire _57695 = _3599 ^ _57694;
  wire _57696 = _57693 ^ _57695;
  wire _57697 = uncoded_block[872] ^ uncoded_block[890];
  wire _57698 = _12150 ^ _57697;
  wire _57699 = _428 ^ _7663;
  wire _57700 = _57698 ^ _57699;
  wire _57701 = _57696 ^ _57700;
  wire _57702 = _19252 ^ _21182;
  wire _57703 = uncoded_block[929] ^ uncoded_block[939];
  wire _57704 = uncoded_block[944] ^ uncoded_block[961];
  wire _57705 = _57703 ^ _57704;
  wire _57706 = _57702 ^ _57705;
  wire _57707 = _12180 ^ _7088;
  wire _57708 = _57707 ^ _29394;
  wire _57709 = _57706 ^ _57708;
  wire _57710 = _57701 ^ _57709;
  wire _57711 = _57691 ^ _57710;
  wire _57712 = _4401 ^ _483;
  wire _57713 = _57712 ^ _57134;
  wire _57714 = uncoded_block[1043] ^ uncoded_block[1060];
  wire _57715 = _57714 ^ _8888;
  wire _57716 = uncoded_block[1080] ^ uncoded_block[1089];
  wire _57717 = _29859 ^ _57716;
  wire _57718 = _57715 ^ _57717;
  wire _57719 = _57713 ^ _57718;
  wire _57720 = _537 ^ _8910;
  wire _57721 = uncoded_block[1106] ^ uncoded_block[1114];
  wire _57722 = uncoded_block[1127] ^ uncoded_block[1135];
  wire _57723 = _57721 ^ _57722;
  wire _57724 = _57720 ^ _57723;
  wire _57725 = uncoded_block[1138] ^ uncoded_block[1146];
  wire _57726 = _57725 ^ _5866;
  wire _57727 = _11157 ^ _3734;
  wire _57728 = _57726 ^ _57727;
  wire _57729 = _57724 ^ _57728;
  wire _57730 = _57719 ^ _57729;
  wire _57731 = uncoded_block[1166] ^ uncoded_block[1172];
  wire _57732 = _57731 ^ _2195;
  wire _57733 = uncoded_block[1194] ^ uncoded_block[1200];
  wire _57734 = _51363 ^ _57733;
  wire _57735 = _57732 ^ _57734;
  wire _57736 = uncoded_block[1211] ^ uncoded_block[1219];
  wire _57737 = _16399 ^ _57736;
  wire _57738 = uncoded_block[1222] ^ uncoded_block[1237];
  wire _57739 = _57738 ^ _11737;
  wire _57740 = _57737 ^ _57739;
  wire _57741 = _57735 ^ _57740;
  wire _57742 = _6546 ^ _3784;
  wire _57743 = _57742 ^ _24473;
  wire _57744 = _5907 ^ _3793;
  wire _57745 = _57744 ^ _24483;
  wire _57746 = _57743 ^ _57745;
  wire _57747 = _57741 ^ _57746;
  wire _57748 = _57730 ^ _57747;
  wire _57749 = _57711 ^ _57748;
  wire _57750 = _57676 ^ _57749;
  wire _57751 = _35380 ^ _1482;
  wire _57752 = uncoded_block[1314] ^ uncoded_block[1323];
  wire _57753 = uncoded_block[1334] ^ uncoded_block[1342];
  wire _57754 = _57752 ^ _57753;
  wire _57755 = _57751 ^ _57754;
  wire _57756 = uncoded_block[1345] ^ uncoded_block[1361];
  wire _57757 = _57756 ^ _4564;
  wire _57758 = _35792 ^ _35016;
  wire _57759 = _57757 ^ _57758;
  wire _57760 = _57755 ^ _57759;
  wire _57761 = uncoded_block[1408] ^ uncoded_block[1411];
  wire _57762 = _57761 ^ _17470;
  wire _57763 = _1544 ^ _1550;
  wire _57764 = _57762 ^ _57763;
  wire _57765 = uncoded_block[1470] ^ uncoded_block[1480];
  wire _57766 = _57765 ^ _54173;
  wire _57767 = _7864 ^ _7259;
  wire _57768 = _57766 ^ _57767;
  wire _57769 = _57764 ^ _57768;
  wire _57770 = _57760 ^ _57769;
  wire _57771 = _5336 ^ _56921;
  wire _57772 = _12914 ^ _5350;
  wire _57773 = _57771 ^ _57772;
  wire _57774 = _1590 ^ _26792;
  wire _57775 = uncoded_block[1554] ^ uncoded_block[1564];
  wire _57776 = _57775 ^ _37871;
  wire _57777 = _57774 ^ _57776;
  wire _57778 = _57773 ^ _57777;
  wire _57779 = uncoded_block[1570] ^ uncoded_block[1578];
  wire _57780 = _57779 ^ _2383;
  wire _57781 = _32567 ^ _25454;
  wire _57782 = _57780 ^ _57781;
  wire _57783 = _29550 ^ _54931;
  wire _57784 = uncoded_block[1616] ^ uncoded_block[1622];
  wire _57785 = _57784 ^ _3161;
  wire _57786 = _57783 ^ _57785;
  wire _57787 = _57782 ^ _57786;
  wire _57788 = _57778 ^ _57787;
  wire _57789 = _57770 ^ _57788;
  wire _57790 = uncoded_block[1644] ^ uncoded_block[1650];
  wire _57791 = _6048 ^ _57790;
  wire _57792 = _24579 ^ _57242;
  wire _57793 = _57791 ^ _57792;
  wire _57794 = _11324 ^ _2437;
  wire _57795 = _854 ^ _860;
  wire _57796 = _57794 ^ _57795;
  wire _57797 = _57793 ^ _57796;
  wire _57798 = _57797 ^ uncoded_block[1722];
  wire _57799 = _57789 ^ _57798;
  wire _57800 = _57750 ^ _57799;
  wire _57801 = uncoded_block[1] ^ uncoded_block[6];
  wire _57802 = _57801 ^ _32609;
  wire _57803 = uncoded_block[14] ^ uncoded_block[24];
  wire _57804 = _57803 ^ _22333;
  wire _57805 = _57802 ^ _57804;
  wire _57806 = _19006 ^ _12428;
  wire _57807 = _28757 ^ _6742;
  wire _57808 = _57806 ^ _57807;
  wire _57809 = _57805 ^ _57808;
  wire _57810 = _6744 ^ _12438;
  wire _57811 = _28765 ^ _6754;
  wire _57812 = _57810 ^ _57811;
  wire _57813 = uncoded_block[105] ^ uncoded_block[111];
  wire _57814 = _57271 ^ _57813;
  wire _57815 = uncoded_block[118] ^ uncoded_block[124];
  wire _57816 = _43278 ^ _57815;
  wire _57817 = _57814 ^ _57816;
  wire _57818 = _57812 ^ _57817;
  wire _57819 = _57809 ^ _57818;
  wire _57820 = uncoded_block[138] ^ uncoded_block[148];
  wire _57821 = _21898 ^ _57820;
  wire _57822 = uncoded_block[161] ^ uncoded_block[167];
  wire _57823 = _2514 ^ _57822;
  wire _57824 = _57821 ^ _57823;
  wire _57825 = _20979 ^ _5477;
  wire _57826 = uncoded_block[185] ^ uncoded_block[198];
  wire _57827 = _57826 ^ _2537;
  wire _57828 = _57825 ^ _57827;
  wire _57829 = _57824 ^ _57828;
  wire _57830 = _28043 ^ _21459;
  wire _57831 = uncoded_block[216] ^ uncoded_block[231];
  wire _57832 = _57831 ^ _33088;
  wire _57833 = _57830 ^ _57832;
  wire _57834 = _6180 ^ _1785;
  wire _57835 = _15657 ^ _20523;
  wire _57836 = _57834 ^ _57835;
  wire _57837 = _57833 ^ _57836;
  wire _57838 = _57829 ^ _57837;
  wire _57839 = _57819 ^ _57838;
  wire _57840 = _46202 ^ _30104;
  wire _57841 = _20038 ^ _1807;
  wire _57842 = _57840 ^ _57841;
  wire _57843 = uncoded_block[306] ^ uncoded_block[315];
  wire _57844 = _8637 ^ _57843;
  wire _57845 = uncoded_block[316] ^ uncoded_block[322];
  wire _57846 = _57845 ^ _41885;
  wire _57847 = _57844 ^ _57846;
  wire _57848 = _57842 ^ _57847;
  wire _57849 = _34751 ^ _1018;
  wire _57850 = uncoded_block[342] ^ uncoded_block[347];
  wire _57851 = _57850 ^ _2602;
  wire _57852 = _57849 ^ _57851;
  wire _57853 = uncoded_block[369] ^ uncoded_block[376];
  wire _57854 = uncoded_block[379] ^ uncoded_block[386];
  wire _57855 = _57853 ^ _57854;
  wire _57856 = _57855 ^ _40743;
  wire _57857 = _57852 ^ _57856;
  wire _57858 = _57848 ^ _57857;
  wire _57859 = _37991 ^ _13650;
  wire _57860 = _26924 ^ _57859;
  wire _57861 = _27344 ^ _9271;
  wire _57862 = uncoded_block[447] ^ uncoded_block[458];
  wire _57863 = _23349 ^ _57862;
  wire _57864 = _57861 ^ _57863;
  wire _57865 = _57860 ^ _57864;
  wire _57866 = _21522 ^ _4185;
  wire _57867 = uncoded_block[466] ^ uncoded_block[480];
  wire _57868 = _57867 ^ _8694;
  wire _57869 = _57866 ^ _57868;
  wire _57870 = _5604 ^ _1097;
  wire _57871 = _57870 ^ _9296;
  wire _57872 = _57869 ^ _57871;
  wire _57873 = _57865 ^ _57872;
  wire _57874 = _57858 ^ _57873;
  wire _57875 = _57839 ^ _57874;
  wire _57876 = uncoded_block[513] ^ uncoded_block[523];
  wire _57877 = _57876 ^ _3447;
  wire _57878 = uncoded_block[533] ^ uncoded_block[539];
  wire _57879 = _57878 ^ _5628;
  wire _57880 = _57877 ^ _57879;
  wire _57881 = uncoded_block[557] ^ uncoded_block[572];
  wire _57882 = _41147 ^ _57881;
  wire _57883 = _4941 ^ _55572;
  wire _57884 = _57882 ^ _57883;
  wire _57885 = _57880 ^ _57884;
  wire _57886 = _18222 ^ _39621;
  wire _57887 = _3486 ^ _15252;
  wire _57888 = _57886 ^ _57887;
  wire _57889 = uncoded_block[605] ^ uncoded_block[616];
  wire _57890 = _57889 ^ _1153;
  wire _57891 = _57890 ^ _57667;
  wire _57892 = _57888 ^ _57891;
  wire _57893 = _57885 ^ _57892;
  wire _57894 = uncoded_block[650] ^ uncoded_block[659];
  wire _57895 = _29743 ^ _57894;
  wire _57896 = uncoded_block[660] ^ uncoded_block[669];
  wire _57897 = _57896 ^ _14759;
  wire _57898 = _57895 ^ _57897;
  wire _57899 = _3521 ^ _1971;
  wire _57900 = _2755 ^ _12644;
  wire _57901 = _57899 ^ _57900;
  wire _57902 = _57898 ^ _57901;
  wire _57903 = uncoded_block[707] ^ uncoded_block[719];
  wire _57904 = _57903 ^ _4287;
  wire _57905 = _57904 ^ _1997;
  wire _57906 = _14264 ^ _8778;
  wire _57907 = _4298 ^ _5027;
  wire _57908 = _57906 ^ _57907;
  wire _57909 = _57905 ^ _57908;
  wire _57910 = _57902 ^ _57909;
  wire _57911 = _57893 ^ _57910;
  wire _57912 = uncoded_block[771] ^ uncoded_block[778];
  wire _57913 = uncoded_block[782] ^ uncoded_block[789];
  wire _57914 = _57912 ^ _57913;
  wire _57915 = _25696 ^ _2801;
  wire _57916 = _57914 ^ _57915;
  wire _57917 = _31971 ^ _57692;
  wire _57918 = _8229 ^ _57917;
  wire _57919 = _57916 ^ _57918;
  wire _57920 = uncoded_block[844] ^ uncoded_block[852];
  wire _57921 = _57920 ^ _9945;
  wire _57922 = uncoded_block[867] ^ uncoded_block[872];
  wire _57923 = _39676 ^ _57922;
  wire _57924 = _57921 ^ _57923;
  wire _57925 = _33671 ^ _35678;
  wire _57926 = _5085 ^ _45355;
  wire _57927 = _57925 ^ _57926;
  wire _57928 = _57924 ^ _57927;
  wire _57929 = _57919 ^ _57928;
  wire _57930 = uncoded_block[906] ^ uncoded_block[913];
  wire _57931 = _57930 ^ _23917;
  wire _57932 = _5766 ^ _13809;
  wire _57933 = _57931 ^ _57932;
  wire _57934 = _4381 ^ _8845;
  wire _57935 = _36515 ^ _32425;
  wire _57936 = _57934 ^ _57935;
  wire _57937 = _57933 ^ _57936;
  wire _57938 = _32427 ^ _6457;
  wire _57939 = uncoded_block[1009] ^ uncoded_block[1023];
  wire _57940 = _38929 ^ _57939;
  wire _57941 = _57938 ^ _57940;
  wire _57942 = _5138 ^ _11668;
  wire _57943 = _57942 ^ _34111;
  wire _57944 = _57941 ^ _57943;
  wire _57945 = _57937 ^ _57944;
  wire _57946 = _57929 ^ _57945;
  wire _57947 = _57911 ^ _57946;
  wire _57948 = _57875 ^ _57947;
  wire _57949 = uncoded_block[1057] ^ uncoded_block[1064];
  wire _57950 = _4430 ^ _57949;
  wire _57951 = _5828 ^ _20251;
  wire _57952 = _57950 ^ _57951;
  wire _57953 = uncoded_block[1083] ^ uncoded_block[1094];
  wire _57954 = _57953 ^ _5169;
  wire _57955 = _19794 ^ _552;
  wire _57956 = _57954 ^ _57955;
  wire _57957 = _57952 ^ _57956;
  wire _57958 = uncoded_block[1121] ^ uncoded_block[1128];
  wire _57959 = _32873 ^ _57958;
  wire _57960 = uncoded_block[1133] ^ uncoded_block[1141];
  wire _57961 = _57960 ^ _10597;
  wire _57962 = _57959 ^ _57961;
  wire _57963 = _8356 ^ _49385;
  wire _57964 = _27111 ^ _27539;
  wire _57965 = _57963 ^ _57964;
  wire _57966 = _57962 ^ _57965;
  wire _57967 = _57957 ^ _57966;
  wire _57968 = uncoded_block[1192] ^ uncoded_block[1203];
  wire _57969 = uncoded_block[1204] ^ uncoded_block[1214];
  wire _57970 = _57968 ^ _57969;
  wire _57971 = uncoded_block[1224] ^ uncoded_block[1234];
  wire _57972 = _15921 ^ _57971;
  wire _57973 = _57970 ^ _57972;
  wire _57974 = _2989 ^ _14416;
  wire _57975 = _6550 ^ _19834;
  wire _57976 = _57974 ^ _57975;
  wire _57977 = _57973 ^ _57976;
  wire _57978 = uncoded_block[1281] ^ uncoded_block[1287];
  wire _57979 = _57978 ^ _9545;
  wire _57980 = _7799 ^ _26276;
  wire _57981 = _57979 ^ _57980;
  wire _57982 = _3811 ^ _7805;
  wire _57983 = uncoded_block[1322] ^ uncoded_block[1329];
  wire _57984 = _57983 ^ _5256;
  wire _57985 = _57982 ^ _57984;
  wire _57986 = _57981 ^ _57985;
  wire _57987 = _57977 ^ _57986;
  wire _57988 = _57967 ^ _57987;
  wire _57989 = _1495 ^ _1497;
  wire _57990 = _8417 ^ _4558;
  wire _57991 = _57989 ^ _57990;
  wire _57992 = uncoded_block[1361] ^ uncoded_block[1368];
  wire _57993 = _4559 ^ _57992;
  wire _57994 = uncoded_block[1370] ^ uncoded_block[1377];
  wire _57995 = _57994 ^ _16451;
  wire _57996 = _57993 ^ _57995;
  wire _57997 = _57991 ^ _57996;
  wire _57998 = _5288 ^ _5955;
  wire _57999 = _10678 ^ _26301;
  wire _58000 = _57998 ^ _57999;
  wire _58001 = uncoded_block[1422] ^ uncoded_block[1433];
  wire _58002 = _58001 ^ _3857;
  wire _58003 = uncoded_block[1446] ^ uncoded_block[1452];
  wire _58004 = _4590 ^ _58003;
  wire _58005 = _58002 ^ _58004;
  wire _58006 = _58000 ^ _58005;
  wire _58007 = _57997 ^ _58006;
  wire _58008 = _2335 ^ _3096;
  wire _58009 = _42516 ^ _58008;
  wire _58010 = _16977 ^ _31294;
  wire _58011 = _25426 ^ _11264;
  wire _58012 = _58010 ^ _58011;
  wire _58013 = _58009 ^ _58012;
  wire _58014 = _15002 ^ _26321;
  wire _58015 = uncoded_block[1527] ^ uncoded_block[1533];
  wire _58016 = _3118 ^ _58015;
  wire _58017 = _58014 ^ _58016;
  wire _58018 = uncoded_block[1553] ^ uncoded_block[1559];
  wire _58019 = _16995 ^ _58018;
  wire _58020 = uncoded_block[1564] ^ uncoded_block[1580];
  wire _58021 = _3139 ^ _58020;
  wire _58022 = _58019 ^ _58021;
  wire _58023 = _58017 ^ _58022;
  wire _58024 = _58013 ^ _58023;
  wire _58025 = _58007 ^ _58024;
  wire _58026 = _57988 ^ _58025;
  wire _58027 = uncoded_block[1595] ^ uncoded_block[1617];
  wire _58028 = _16025 ^ _58027;
  wire _58029 = uncoded_block[1639] ^ uncoded_block[1647];
  wire _58030 = _17022 ^ _58029;
  wire _58031 = _58028 ^ _58030;
  wire _58032 = _14530 ^ _10761;
  wire _58033 = uncoded_block[1662] ^ uncoded_block[1667];
  wire _58034 = uncoded_block[1672] ^ uncoded_block[1684];
  wire _58035 = _58033 ^ _58034;
  wire _58036 = _58032 ^ _58035;
  wire _58037 = _58031 ^ _58036;
  wire _58038 = _4694 ^ _3968;
  wire _58039 = _11327 ^ _2438;
  wire _58040 = _58038 ^ _58039;
  wire _58041 = _3200 ^ uncoded_block[1721];
  wire _58042 = _58040 ^ _58041;
  wire _58043 = _58037 ^ _58042;
  wire _58044 = _58026 ^ _58043;
  wire _58045 = _57948 ^ _58044;
  wire _58046 = _10787 ^ _30034;
  wire _58047 = _3998 ^ _2458;
  wire _58048 = _58046 ^ _58047;
  wire _58049 = _35096 ^ _25941;
  wire _58050 = uncoded_block[34] ^ uncoded_block[41];
  wire _58051 = _58050 ^ _12425;
  wire _58052 = _58049 ^ _58051;
  wire _58053 = _58048 ^ _58052;
  wire _58054 = uncoded_block[57] ^ uncoded_block[70];
  wire _58055 = _48418 ^ _58054;
  wire _58056 = _897 ^ _28765;
  wire _58057 = _58055 ^ _58056;
  wire _58058 = _41 ^ _2487;
  wire _58059 = _7374 ^ _14068;
  wire _58060 = _58058 ^ _58059;
  wire _58061 = _58057 ^ _58060;
  wire _58062 = _58053 ^ _58061;
  wire _58063 = uncoded_block[106] ^ uncoded_block[116];
  wire _58064 = _11909 ^ _58063;
  wire _58065 = _2497 ^ _25070;
  wire _58066 = _58064 ^ _58065;
  wire _58067 = uncoded_block[124] ^ uncoded_block[130];
  wire _58068 = _58067 ^ _1735;
  wire _58069 = _58068 ^ _10260;
  wire _58070 = _58066 ^ _58069;
  wire _58071 = _15620 ^ _24178;
  wire _58072 = _58071 ^ _55478;
  wire _58073 = uncoded_block[155] ^ uncoded_block[169];
  wire _58074 = _5469 ^ _58073;
  wire _58075 = _6147 ^ _82;
  wire _58076 = _58074 ^ _58075;
  wire _58077 = _58072 ^ _58076;
  wire _58078 = _58070 ^ _58077;
  wire _58079 = _58062 ^ _58078;
  wire _58080 = _49664 ^ _6797;
  wire _58081 = _3283 ^ _25983;
  wire _58082 = _58080 ^ _58081;
  wire _58083 = _6806 ^ _3292;
  wire _58084 = _9202 ^ _17617;
  wire _58085 = _58083 ^ _58084;
  wire _58086 = _58082 ^ _58085;
  wire _58087 = uncoded_block[226] ^ uncoded_block[231];
  wire _58088 = _58087 ^ _2550;
  wire _58089 = _58088 ^ _50046;
  wire _58090 = _7432 ^ _13053;
  wire _58091 = _3311 ^ _120;
  wire _58092 = _58090 ^ _58091;
  wire _58093 = _58089 ^ _58092;
  wire _58094 = _58086 ^ _58093;
  wire _58095 = uncoded_block[271] ^ uncoded_block[277];
  wire _58096 = _4099 ^ _58095;
  wire _58097 = _20527 ^ _7446;
  wire _58098 = _58096 ^ _58097;
  wire _58099 = _28065 ^ _8052;
  wire _58100 = _43316 ^ _58099;
  wire _58101 = _58098 ^ _58100;
  wire _58102 = _3337 ^ _15168;
  wire _58103 = uncoded_block[325] ^ uncoded_block[328];
  wire _58104 = _1008 ^ _58103;
  wire _58105 = _58102 ^ _58104;
  wire _58106 = _33112 ^ _2592;
  wire _58107 = _58106 ^ _33539;
  wire _58108 = _58105 ^ _58107;
  wire _58109 = _58101 ^ _58108;
  wire _58110 = _58094 ^ _58109;
  wire _58111 = _58079 ^ _58110;
  wire _58112 = _8069 ^ _39567;
  wire _58113 = _10898 ^ _10901;
  wire _58114 = _58112 ^ _58113;
  wire _58115 = _13644 ^ _4152;
  wire _58116 = _28845 ^ _6244;
  wire _58117 = _58115 ^ _58116;
  wire _58118 = _58114 ^ _58117;
  wire _58119 = _11473 ^ _43717;
  wire _58120 = _14689 ^ _16187;
  wire _58121 = _58119 ^ _58120;
  wire _58122 = _21516 ^ _12559;
  wire _58123 = uncoded_block[446] ^ uncoded_block[451];
  wire _58124 = uncoded_block[452] ^ uncoded_block[462];
  wire _58125 = _58123 ^ _58124;
  wire _58126 = _58122 ^ _58125;
  wire _58127 = _58121 ^ _58126;
  wire _58128 = _58118 ^ _58127;
  wire _58129 = _13665 ^ _2657;
  wire _58130 = _58129 ^ _40762;
  wire _58131 = uncoded_block[498] ^ uncoded_block[503];
  wire _58132 = _6919 ^ _58131;
  wire _58133 = _20088 ^ _4908;
  wire _58134 = _58132 ^ _58133;
  wire _58135 = _58130 ^ _58134;
  wire _58136 = uncoded_block[512] ^ uncoded_block[518];
  wire _58137 = _58136 ^ _8708;
  wire _58138 = _10948 ^ _1905;
  wire _58139 = _58137 ^ _58138;
  wire _58140 = uncoded_block[561] ^ uncoded_block[567];
  wire _58141 = _14204 ^ _58140;
  wire _58142 = _13690 ^ _58141;
  wire _58143 = _58139 ^ _58142;
  wire _58144 = _58135 ^ _58143;
  wire _58145 = _58128 ^ _58144;
  wire _58146 = _12057 ^ _1933;
  wire _58147 = uncoded_block[595] ^ uncoded_block[599];
  wire _58148 = _58147 ^ _15252;
  wire _58149 = _58146 ^ _58148;
  wire _58150 = uncoded_block[608] ^ uncoded_block[613];
  wire _58151 = _58150 ^ _21098;
  wire _58152 = _4243 ^ _4247;
  wire _58153 = _58151 ^ _58152;
  wire _58154 = _58149 ^ _58153;
  wire _58155 = _1157 ^ _11543;
  wire _58156 = _10985 ^ _10427;
  wire _58157 = _58155 ^ _58156;
  wire _58158 = _18705 ^ _2742;
  wire _58159 = _58158 ^ _25661;
  wire _58160 = _58157 ^ _58159;
  wire _58161 = _58154 ^ _58160;
  wire _58162 = _40802 ^ _36026;
  wire _58163 = uncoded_block[693] ^ uncoded_block[698];
  wire _58164 = _26557 ^ _58163;
  wire _58165 = uncoded_block[709] ^ uncoded_block[716];
  wire _58166 = _58165 ^ _12648;
  wire _58167 = _58164 ^ _58166;
  wire _58168 = _58162 ^ _58167;
  wire _58169 = uncoded_block[726] ^ uncoded_block[731];
  wire _58170 = _58169 ^ _7002;
  wire _58171 = _1995 ^ _36040;
  wire _58172 = _58170 ^ _58171;
  wire _58173 = _2775 ^ _12663;
  wire _58174 = _4298 ^ _9914;
  wire _58175 = _58173 ^ _58174;
  wire _58176 = _58172 ^ _58175;
  wire _58177 = _58168 ^ _58176;
  wire _58178 = _58161 ^ _58177;
  wire _58179 = _58145 ^ _58178;
  wire _58180 = _58111 ^ _58179;
  wire _58181 = _7616 ^ _22063;
  wire _58182 = uncoded_block[793] ^ uncoded_block[801];
  wire _58183 = _43031 ^ _58182;
  wire _58184 = _58181 ^ _58183;
  wire _58185 = _5042 ^ _4324;
  wire _58186 = _37301 ^ _58185;
  wire _58187 = _58184 ^ _58186;
  wire _58188 = _30246 ^ _21158;
  wire _58189 = _42703 ^ _33239;
  wire _58190 = _6406 ^ _408;
  wire _58191 = _58189 ^ _58190;
  wire _58192 = _58188 ^ _58191;
  wire _58193 = _58187 ^ _58192;
  wire _58194 = _2827 ^ _18302;
  wire _58195 = _12151 ^ _4351;
  wire _58196 = _58194 ^ _58195;
  wire _58197 = uncoded_block[890] ^ uncoded_block[899];
  wire _58198 = _4352 ^ _58197;
  wire _58199 = uncoded_block[902] ^ uncoded_block[907];
  wire _58200 = _58199 ^ _1285;
  wire _58201 = _58198 ^ _58200;
  wire _58202 = _58196 ^ _58201;
  wire _58203 = _6430 ^ _17318;
  wire _58204 = _29379 ^ _21649;
  wire _58205 = _58203 ^ _58204;
  wire _58206 = _8839 ^ _22559;
  wire _58207 = _5104 ^ _1307;
  wire _58208 = _58206 ^ _58207;
  wire _58209 = _58205 ^ _58208;
  wire _58210 = _58202 ^ _58209;
  wire _58211 = _58193 ^ _58210;
  wire _58212 = _1308 ^ _22112;
  wire _58213 = _19268 ^ _28233;
  wire _58214 = _58212 ^ _58213;
  wire _58215 = _28235 ^ _2106;
  wire _58216 = _58214 ^ _58215;
  wire _58217 = _23945 ^ _22122;
  wire _58218 = _58217 ^ _27078;
  wire _58219 = _2894 ^ _2126;
  wire _58220 = _2127 ^ _12198;
  wire _58221 = _58219 ^ _58220;
  wire _58222 = _58218 ^ _58221;
  wire _58223 = _58216 ^ _58222;
  wire _58224 = _6475 ^ _515;
  wire _58225 = _58224 ^ _15872;
  wire _58226 = _11125 ^ _2925;
  wire _58227 = _3690 ^ _58226;
  wire _58228 = _58225 ^ _58227;
  wire _58229 = _26225 ^ _11137;
  wire _58230 = _5843 ^ _545;
  wire _58231 = _58229 ^ _58230;
  wire _58232 = _8914 ^ _36134;
  wire _58233 = uncoded_block[1135] ^ uncoded_block[1145];
  wire _58234 = _13866 ^ _58233;
  wire _58235 = _58232 ^ _58234;
  wire _58236 = _58231 ^ _58235;
  wire _58237 = _58228 ^ _58236;
  wire _58238 = _58223 ^ _58237;
  wire _58239 = _58211 ^ _58238;
  wire _58240 = _5184 ^ _29439;
  wire _58241 = _58240 ^ _37776;
  wire _58242 = _10046 ^ _52928;
  wire _58243 = _31637 ^ _35354;
  wire _58244 = _58242 ^ _58243;
  wire _58245 = _58241 ^ _58244;
  wire _58246 = _597 ^ _2207;
  wire _58247 = _6529 ^ _2981;
  wire _58248 = _58246 ^ _58247;
  wire _58249 = _606 ^ _2986;
  wire _58250 = _15927 ^ _5221;
  wire _58251 = _58249 ^ _58250;
  wire _58252 = _58248 ^ _58251;
  wire _58253 = _58245 ^ _58252;
  wire _58254 = uncoded_block[1247] ^ uncoded_block[1250];
  wire _58255 = _11734 ^ _58254;
  wire _58256 = _3784 ^ _53846;
  wire _58257 = _58255 ^ _58256;
  wire _58258 = _9533 ^ _16419;
  wire _58259 = _58258 ^ _19364;
  wire _58260 = _58257 ^ _58259;
  wire _58261 = uncoded_block[1289] ^ uncoded_block[1296];
  wire _58262 = _58261 ^ _3017;
  wire _58263 = _20812 ^ _6572;
  wire _58264 = _58262 ^ _58263;
  wire _58265 = _20314 ^ _14432;
  wire _58266 = _2262 ^ _1487;
  wire _58267 = _58265 ^ _58266;
  wire _58268 = _58264 ^ _58267;
  wire _58269 = _58260 ^ _58268;
  wire _58270 = _58253 ^ _58269;
  wire _58271 = uncoded_block[1336] ^ uncoded_block[1343];
  wire _58272 = _4551 ^ _58271;
  wire _58273 = _50288 ^ _58272;
  wire _58274 = _13401 ^ _16942;
  wire _58275 = _58274 ^ _16443;
  wire _58276 = _58273 ^ _58275;
  wire _58277 = uncoded_block[1381] ^ uncoded_block[1387];
  wire _58278 = _5275 ^ _58277;
  wire _58279 = _692 ^ _3065;
  wire _58280 = _58278 ^ _58279;
  wire _58281 = _4572 ^ _1519;
  wire _58282 = _1523 ^ _704;
  wire _58283 = _58281 ^ _58282;
  wire _58284 = _58280 ^ _58283;
  wire _58285 = _58276 ^ _58284;
  wire _58286 = _13429 ^ _1530;
  wire _58287 = _9595 ^ _20357;
  wire _58288 = _58286 ^ _58287;
  wire _58289 = _26763 ^ _12332;
  wire _58290 = uncoded_block[1463] ^ uncoded_block[1471];
  wire _58291 = _723 ^ _58290;
  wire _58292 = _58289 ^ _58291;
  wire _58293 = _58288 ^ _58292;
  wire _58294 = _10704 ^ _2349;
  wire _58295 = _9614 ^ _12898;
  wire _58296 = _58294 ^ _58295;
  wire _58297 = _3109 ^ _7259;
  wire _58298 = _58297 ^ _56128;
  wire _58299 = _58296 ^ _58298;
  wire _58300 = _58293 ^ _58299;
  wire _58301 = _58285 ^ _58300;
  wire _58302 = _58270 ^ _58301;
  wire _58303 = _58239 ^ _58302;
  wire _58304 = _58180 ^ _58303;
  wire _58305 = _16988 ^ _8473;
  wire _58306 = _34223 ^ _58305;
  wire _58307 = _23198 ^ _26789;
  wire _58308 = _58306 ^ _58307;
  wire _58309 = uncoded_block[1540] ^ uncoded_block[1544];
  wire _58310 = _58309 ^ _18492;
  wire _58311 = uncoded_block[1554] ^ uncoded_block[1561];
  wire _58312 = _7277 ^ _58311;
  wire _58313 = _58310 ^ _58312;
  wire _58314 = uncoded_block[1574] ^ uncoded_block[1579];
  wire _58315 = _4644 ^ _58314;
  wire _58316 = _784 ^ _3927;
  wire _58317 = _58315 ^ _58316;
  wire _58318 = _58313 ^ _58317;
  wire _58319 = _58308 ^ _58318;
  wire _58320 = _791 ^ _11295;
  wire _58321 = _9088 ^ _49971;
  wire _58322 = _58320 ^ _58321;
  wire _58323 = _3946 ^ _57234;
  wire _58324 = _48018 ^ _58323;
  wire _58325 = _58322 ^ _58324;
  wire _58326 = uncoded_block[1652] ^ uncoded_block[1666];
  wire _58327 = _2412 ^ _58326;
  wire _58328 = _2422 ^ _7323;
  wire _58329 = _58327 ^ _58328;
  wire _58330 = uncoded_block[1675] ^ uncoded_block[1684];
  wire _58331 = _58330 ^ _839;
  wire _58332 = _25037 ^ _8536;
  wire _58333 = _58331 ^ _58332;
  wire _58334 = _58329 ^ _58333;
  wire _58335 = _58325 ^ _58334;
  wire _58336 = _58319 ^ _58335;
  wire _58337 = _25928 ^ _12976;
  wire _58338 = _853 ^ _58337;
  wire _58339 = _58338 ^ uncoded_block[1722];
  wire _58340 = _58336 ^ _58339;
  wire _58341 = _58304 ^ _58340;
  wire _58342 = _18539 ^ _6724;
  wire _58343 = _14560 ^ _19963;
  wire _58344 = _58342 ^ _58343;
  wire _58345 = _11 ^ _6095;
  wire _58346 = _35869 ^ _58345;
  wire _58347 = _58344 ^ _58346;
  wire _58348 = _15590 ^ _7965;
  wire _58349 = _58348 ^ _20460;
  wire _58350 = _3233 ^ _1700;
  wire _58351 = _58350 ^ _14580;
  wire _58352 = _58349 ^ _58351;
  wire _58353 = _58347 ^ _58352;
  wire _58354 = _19011 ^ _34;
  wire _58355 = uncoded_block[76] ^ uncoded_block[80];
  wire _58356 = _35 ^ _58355;
  wire _58357 = _58354 ^ _58356;
  wire _58358 = _2487 ^ _4026;
  wire _58359 = _35502 ^ _58358;
  wire _58360 = _58357 ^ _58359;
  wire _58361 = _23708 ^ _11911;
  wire _58362 = _46546 ^ _6126;
  wire _58363 = _10816 ^ _6128;
  wire _58364 = _58362 ^ _58363;
  wire _58365 = _58361 ^ _58364;
  wire _58366 = _58360 ^ _58365;
  wire _58367 = _58353 ^ _58366;
  wire _58368 = _10819 ^ _20961;
  wire _58369 = _4754 ^ _47307;
  wire _58370 = _58368 ^ _58369;
  wire _58371 = uncoded_block[142] ^ uncoded_block[148];
  wire _58372 = _58371 ^ _20488;
  wire _58373 = _4049 ^ _21906;
  wire _58374 = _58372 ^ _58373;
  wire _58375 = _58370 ^ _58374;
  wire _58376 = uncoded_block[162] ^ uncoded_block[168];
  wire _58377 = _58376 ^ _1752;
  wire _58378 = _4057 ^ _8009;
  wire _58379 = _58377 ^ _58378;
  wire _58380 = _20500 ^ _11402;
  wire _58381 = _55485 ^ _58380;
  wire _58382 = _58379 ^ _58381;
  wire _58383 = _58375 ^ _58382;
  wire _58384 = uncoded_block[207] ^ uncoded_block[210];
  wire _58385 = _58384 ^ _3295;
  wire _58386 = _17610 ^ _58385;
  wire _58387 = _21461 ^ _20506;
  wire _58388 = _58386 ^ _58387;
  wire _58389 = _11410 ^ _1774;
  wire _58390 = _2550 ^ _7423;
  wire _58391 = _58389 ^ _58390;
  wire _58392 = _9756 ^ _113;
  wire _58393 = uncoded_block[245] ^ uncoded_block[250];
  wire _58394 = _58393 ^ _2557;
  wire _58395 = _58392 ^ _58394;
  wire _58396 = _58391 ^ _58395;
  wire _58397 = _58388 ^ _58396;
  wire _58398 = _58383 ^ _58397;
  wire _58399 = _58367 ^ _58398;
  wire _58400 = _49200 ^ _30977;
  wire _58401 = _4099 ^ _3320;
  wire _58402 = _58401 ^ _11965;
  wire _58403 = _58400 ^ _58402;
  wire _58404 = _134 ^ _31842;
  wire _58405 = _58097 ^ _58404;
  wire _58406 = _35933 ^ _6845;
  wire _58407 = _19076 ^ _58406;
  wire _58408 = _58405 ^ _58407;
  wire _58409 = _58403 ^ _58408;
  wire _58410 = _22866 ^ _15168;
  wire _58411 = _58410 ^ _13080;
  wire _58412 = _11983 ^ _3352;
  wire _58413 = _30560 ^ _58412;
  wire _58414 = _58411 ^ _58413;
  wire _58415 = _3355 ^ _2596;
  wire _58416 = _46217 ^ _58415;
  wire _58417 = _15179 ^ _2601;
  wire _58418 = _6864 ^ _5548;
  wire _58419 = _58417 ^ _58418;
  wire _58420 = _58416 ^ _58419;
  wire _58421 = _58414 ^ _58420;
  wire _58422 = _58409 ^ _58421;
  wire _58423 = _19591 ^ _4855;
  wire _58424 = _1038 ^ _3380;
  wire _58425 = _13644 ^ _1847;
  wire _58426 = _58424 ^ _58425;
  wire _58427 = _58423 ^ _58426;
  wire _58428 = _1849 ^ _181;
  wire _58429 = uncoded_block[406] ^ uncoded_block[410];
  wire _58430 = _183 ^ _58429;
  wire _58431 = _58428 ^ _58430;
  wire _58432 = _24245 ^ _4874;
  wire _58433 = _197 ^ _2638;
  wire _58434 = _58432 ^ _58433;
  wire _58435 = _58431 ^ _58434;
  wire _58436 = _58427 ^ _58435;
  wire _58437 = _10352 ^ _3405;
  wire _58438 = _21052 ^ _33565;
  wire _58439 = _58437 ^ _58438;
  wire _58440 = uncoded_block[468] ^ uncoded_block[474];
  wire _58441 = _7507 ^ _58440;
  wire _58442 = _55913 ^ _58441;
  wire _58443 = _58439 ^ _58442;
  wire _58444 = _21526 ^ _5593;
  wire _58445 = _16200 ^ _14183;
  wire _58446 = _58444 ^ _58445;
  wire _58447 = _27361 ^ _23370;
  wire _58448 = _16204 ^ _58447;
  wire _58449 = _58446 ^ _58448;
  wire _58450 = _58443 ^ _58449;
  wire _58451 = _58436 ^ _58450;
  wire _58452 = _58422 ^ _58451;
  wire _58453 = _58399 ^ _58452;
  wire _58454 = _4918 ^ _9301;
  wire _58455 = _4214 ^ _16215;
  wire _58456 = _58454 ^ _58455;
  wire _58457 = uncoded_block[553] ^ uncoded_block[561];
  wire _58458 = _4931 ^ _58457;
  wire _58459 = _45269 ^ _58458;
  wire _58460 = _58456 ^ _58459;
  wire _58461 = _3464 ^ _32327;
  wire _58462 = _8727 ^ _3472;
  wire _58463 = _58461 ^ _58462;
  wire _58464 = _4946 ^ _37247;
  wire _58465 = _1134 ^ _58464;
  wire _58466 = _58463 ^ _58465;
  wire _58467 = _58460 ^ _58466;
  wire _58468 = _4234 ^ _3480;
  wire _58469 = _10408 ^ _3489;
  wire _58470 = _58468 ^ _58469;
  wire _58471 = uncoded_block[606] ^ uncoded_block[609];
  wire _58472 = _58471 ^ _4242;
  wire _58473 = _281 ^ _1946;
  wire _58474 = _58472 ^ _58473;
  wire _58475 = _58470 ^ _58474;
  wire _58476 = _2720 ^ _1156;
  wire _58477 = _4249 ^ _9343;
  wire _58478 = _58476 ^ _58477;
  wire _58479 = _36017 ^ _10427;
  wire _58480 = _304 ^ _2738;
  wire _58481 = _58479 ^ _58480;
  wire _58482 = _58478 ^ _58481;
  wire _58483 = _58475 ^ _58482;
  wire _58484 = _58467 ^ _58483;
  wire _58485 = _16751 ^ _8760;
  wire _58486 = _7583 ^ _58485;
  wire _58487 = _10440 ^ _18247;
  wire _58488 = _321 ^ _4271;
  wire _58489 = _58487 ^ _58488;
  wire _58490 = _58486 ^ _58489;
  wire _58491 = _5681 ^ _330;
  wire _58492 = _22499 ^ _17266;
  wire _58493 = _50150 ^ _58492;
  wire _58494 = _58491 ^ _58493;
  wire _58495 = _58490 ^ _58494;
  wire _58496 = _340 ^ _12648;
  wire _58497 = _3544 ^ _5693;
  wire _58498 = _58496 ^ _58497;
  wire _58499 = _1991 ^ _23870;
  wire _58500 = _3550 ^ _5013;
  wire _58501 = _58499 ^ _58500;
  wire _58502 = _58498 ^ _58501;
  wire _58503 = _49300 ^ _12664;
  wire _58504 = _58503 ^ _8211;
  wire _58505 = _15799 ^ _3562;
  wire _58506 = _368 ^ _5715;
  wire _58507 = _58505 ^ _58506;
  wire _58508 = _58504 ^ _58507;
  wire _58509 = _58502 ^ _58508;
  wire _58510 = _58495 ^ _58509;
  wire _58511 = _58484 ^ _58510;
  wire _58512 = _1224 ^ _7626;
  wire _58513 = _26588 ^ _7029;
  wire _58514 = _58512 ^ _58513;
  wire _58515 = _5045 ^ _4325;
  wire _58516 = _41215 ^ _58515;
  wire _58517 = _58514 ^ _58516;
  wire _58518 = _15320 ^ _1247;
  wire _58519 = _58518 ^ _25707;
  wire _58520 = _25710 ^ _46711;
  wire _58521 = _17296 ^ _58520;
  wire _58522 = _58519 ^ _58521;
  wire _58523 = _58517 ^ _58522;
  wire _58524 = _15824 ^ _414;
  wire _58525 = uncoded_block[873] ^ uncoded_block[878];
  wire _58526 = _57922 ^ _58525;
  wire _58527 = _58524 ^ _58526;
  wire _58528 = _421 ^ _11059;
  wire _58529 = _11060 ^ _8250;
  wire _58530 = _58528 ^ _58529;
  wire _58531 = _58527 ^ _58530;
  wire _58532 = _28965 ^ _15345;
  wire _58533 = _9424 ^ _23917;
  wire _58534 = _58532 ^ _58533;
  wire _58535 = _439 ^ _5766;
  wire _58536 = _8260 ^ _3637;
  wire _58537 = _58535 ^ _58536;
  wire _58538 = _58534 ^ _58537;
  wire _58539 = _58531 ^ _58538;
  wire _58540 = _58523 ^ _58539;
  wire _58541 = _15848 ^ _9971;
  wire _58542 = uncoded_block[943] ^ uncoded_block[949];
  wire _58543 = _58542 ^ _2869;
  wire _58544 = _58541 ^ _58543;
  wire _58545 = _2090 ^ _10529;
  wire _58546 = _58545 ^ _12181;
  wire _58547 = _58544 ^ _58546;
  wire _58548 = _11649 ^ _4391;
  wire _58549 = _58548 ^ _50209;
  wire _58550 = _24853 ^ _8859;
  wire _58551 = _10543 ^ _13277;
  wire _58552 = _58550 ^ _58551;
  wire _58553 = _58549 ^ _58552;
  wire _58554 = _58547 ^ _58553;
  wire _58555 = _2111 ^ _6459;
  wire _58556 = _58555 ^ _40501;
  wire _58557 = _5131 ^ _1334;
  wire _58558 = uncoded_block[1023] ^ uncoded_block[1031];
  wire _58559 = _58558 ^ _11668;
  wire _58560 = _58557 ^ _58559;
  wire _58561 = _58556 ^ _58560;
  wire _58562 = _1345 ^ _2910;
  wire _58563 = _515 ^ _518;
  wire _58564 = _58562 ^ _58563;
  wire _58565 = _6483 ^ _2140;
  wire _58566 = _32444 ^ _58565;
  wire _58567 = _58564 ^ _58566;
  wire _58568 = _58561 ^ _58567;
  wire _58569 = _58554 ^ _58568;
  wire _58570 = _58540 ^ _58569;
  wire _58571 = _58511 ^ _58570;
  wire _58572 = _58453 ^ _58571;
  wire _58573 = _2143 ^ _3692;
  wire _58574 = _58573 ^ _23971;
  wire _58575 = _51984 ^ _16369;
  wire _58576 = _58574 ^ _58575;
  wire _58577 = _26227 ^ _2164;
  wire _58578 = _58577 ^ _8918;
  wire _58579 = _12782 ^ _11147;
  wire _58580 = _36134 ^ _558;
  wire _58581 = _58579 ^ _58580;
  wire _58582 = _58578 ^ _58581;
  wire _58583 = _58576 ^ _58582;
  wire _58584 = _9494 ^ _14380;
  wire _58585 = _58584 ^ _26235;
  wire _58586 = _38963 ^ _5188;
  wire _58587 = _58586 ^ _5191;
  wire _58588 = _58585 ^ _58587;
  wire _58589 = _22627 ^ _15907;
  wire _58590 = _1408 ^ _52928;
  wire _58591 = _58589 ^ _58590;
  wire _58592 = _10053 ^ _2971;
  wire _58593 = _26687 ^ _58592;
  wire _58594 = _58591 ^ _58593;
  wire _58595 = _58588 ^ _58594;
  wire _58596 = _58583 ^ _58595;
  wire _58597 = _38970 ^ _8951;
  wire _58598 = _58597 ^ _27551;
  wire _58599 = _23106 ^ _31222;
  wire _58600 = _58598 ^ _58599;
  wire _58601 = _5219 ^ _3772;
  wire _58602 = _38977 ^ _58601;
  wire _58603 = _2994 ^ _8963;
  wire _58604 = uncoded_block[1248] ^ uncoded_block[1253];
  wire _58605 = _58604 ^ _5902;
  wire _58606 = _58603 ^ _58605;
  wire _58607 = _58602 ^ _58606;
  wire _58608 = _58600 ^ _58607;
  wire _58609 = _1458 ^ _628;
  wire _58610 = _42769 ^ _58609;
  wire _58611 = _1463 ^ _6556;
  wire _58612 = _638 ^ _5243;
  wire _58613 = _58611 ^ _58612;
  wire _58614 = _58610 ^ _58613;
  wire _58615 = _11195 ^ _30797;
  wire _58616 = uncoded_block[1297] ^ uncoded_block[1303];
  wire _58617 = _3015 ^ _58616;
  wire _58618 = _58615 ^ _58617;
  wire _58619 = _1479 ^ _18423;
  wire _58620 = uncoded_block[1318] ^ uncoded_block[1324];
  wire _58621 = _3811 ^ _58620;
  wire _58622 = _58619 ^ _58621;
  wire _58623 = _58618 ^ _58622;
  wire _58624 = _58614 ^ _58623;
  wire _58625 = _58608 ^ _58624;
  wire _58626 = _58596 ^ _58625;
  wire _58627 = _44316 ^ _8413;
  wire _58628 = uncoded_block[1343] ^ uncoded_block[1350];
  wire _58629 = _13399 ^ _58628;
  wire _58630 = _58627 ^ _58629;
  wire _58631 = _11773 ^ _57192;
  wire _58632 = _28331 ^ _58631;
  wire _58633 = _58630 ^ _58632;
  wire _58634 = uncoded_block[1382] ^ uncoded_block[1385];
  wire _58635 = _7219 ^ _58634;
  wire _58636 = _58635 ^ _7223;
  wire _58637 = _28340 ^ _4572;
  wire _58638 = _3841 ^ _14457;
  wire _58639 = _58637 ^ _58638;
  wire _58640 = _58636 ^ _58639;
  wire _58641 = _58633 ^ _58640;
  wire _58642 = _5296 ^ _17960;
  wire _58643 = _9586 ^ _58642;
  wire _58644 = _16463 ^ _9022;
  wire _58645 = _11239 ^ _15498;
  wire _58646 = _58644 ^ _58645;
  wire _58647 = _58643 ^ _58646;
  wire _58648 = _25863 ^ _37449;
  wire _58649 = _11246 ^ _11249;
  wire _58650 = _9602 ^ _23614;
  wire _58651 = _58649 ^ _58650;
  wire _58652 = _58648 ^ _58651;
  wire _58653 = _58647 ^ _58652;
  wire _58654 = _58641 ^ _58653;
  wire _58655 = _41757 ^ _15994;
  wire _58656 = _10706 ^ _2349;
  wire _58657 = _58655 ^ _58656;
  wire _58658 = _1565 ^ _6631;
  wire _58659 = _2352 ^ _11813;
  wire _58660 = _58658 ^ _58659;
  wire _58661 = _58657 ^ _58660;
  wire _58662 = _24539 ^ _5334;
  wire _58663 = _58662 ^ _39049;
  wire _58664 = _5337 ^ _33818;
  wire _58665 = _9626 ^ _53901;
  wire _58666 = _58664 ^ _58665;
  wire _58667 = _58663 ^ _58666;
  wire _58668 = _58661 ^ _58667;
  wire _58669 = uncoded_block[1535] ^ uncoded_block[1541];
  wire _58670 = _58669 ^ _2370;
  wire _58671 = _58670 ^ _35051;
  wire _58672 = _39056 ^ _18006;
  wire _58673 = _58671 ^ _58672;
  wire _58674 = _2383 ^ _40243;
  wire _58675 = _17008 ^ _58674;
  wire _58676 = _25454 ^ _4654;
  wire _58677 = _12937 ^ _8502;
  wire _58678 = _58676 ^ _58677;
  wire _58679 = _58675 ^ _58678;
  wire _58680 = _58673 ^ _58679;
  wire _58681 = _58668 ^ _58680;
  wire _58682 = _58654 ^ _58681;
  wire _58683 = _58626 ^ _58682;
  wire _58684 = _11849 ^ _4662;
  wire _58685 = _29997 ^ _7911;
  wire _58686 = _58684 ^ _58685;
  wire _58687 = _14006 ^ _2404;
  wire _58688 = _812 ^ _5392;
  wire _58689 = _58687 ^ _58688;
  wire _58690 = _58686 ^ _58689;
  wire _58691 = _2408 ^ _5394;
  wire _58692 = _2412 ^ _24578;
  wire _58693 = _58691 ^ _58692;
  wire _58694 = _12390 ^ _4680;
  wire _58695 = _58694 ^ _35848;
  wire _58696 = _58693 ^ _58695;
  wire _58697 = _58690 ^ _58696;
  wire _58698 = _41009 ^ _11321;
  wire _58699 = uncoded_block[1682] ^ uncoded_block[1687];
  wire _58700 = _10766 ^ _58699;
  wire _58701 = _58698 ^ _58700;
  wire _58702 = uncoded_block[1696] ^ uncoded_block[1700];
  wire _58703 = _840 ^ _58702;
  wire _58704 = _4700 ^ _53943;
  wire _58705 = _58703 ^ _58704;
  wire _58706 = _58701 ^ _58705;
  wire _58707 = _43251 ^ _6720;
  wire _58708 = _58706 ^ _58707;
  wire _58709 = _58697 ^ _58708;
  wire _58710 = _58683 ^ _58709;
  wire _58711 = _58572 ^ _58710;
  wire _58712 = _3210 ^ _19959;
  wire _58713 = _46150 ^ _56963;
  wire _58714 = _58712 ^ _58713;
  wire _58715 = _21416 ^ _1699;
  wire _58716 = _32614 ^ _58715;
  wire _58717 = _58714 ^ _58716;
  wire _58718 = uncoded_block[60] ^ uncoded_block[69];
  wire _58719 = _58718 ^ _897;
  wire _58720 = _58719 ^ _14061;
  wire _58721 = uncoded_block[94] ^ uncoded_block[99];
  wire _58722 = _58721 ^ _6763;
  wire _58723 = _33050 ^ _58722;
  wire _58724 = _58720 ^ _58723;
  wire _58725 = _58717 ^ _58724;
  wire _58726 = _9721 ^ _10256;
  wire _58727 = uncoded_block[129] ^ uncoded_block[137];
  wire _58728 = _917 ^ _58727;
  wire _58729 = _58726 ^ _58728;
  wire _58730 = uncoded_block[140] ^ uncoded_block[146];
  wire _58731 = uncoded_block[156] ^ uncoded_block[161];
  wire _58732 = _58730 ^ _58731;
  wire _58733 = _19536 ^ _2517;
  wire _58734 = _58732 ^ _58733;
  wire _58735 = _58729 ^ _58734;
  wire _58736 = _13032 ^ _5477;
  wire _58737 = uncoded_block[182] ^ uncoded_block[188];
  wire _58738 = uncoded_block[190] ^ uncoded_block[198];
  wire _58739 = _58737 ^ _58738;
  wire _58740 = _58736 ^ _58739;
  wire _58741 = _32248 ^ _58384;
  wire _58742 = _956 ^ _3299;
  wire _58743 = _58741 ^ _58742;
  wire _58744 = _58740 ^ _58743;
  wire _58745 = _58735 ^ _58744;
  wire _58746 = _58725 ^ _58745;
  wire _58747 = uncoded_block[230] ^ uncoded_block[236];
  wire _58748 = uncoded_block[240] ^ uncoded_block[245];
  wire _58749 = _58747 ^ _58748;
  wire _58750 = uncoded_block[246] ^ uncoded_block[250];
  wire _58751 = _58750 ^ _1785;
  wire _58752 = _58749 ^ _58751;
  wire _58753 = _1789 ^ _127;
  wire _58754 = uncoded_block[275] ^ uncoded_block[279];
  wire _58755 = _1793 ^ _58754;
  wire _58756 = _58753 ^ _58755;
  wire _58757 = _58752 ^ _58756;
  wire _58758 = _11424 ^ _3327;
  wire _58759 = _4819 ^ _28065;
  wire _58760 = _58758 ^ _58759;
  wire _58761 = uncoded_block[307] ^ uncoded_block[317];
  wire _58762 = _6845 ^ _58761;
  wire _58763 = _29245 ^ _1819;
  wire _58764 = _58762 ^ _58763;
  wire _58765 = _58760 ^ _58764;
  wire _58766 = _58757 ^ _58765;
  wire _58767 = _6217 ^ _4131;
  wire _58768 = _58767 ^ _18155;
  wire _58769 = uncoded_block[357] ^ uncoded_block[376];
  wire _58770 = _58769 ^ _1841;
  wire _58771 = _1039 ^ _177;
  wire _58772 = _58770 ^ _58771;
  wire _58773 = _58768 ^ _58772;
  wire _58774 = _33128 ^ _16177;
  wire _58775 = uncoded_block[408] ^ uncoded_block[417];
  wire _58776 = _58775 ^ _11479;
  wire _58777 = _58774 ^ _58776;
  wire _58778 = _3411 ^ _5584;
  wire _58779 = _37610 ^ _58778;
  wire _58780 = _58777 ^ _58779;
  wire _58781 = _58773 ^ _58780;
  wire _58782 = _58766 ^ _58781;
  wire _58783 = _58746 ^ _58782;
  wire _58784 = _1079 ^ _58440;
  wire _58785 = _4891 ^ _58784;
  wire _58786 = _33570 ^ _32309;
  wire _58787 = _21987 ^ _7529;
  wire _58788 = _58786 ^ _58787;
  wire _58789 = _58785 ^ _58788;
  wire _58790 = _3437 ^ _29289;
  wire _58791 = _4918 ^ _4921;
  wire _58792 = _58790 ^ _58791;
  wire _58793 = _33587 ^ _14198;
  wire _58794 = _48151 ^ _3467;
  wire _58795 = _58793 ^ _58794;
  wire _58796 = _58792 ^ _58795;
  wire _58797 = _58789 ^ _58796;
  wire _58798 = _8727 ^ _10400;
  wire _58799 = _58798 ^ _16229;
  wire _58800 = _2706 ^ _14218;
  wire _58801 = _16238 ^ _17238;
  wire _58802 = _58800 ^ _58801;
  wire _58803 = _58799 ^ _58802;
  wire _58804 = _43761 ^ _3502;
  wire _58805 = uncoded_block[651] ^ uncoded_block[660];
  wire _58806 = _10425 ^ _58805;
  wire _58807 = _58804 ^ _58806;
  wire _58808 = _13190 ^ _16752;
  wire _58809 = _58808 ^ _6350;
  wire _58810 = _58807 ^ _58809;
  wire _58811 = _58803 ^ _58810;
  wire _58812 = _58797 ^ _58811;
  wire _58813 = _35635 ^ _44559;
  wire _58814 = _41180 ^ _11562;
  wire _58815 = _58813 ^ _58814;
  wire _58816 = _3533 ^ _33204;
  wire _58817 = uncoded_block[731] ^ uncoded_block[737];
  wire _58818 = _1194 ^ _58817;
  wire _58819 = _58816 ^ _58818;
  wire _58820 = _58815 ^ _58819;
  wire _58821 = uncoded_block[748] ^ uncoded_block[754];
  wire _58822 = _13208 ^ _58821;
  wire _58823 = _58822 ^ _14781;
  wire _58824 = uncoded_block[771] ^ uncoded_block[776];
  wire _58825 = _58824 ^ _17284;
  wire _58826 = _43418 ^ _58825;
  wire _58827 = _58823 ^ _58826;
  wire _58828 = _58820 ^ _58827;
  wire _58829 = _4309 ^ _1224;
  wire _58830 = _4314 ^ _54752;
  wire _58831 = _58829 ^ _58830;
  wire _58832 = _24807 ^ _33655;
  wire _58833 = _58831 ^ _58832;
  wire _58834 = _1253 ^ _11043;
  wire _58835 = _9405 ^ _2046;
  wire _58836 = _58834 ^ _58835;
  wire _58837 = _34476 ^ _17304;
  wire _58838 = uncoded_block[889] ^ uncoded_block[900];
  wire _58839 = _53198 ^ _58838;
  wire _58840 = _58837 ^ _58839;
  wire _58841 = _58836 ^ _58840;
  wire _58842 = _58833 ^ _58841;
  wire _58843 = _58828 ^ _58842;
  wire _58844 = _58812 ^ _58843;
  wire _58845 = _58783 ^ _58844;
  wire _58846 = uncoded_block[917] ^ uncoded_block[924];
  wire _58847 = _435 ^ _58846;
  wire _58848 = _7664 ^ _58847;
  wire _58849 = _41240 ^ _9971;
  wire _58850 = _9433 ^ _21191;
  wire _58851 = _58849 ^ _58850;
  wire _58852 = _58848 ^ _58851;
  wire _58853 = _2871 ^ _8847;
  wire _58854 = uncoded_block[974] ^ uncoded_block[981];
  wire _58855 = uncoded_block[983] ^ uncoded_block[991];
  wire _58856 = _58854 ^ _58855;
  wire _58857 = _58853 ^ _58856;
  wire _58858 = _6459 ^ _21206;
  wire _58859 = _37346 ^ _58858;
  wire _58860 = _58857 ^ _58859;
  wire _58861 = _58852 ^ _58860;
  wire _58862 = _1331 ^ _27494;
  wire _58863 = _14857 ^ _1346;
  wire _58864 = _58862 ^ _58863;
  wire _58865 = uncoded_block[1050] ^ uncoded_block[1055];
  wire _58866 = _54805 ^ _58865;
  wire _58867 = _38944 ^ _2921;
  wire _58868 = _58866 ^ _58867;
  wire _58869 = _58864 ^ _58868;
  wire _58870 = uncoded_block[1071] ^ uncoded_block[1080];
  wire _58871 = _5828 ^ _58870;
  wire _58872 = _10575 ^ _11687;
  wire _58873 = _58871 ^ _58872;
  wire _58874 = _23508 ^ _5843;
  wire _58875 = uncoded_block[1100] ^ uncoded_block[1114];
  wire _58876 = _58875 ^ _13322;
  wire _58877 = _58874 ^ _58876;
  wire _58878 = _58873 ^ _58877;
  wire _58879 = _58869 ^ _58878;
  wire _58880 = _58861 ^ _58879;
  wire _58881 = _10587 ^ _5859;
  wire _58882 = uncoded_block[1143] ^ uncoded_block[1148];
  wire _58883 = _58882 ^ _2956;
  wire _58884 = _58881 ^ _58883;
  wire _58885 = _8937 ^ _2964;
  wire _58886 = uncoded_block[1169] ^ uncoded_block[1177];
  wire _58887 = uncoded_block[1179] ^ uncoded_block[1186];
  wire _58888 = _58886 ^ _58887;
  wire _58889 = _58885 ^ _58888;
  wire _58890 = _58884 ^ _58889;
  wire _58891 = _6525 ^ _7163;
  wire _58892 = _21716 ^ _58891;
  wire _58893 = _27911 ^ _608;
  wire _58894 = _30773 ^ _40166;
  wire _58895 = _58893 ^ _58894;
  wire _58896 = _58892 ^ _58895;
  wire _58897 = _58890 ^ _58896;
  wire _58898 = _13360 ^ _5221;
  wire _58899 = _23114 ^ _32082;
  wire _58900 = _58898 ^ _58899;
  wire _58901 = _7781 ^ _5235;
  wire _58902 = uncoded_block[1270] ^ uncoded_block[1274];
  wire _58903 = _3008 ^ _58902;
  wire _58904 = _58901 ^ _58903;
  wire _58905 = _58900 ^ _58904;
  wire _58906 = _10638 ^ _16924;
  wire _58907 = _18866 ^ _21741;
  wire _58908 = _58906 ^ _58907;
  wire _58909 = _5248 ^ _1482;
  wire _58910 = uncoded_block[1313] ^ uncoded_block[1324];
  wire _58911 = _58910 ^ _10655;
  wire _58912 = _58909 ^ _58911;
  wire _58913 = _58908 ^ _58912;
  wire _58914 = _58905 ^ _58913;
  wire _58915 = _58897 ^ _58914;
  wire _58916 = _58880 ^ _58915;
  wire _58917 = _14437 ^ _5262;
  wire _58918 = uncoded_block[1350] ^ uncoded_block[1355];
  wire _58919 = _3039 ^ _58918;
  wire _58920 = _58917 ^ _58919;
  wire _58921 = _15477 ^ _677;
  wire _58922 = _10665 ^ _11226;
  wire _58923 = _58921 ^ _58922;
  wire _58924 = _58920 ^ _58923;
  wire _58925 = _7824 ^ _3834;
  wire _58926 = _10108 ^ _691;
  wire _58927 = _58925 ^ _58926;
  wire _58928 = _35016 ^ _9016;
  wire _58929 = uncoded_block[1408] ^ uncoded_block[1417];
  wire _58930 = _58929 ^ _7842;
  wire _58931 = _58928 ^ _58930;
  wire _58932 = _58927 ^ _58931;
  wire _58933 = _58924 ^ _58932;
  wire _58934 = uncoded_block[1428] ^ uncoded_block[1432];
  wire _58935 = _5967 ^ _58934;
  wire _58936 = _20355 ^ _14983;
  wire _58937 = _58935 ^ _58936;
  wire _58938 = _720 ^ _13440;
  wire _58939 = uncoded_block[1474] ^ uncoded_block[1481];
  wire _58940 = _22254 ^ _58939;
  wire _58941 = _58938 ^ _58940;
  wire _58942 = _58937 ^ _58941;
  wire _58943 = uncoded_block[1491] ^ uncoded_block[1498];
  wire _58944 = _50324 ^ _58943;
  wire _58945 = uncoded_block[1509] ^ uncoded_block[1519];
  wire _58946 = _11813 ^ _58945;
  wire _58947 = _58944 ^ _58946;
  wire _58948 = _23194 ^ _53901;
  wire _58949 = _58948 ^ _47237;
  wire _58950 = _58947 ^ _58949;
  wire _58951 = _58942 ^ _58950;
  wire _58952 = _58933 ^ _58951;
  wire _58953 = _1589 ^ _5355;
  wire _58954 = _7275 ^ _16016;
  wire _58955 = _58953 ^ _58954;
  wire _58956 = _26794 ^ _16019;
  wire _58957 = uncoded_block[1579] ^ uncoded_block[1590];
  wire _58958 = _15535 ^ _58957;
  wire _58959 = _58956 ^ _58958;
  wire _58960 = _58955 ^ _58959;
  wire _58961 = _3146 ^ _4654;
  wire _58962 = _6674 ^ _40633;
  wire _58963 = _58961 ^ _58962;
  wire _58964 = uncoded_block[1620] ^ uncoded_block[1625];
  wire _58965 = _49471 ^ _58964;
  wire _58966 = uncoded_block[1638] ^ uncoded_block[1649];
  wire _58967 = _18511 ^ _58966;
  wire _58968 = _58965 ^ _58967;
  wire _58969 = _58963 ^ _58968;
  wire _58970 = _58960 ^ _58969;
  wire _58971 = _8515 ^ _36687;
  wire _58972 = _17032 ^ _37892;
  wire _58973 = _58971 ^ _58972;
  wire _58974 = _37895 ^ _39083;
  wire _58975 = _9118 ^ _10214;
  wire _58976 = _58974 ^ _58975;
  wire _58977 = _58973 ^ _58976;
  wire _58978 = _41018 ^ uncoded_block[1722];
  wire _58979 = _58977 ^ _58978;
  wire _58980 = _58970 ^ _58979;
  wire _58981 = _58952 ^ _58980;
  wire _58982 = _58916 ^ _58981;
  wire _58983 = _58845 ^ _58982;
  wire _58984 = uncoded_block[10] ^ uncoded_block[18];
  wire _58985 = _24147 ^ _58984;
  wire _58986 = _56963 ^ _11344;
  wire _58987 = _58985 ^ _58986;
  wire _58988 = _37116 ^ _19006;
  wire _58989 = _58988 ^ _32213;
  wire _58990 = _58987 ^ _58989;
  wire _58991 = uncoded_block[59] ^ uncoded_block[68];
  wire _58992 = _58991 ^ _4733;
  wire _58993 = uncoded_block[80] ^ uncoded_block[83];
  wire _58994 = _14060 ^ _58993;
  wire _58995 = _58992 ^ _58994;
  wire _58996 = _15603 ^ _9718;
  wire _58997 = uncoded_block[101] ^ uncoded_block[109];
  wire _58998 = uncoded_block[110] ^ uncoded_block[116];
  wire _58999 = _58997 ^ _58998;
  wire _59000 = _58996 ^ _58999;
  wire _59001 = _58995 ^ _59000;
  wire _59002 = _58990 ^ _59001;
  wire _59003 = _2498 ^ _33058;
  wire _59004 = uncoded_block[128] ^ uncoded_block[133];
  wire _59005 = _59004 ^ _4760;
  wire _59006 = _59003 ^ _59005;
  wire _59007 = _58371 ^ _29208;
  wire _59008 = _41061 ^ _85;
  wire _59009 = _59007 ^ _59008;
  wire _59010 = _59006 ^ _59009;
  wire _59011 = uncoded_block[194] ^ uncoded_block[198];
  wire _59012 = _88 ^ _59011;
  wire _59013 = _10849 ^ _8021;
  wire _59014 = _59012 ^ _59013;
  wire _59015 = uncoded_block[214] ^ uncoded_block[223];
  wire _59016 = _7415 ^ _59015;
  wire _59017 = _2545 ^ _25104;
  wire _59018 = _59016 ^ _59017;
  wire _59019 = _59014 ^ _59018;
  wire _59020 = _59010 ^ _59019;
  wire _59021 = _59002 ^ _59020;
  wire _59022 = _4800 ^ _1786;
  wire _59023 = _120 ^ _3321;
  wire _59024 = _59022 ^ _59023;
  wire _59025 = _4814 ^ _1803;
  wire _59026 = uncoded_block[289] ^ uncoded_block[295];
  wire _59027 = _59026 ^ _8051;
  wire _59028 = _59025 ^ _59027;
  wire _59029 = _59024 ^ _59028;
  wire _59030 = uncoded_block[305] ^ uncoded_block[315];
  wire _59031 = _59030 ^ _2580;
  wire _59032 = _13081 ^ _2587;
  wire _59033 = _59031 ^ _59032;
  wire _59034 = _46597 ^ _16161;
  wire _59035 = uncoded_block[350] ^ uncoded_block[354];
  wire _59036 = _59035 ^ _23330;
  wire _59037 = _59034 ^ _59036;
  wire _59038 = _59033 ^ _59037;
  wire _59039 = _59029 ^ _59038;
  wire _59040 = _17658 ^ _4141;
  wire _59041 = uncoded_block[382] ^ uncoded_block[393];
  wire _59042 = _59041 ^ _1847;
  wire _59043 = _59040 ^ _59042;
  wire _59044 = uncoded_block[404] ^ uncoded_block[418];
  wire _59045 = _10341 ^ _59044;
  wire _59046 = uncoded_block[422] ^ uncoded_block[433];
  wire _59047 = _59046 ^ _2640;
  wire _59048 = _59045 ^ _59047;
  wire _59049 = _59043 ^ _59048;
  wire _59050 = _16187 ^ _21974;
  wire _59051 = _9275 ^ _6900;
  wire _59052 = _59050 ^ _59051;
  wire _59053 = uncoded_block[458] ^ uncoded_block[473];
  wire _59054 = _1870 ^ _59053;
  wire _59055 = _4189 ^ _9832;
  wire _59056 = _59054 ^ _59055;
  wire _59057 = _59052 ^ _59056;
  wire _59058 = _59049 ^ _59057;
  wire _59059 = _59039 ^ _59058;
  wire _59060 = _59021 ^ _59059;
  wire _59061 = uncoded_block[496] ^ uncoded_block[502];
  wire _59062 = uncoded_block[505] ^ uncoded_block[517];
  wire _59063 = _59061 ^ _59062;
  wire _59064 = uncoded_block[525] ^ uncoded_block[533];
  wire _59065 = _9841 ^ _59064;
  wire _59066 = _59063 ^ _59065;
  wire _59067 = _1115 ^ _28882;
  wire _59068 = uncoded_block[546] ^ uncoded_block[551];
  wire _59069 = _59068 ^ _4934;
  wire _59070 = _59067 ^ _59069;
  wire _59071 = _59066 ^ _59070;
  wire _59072 = uncoded_block[573] ^ uncoded_block[581];
  wire _59073 = _18682 ^ _59072;
  wire _59074 = _22012 ^ _34013;
  wire _59075 = _59073 ^ _59074;
  wire _59076 = uncoded_block[606] ^ uncoded_block[614];
  wire _59077 = _41941 ^ _59076;
  wire _59078 = _13713 ^ _6331;
  wire _59079 = _59077 ^ _59078;
  wire _59080 = _59075 ^ _59079;
  wire _59081 = _59071 ^ _59080;
  wire _59082 = _3502 ^ _297;
  wire _59083 = _302 ^ _16747;
  wire _59084 = _59082 ^ _59083;
  wire _59085 = _57381 ^ _50508;
  wire _59086 = _59084 ^ _59085;
  wire _59087 = _22963 ^ _322;
  wire _59088 = _4272 ^ _34840;
  wire _59089 = _59087 ^ _59088;
  wire _59090 = uncoded_block[734] ^ uncoded_block[742];
  wire _59091 = _36036 ^ _59090;
  wire _59092 = _7013 ^ _43417;
  wire _59093 = _59091 ^ _59092;
  wire _59094 = _59089 ^ _59093;
  wire _59095 = _59086 ^ _59094;
  wire _59096 = _59081 ^ _59095;
  wire _59097 = _11019 ^ _12117;
  wire _59098 = _59097 ^ _48582;
  wire _59099 = _34059 ^ _57406;
  wire _59100 = uncoded_block[814] ^ uncoded_block[821];
  wire _59101 = _8793 ^ _59100;
  wire _59102 = _59099 ^ _59101;
  wire _59103 = _59098 ^ _59102;
  wire _59104 = _17797 ^ _1250;
  wire _59105 = uncoded_block[854] ^ uncoded_block[864];
  wire _59106 = _1253 ^ _59105;
  wire _59107 = _59104 ^ _59106;
  wire _59108 = uncoded_block[871] ^ uncoded_block[882];
  wire _59109 = _16811 ^ _59108;
  wire _59110 = uncoded_block[886] ^ uncoded_block[897];
  wire _59111 = _59110 ^ _49819;
  wire _59112 = _59109 ^ _59111;
  wire _59113 = _59107 ^ _59112;
  wire _59114 = _59103 ^ _59113;
  wire _59115 = _435 ^ _3631;
  wire _59116 = _31995 ^ _16321;
  wire _59117 = _59115 ^ _59116;
  wire _59118 = uncoded_block[941] ^ uncoded_block[949];
  wire _59119 = _24383 ^ _59118;
  wire _59120 = _4381 ^ _45753;
  wire _59121 = _59119 ^ _59120;
  wire _59122 = _59117 ^ _59121;
  wire _59123 = _1310 ^ _11087;
  wire _59124 = uncoded_block[969] ^ uncoded_block[974];
  wire _59125 = _59124 ^ _57438;
  wire _59126 = _59123 ^ _59125;
  wire _59127 = uncoded_block[993] ^ uncoded_block[1004];
  wire _59128 = _59127 ^ _43085;
  wire _59129 = uncoded_block[1012] ^ uncoded_block[1019];
  wire _59130 = _59129 ^ _4415;
  wire _59131 = _59128 ^ _59130;
  wire _59132 = _59126 ^ _59131;
  wire _59133 = _59122 ^ _59132;
  wire _59134 = _59114 ^ _59133;
  wire _59135 = _59096 ^ _59134;
  wire _59136 = _59060 ^ _59135;
  wire _59137 = _31172 ^ _50575;
  wire _59138 = uncoded_block[1049] ^ uncoded_block[1058];
  wire _59139 = _6475 ^ _59138;
  wire _59140 = _59137 ^ _59139;
  wire _59141 = _42044 ^ _12213;
  wire _59142 = uncoded_block[1071] ^ uncoded_block[1082];
  wire _59143 = _59142 ^ _5839;
  wire _59144 = _59141 ^ _59143;
  wire _59145 = _59140 ^ _59144;
  wire _59146 = _58874 ^ _16370;
  wire _59147 = _550 ^ _25323;
  wire _59148 = _1388 ^ _57152;
  wire _59149 = _59147 ^ _59148;
  wire _59150 = _59146 ^ _59149;
  wire _59151 = _59145 ^ _59150;
  wire _59152 = uncoded_block[1129] ^ uncoded_block[1151];
  wire _59153 = _59152 ^ _4469;
  wire _59154 = uncoded_block[1165] ^ uncoded_block[1181];
  wire _59155 = _7149 ^ _59154;
  wire _59156 = _59153 ^ _59155;
  wire _59157 = uncoded_block[1182] ^ uncoded_block[1189];
  wire _59158 = _59157 ^ _5207;
  wire _59159 = uncoded_block[1206] ^ uncoded_block[1212];
  wire _59160 = uncoded_block[1213] ^ uncoded_block[1220];
  wire _59161 = _59159 ^ _59160;
  wire _59162 = _59158 ^ _59161;
  wire _59163 = _59156 ^ _59162;
  wire _59164 = uncoded_block[1227] ^ uncoded_block[1233];
  wire _59165 = _45036 ^ _59164;
  wire _59166 = _3772 ^ _16408;
  wire _59167 = _59165 ^ _59166;
  wire _59168 = uncoded_block[1246] ^ uncoded_block[1253];
  wire _59169 = _59168 ^ _56573;
  wire _59170 = _5235 ^ _58902;
  wire _59171 = _59169 ^ _59170;
  wire _59172 = _59167 ^ _59171;
  wire _59173 = _59163 ^ _59172;
  wire _59174 = _59151 ^ _59173;
  wire _59175 = _11194 ^ _57502;
  wire _59176 = uncoded_block[1292] ^ uncoded_block[1301];
  wire _59177 = _59176 ^ _11759;
  wire _59178 = uncoded_block[1322] ^ uncoded_block[1327];
  wire _59179 = uncoded_block[1335] ^ uncoded_block[1340];
  wire _59180 = _59178 ^ _59179;
  wire _59181 = _59177 ^ _59180;
  wire _59182 = _59175 ^ _59181;
  wire _59183 = uncoded_block[1341] ^ uncoded_block[1347];
  wire _59184 = _59183 ^ _57518;
  wire _59185 = uncoded_block[1357] ^ uncoded_block[1363];
  wire _59186 = _59185 ^ _40581;
  wire _59187 = _59184 ^ _59186;
  wire _59188 = _680 ^ _15966;
  wire _59189 = uncoded_block[1386] ^ uncoded_block[1390];
  wire _59190 = _7219 ^ _59189;
  wire _59191 = _59188 ^ _59190;
  wire _59192 = _59187 ^ _59191;
  wire _59193 = _59182 ^ _59192;
  wire _59194 = _7834 ^ _1517;
  wire _59195 = _5294 ^ _33374;
  wire _59196 = _59194 ^ _59195;
  wire _59197 = _9021 ^ _9588;
  wire _59198 = _21323 ^ _15982;
  wire _59199 = _59197 ^ _59198;
  wire _59200 = _59196 ^ _59199;
  wire _59201 = uncoded_block[1448] ^ uncoded_block[1456];
  wire _59202 = _45085 ^ _59201;
  wire _59203 = _36213 ^ _3094;
  wire _59204 = _59202 ^ _59203;
  wire _59205 = _3879 ^ _3881;
  wire _59206 = uncoded_block[1490] ^ uncoded_block[1496];
  wire _59207 = _3884 ^ _59206;
  wire _59208 = _59205 ^ _59207;
  wire _59209 = _59204 ^ _59208;
  wire _59210 = _59200 ^ _59209;
  wire _59211 = _59193 ^ _59210;
  wire _59212 = _59174 ^ _59211;
  wire _59213 = _7259 ^ _4617;
  wire _59214 = _37053 ^ _59213;
  wire _59215 = _751 ^ _46860;
  wire _59216 = _4623 ^ _6647;
  wire _59217 = _59215 ^ _59216;
  wire _59218 = _59214 ^ _59217;
  wire _59219 = _16496 ^ _27626;
  wire _59220 = uncoded_block[1556] ^ uncoded_block[1562];
  wire _59221 = _50336 ^ _59220;
  wire _59222 = _59219 ^ _59221;
  wire _59223 = _32565 ^ _16515;
  wire _59224 = _11292 ^ _14517;
  wire _59225 = _59223 ^ _59224;
  wire _59226 = _59222 ^ _59225;
  wire _59227 = _59218 ^ _59226;
  wire _59228 = uncoded_block[1617] ^ uncoded_block[1624];
  wire _59229 = _16031 ^ _59228;
  wire _59230 = _807 ^ _3166;
  wire _59231 = _59229 ^ _59230;
  wire _59232 = uncoded_block[1635] ^ uncoded_block[1639];
  wire _59233 = uncoded_block[1641] ^ uncoded_block[1648];
  wire _59234 = _59232 ^ _59233;
  wire _59235 = _3953 ^ _820;
  wire _59236 = _59234 ^ _59235;
  wire _59237 = _59231 ^ _59236;
  wire _59238 = uncoded_block[1687] ^ uncoded_block[1693];
  wire _59239 = _11321 ^ _59238;
  wire _59240 = _57578 ^ _59239;
  wire _59241 = _2430 ^ _1670;
  wire _59242 = _5412 ^ uncoded_block[1722];
  wire _59243 = _59241 ^ _59242;
  wire _59244 = _59240 ^ _59243;
  wire _59245 = _59237 ^ _59244;
  wire _59246 = _59227 ^ _59245;
  wire _59247 = _59212 ^ _59246;
  wire _59248 = _59136 ^ _59247;
  wire _59249 = uncoded_block[0] ^ uncoded_block[17];
  wire _59250 = _59249 ^ _3219;
  wire _59251 = _18 ^ _56408;
  wire _59252 = _59250 ^ _59251;
  wire _59253 = _56409 ^ _47675;
  wire _59254 = _9161 ^ _2484;
  wire _59255 = _59253 ^ _59254;
  wire _59256 = _59252 ^ _59255;
  wire _59257 = uncoded_block[116] ^ uncoded_block[124];
  wire _59258 = _1718 ^ _59257;
  wire _59259 = uncoded_block[133] ^ uncoded_block[142];
  wire _59260 = _59259 ^ _70;
  wire _59261 = _59258 ^ _59260;
  wire _59262 = _56421 ^ _56425;
  wire _59263 = _59261 ^ _59262;
  wire _59264 = _59256 ^ _59263;
  wire _59265 = uncoded_block[208] ^ uncoded_block[219];
  wire _59266 = _89 ^ _59265;
  wire _59267 = _50418 ^ _14116;
  wire _59268 = _59266 ^ _59267;
  wire _59269 = _59268 ^ _56441;
  wire _59270 = uncoded_block[294] ^ uncoded_block[316];
  wire _59271 = uncoded_block[324] ^ uncoded_block[331];
  wire _59272 = _59270 ^ _59271;
  wire _59273 = uncoded_block[345] ^ uncoded_block[351];
  wire _59274 = _56444 ^ _59273;
  wire _59275 = _59272 ^ _59274;
  wire _59276 = _50076 ^ _31862;
  wire _59277 = _59276 ^ _56453;
  wire _59278 = _59275 ^ _59277;
  wire _59279 = _59269 ^ _59278;
  wire _59280 = _59264 ^ _59279;
  wire _59281 = _32297 ^ _5577;
  wire _59282 = _56456 ^ _59281;
  wire _59283 = _56462 ^ _56464;
  wire _59284 = _5600 ^ _6919;
  wire _59285 = _59283 ^ _59284;
  wire _59286 = _59282 ^ _59285;
  wire _59287 = uncoded_block[499] ^ uncoded_block[530];
  wire _59288 = _59287 ^ _24279;
  wire _59289 = _56473 ^ _1916;
  wire _59290 = _59288 ^ _59289;
  wire _59291 = _8139 ^ _52447;
  wire _59292 = _26096 ^ _4236;
  wire _59293 = _59291 ^ _59292;
  wire _59294 = _59290 ^ _59293;
  wire _59295 = _59286 ^ _59294;
  wire _59296 = uncoded_block[606] ^ uncoded_block[624];
  wire _59297 = _11535 ^ _59296;
  wire _59298 = _59297 ^ _56485;
  wire _59299 = uncoded_block[648] ^ uncoded_block[655];
  wire _59300 = _16241 ^ _59299;
  wire _59301 = _15270 ^ _56495;
  wire _59302 = _59300 ^ _59301;
  wire _59303 = _59298 ^ _59302;
  wire _59304 = uncoded_block[693] ^ uncoded_block[713];
  wire _59305 = _59304 ^ _38450;
  wire _59306 = _2768 ^ _9908;
  wire _59307 = _59305 ^ _59306;
  wire _59308 = uncoded_block[750] ^ uncoded_block[760];
  wire _59309 = _5013 ^ _59308;
  wire _59310 = _17776 ^ _56505;
  wire _59311 = _59309 ^ _59310;
  wire _59312 = _59307 ^ _59311;
  wire _59313 = _59303 ^ _59312;
  wire _59314 = _59295 ^ _59313;
  wire _59315 = _59280 ^ _59314;
  wire _59316 = uncoded_block[801] ^ uncoded_block[809];
  wire _59317 = _56506 ^ _59316;
  wire _59318 = uncoded_block[811] ^ uncoded_block[820];
  wire _59319 = _59318 ^ _400;
  wire _59320 = _59317 ^ _59319;
  wire _59321 = uncoded_block[838] ^ uncoded_block[862];
  wire _59322 = _401 ^ _59321;
  wire _59323 = _59322 ^ _56519;
  wire _59324 = _59320 ^ _59323;
  wire _59325 = _5762 ^ _56521;
  wire _59326 = _27049 ^ _59325;
  wire _59327 = uncoded_block[946] ^ uncoded_block[956];
  wire _59328 = _2083 ^ _59327;
  wire _59329 = _12179 ^ _5786;
  wire _59330 = _59328 ^ _59329;
  wire _59331 = _59326 ^ _59330;
  wire _59332 = _59324 ^ _59331;
  wire _59333 = _28980 ^ _56532;
  wire _59334 = _1326 ^ _5129;
  wire _59335 = _59333 ^ _59334;
  wire _59336 = _19286 ^ _2127;
  wire _59337 = uncoded_block[1043] ^ uncoded_block[1046];
  wire _59338 = _59337 ^ _42039;
  wire _59339 = _59336 ^ _59338;
  wire _59340 = _59335 ^ _59339;
  wire _59341 = _22603 ^ _2924;
  wire _59342 = _59341 ^ _56550;
  wire _59343 = _44259 ^ _9484;
  wire _59344 = uncoded_block[1125] ^ uncoded_block[1145];
  wire _59345 = _45790 ^ _59344;
  wire _59346 = _59343 ^ _59345;
  wire _59347 = _59342 ^ _59346;
  wire _59348 = _59340 ^ _59347;
  wire _59349 = _59332 ^ _59348;
  wire _59350 = _5866 ^ _2188;
  wire _59351 = uncoded_block[1170] ^ uncoded_block[1187];
  wire _59352 = _5869 ^ _59351;
  wire _59353 = _59350 ^ _59352;
  wire _59354 = _5882 ^ _1425;
  wire _59355 = _36581 ^ _5218;
  wire _59356 = _59354 ^ _59355;
  wire _59357 = _59353 ^ _59356;
  wire _59358 = _15441 ^ _10630;
  wire _59359 = _21732 ^ _56574;
  wire _59360 = _59358 ^ _59359;
  wire _59361 = uncoded_block[1283] ^ uncoded_block[1298];
  wire _59362 = _3011 ^ _59361;
  wire _59363 = uncoded_block[1303] ^ uncoded_block[1324];
  wire _59364 = _18870 ^ _59363;
  wire _59365 = _59362 ^ _59364;
  wire _59366 = _59360 ^ _59365;
  wire _59367 = _59357 ^ _59366;
  wire _59368 = _56585 ^ _5272;
  wire _59369 = _59368 ^ _56591;
  wire _59370 = _59369 ^ _56598;
  wire _59371 = _29508 ^ _717;
  wire _59372 = _59371 ^ _25868;
  wire _59373 = _4601 ^ _9610;
  wire _59374 = _1558 ^ _8461;
  wire _59375 = _59373 ^ _59374;
  wire _59376 = _59372 ^ _59375;
  wire _59377 = _59370 ^ _59376;
  wire _59378 = _59367 ^ _59377;
  wire _59379 = _59349 ^ _59378;
  wire _59380 = _59315 ^ _59379;
  wire _59381 = uncoded_block[1490] ^ uncoded_block[1498];
  wire _59382 = _59381 ^ _1575;
  wire _59383 = _15004 ^ _1582;
  wire _59384 = _59382 ^ _59383;
  wire _59385 = _56612 ^ _56615;
  wire _59386 = _59384 ^ _59385;
  wire _59387 = uncoded_block[1583] ^ uncoded_block[1592];
  wire _59388 = _59387 ^ _13486;
  wire _59389 = uncoded_block[1599] ^ uncoded_block[1603];
  wire _59390 = _59389 ^ _5382;
  wire _59391 = _59388 ^ _59390;
  wire _59392 = uncoded_block[1621] ^ uncoded_block[1625];
  wire _59393 = _59392 ^ _56625;
  wire _59394 = _56626 ^ _56628;
  wire _59395 = _59393 ^ _59394;
  wire _59396 = _59391 ^ _59395;
  wire _59397 = _59386 ^ _59396;
  wire _59398 = _3967 ^ _11327;
  wire _59399 = _59398 ^ uncoded_block[1714];
  wire _59400 = _59397 ^ _59399;
  wire _59401 = _59380 ^ _59400;
  wire _59402 = uncoded_block[0] ^ uncoded_block[7];
  wire _59403 = uncoded_block[8] ^ uncoded_block[18];
  wire _59404 = _59402 ^ _59403;
  wire _59405 = _2458 ^ _14565;
  wire _59406 = _59404 ^ _59405;
  wire _59407 = _1693 ^ _16;
  wire _59408 = _7965 ^ _10234;
  wire _59409 = _59407 ^ _59408;
  wire _59410 = _59406 ^ _59409;
  wire _59411 = _14575 ^ _19506;
  wire _59412 = _23698 ^ _12438;
  wire _59413 = _59411 ^ _59412;
  wire _59414 = uncoded_block[85] ^ uncoded_block[98];
  wire _59415 = _6750 ^ _59414;
  wire _59416 = uncoded_block[101] ^ uncoded_block[106];
  wire _59417 = _59416 ^ _54596;
  wire _59418 = _59415 ^ _59417;
  wire _59419 = _59413 ^ _59418;
  wire _59420 = _59410 ^ _59419;
  wire _59421 = _4040 ^ _18567;
  wire _59422 = _7999 ^ _13573;
  wire _59423 = _59421 ^ _59422;
  wire _59424 = uncoded_block[153] ^ uncoded_block[165];
  wire _59425 = _59424 ^ _81;
  wire _59426 = _4057 ^ _7403;
  wire _59427 = _59425 ^ _59426;
  wire _59428 = _59423 ^ _59427;
  wire _59429 = _8018 ^ _4779;
  wire _59430 = _25092 ^ _59429;
  wire _59431 = uncoded_block[213] ^ uncoded_block[222];
  wire _59432 = _59431 ^ _4076;
  wire _59433 = _3299 ^ _29225;
  wire _59434 = _59432 ^ _59433;
  wire _59435 = _59430 ^ _59434;
  wire _59436 = _59428 ^ _59435;
  wire _59437 = _59420 ^ _59436;
  wire _59438 = _968 ^ _10860;
  wire _59439 = _116 ^ _3311;
  wire _59440 = _59438 ^ _59439;
  wire _59441 = uncoded_block[272] ^ uncoded_block[277];
  wire _59442 = _3312 ^ _59441;
  wire _59443 = _41876 ^ _11428;
  wire _59444 = _59442 ^ _59443;
  wire _59445 = _59440 ^ _59444;
  wire _59446 = _995 ^ _1000;
  wire _59447 = _25569 ^ _23764;
  wire _59448 = _59446 ^ _59447;
  wire _59449 = _29663 ^ _41885;
  wire _59450 = uncoded_block[339] ^ uncoded_block[347];
  wire _59451 = _1822 ^ _59450;
  wire _59452 = _59449 ^ _59451;
  wire _59453 = _59448 ^ _59452;
  wire _59454 = _59445 ^ _59453;
  wire _59455 = uncoded_block[355] ^ uncoded_block[367];
  wire _59456 = _17651 ^ _59455;
  wire _59457 = _59456 ^ _50798;
  wire _59458 = _33962 ^ _4151;
  wire _59459 = _10340 ^ _7487;
  wire _59460 = _59458 ^ _59459;
  wire _59461 = _59457 ^ _59460;
  wire _59462 = _5565 ^ _3397;
  wire _59463 = _35576 ^ _14690;
  wire _59464 = _59462 ^ _59463;
  wire _59465 = _21974 ^ _10356;
  wire _59466 = uncoded_block[453] ^ uncoded_block[459];
  wire _59467 = _59466 ^ _12023;
  wire _59468 = _59465 ^ _59467;
  wire _59469 = _59464 ^ _59468;
  wire _59470 = _59461 ^ _59469;
  wire _59471 = _59454 ^ _59470;
  wire _59472 = _59437 ^ _59471;
  wire _59473 = uncoded_block[476] ^ uncoded_block[484];
  wire _59474 = _59473 ^ _6276;
  wire _59475 = _1093 ^ _21536;
  wire _59476 = _59474 ^ _59475;
  wire _59477 = _12034 ^ _10945;
  wire _59478 = _59477 ^ _12038;
  wire _59479 = _59476 ^ _59478;
  wire _59480 = _1117 ^ _23382;
  wire _59481 = _59480 ^ _8138;
  wire _59482 = uncoded_block[562] ^ uncoded_block[567];
  wire _59483 = _59482 ^ _39617;
  wire _59484 = _263 ^ _6947;
  wire _59485 = _59483 ^ _59484;
  wire _59486 = _59481 ^ _59485;
  wire _59487 = _59479 ^ _59486;
  wire _59488 = _52450 ^ _8148;
  wire _59489 = uncoded_block[597] ^ uncoded_block[603];
  wire _59490 = _59489 ^ _39233;
  wire _59491 = _59488 ^ _59490;
  wire _59492 = _51584 ^ _4964;
  wire _59493 = _36847 ^ _3502;
  wire _59494 = _59492 ^ _59493;
  wire _59495 = _59491 ^ _59494;
  wire _59496 = _2729 ^ _41955;
  wire _59497 = _57071 ^ _21113;
  wire _59498 = _59496 ^ _59497;
  wire _59499 = _4265 ^ _17745;
  wire _59500 = _319 ^ _31076;
  wire _59501 = _59499 ^ _59500;
  wire _59502 = _59498 ^ _59501;
  wire _59503 = _59495 ^ _59502;
  wire _59504 = _59487 ^ _59503;
  wire _59505 = uncoded_block[704] ^ uncoded_block[710];
  wire _59506 = _1186 ^ _59505;
  wire _59507 = _5002 ^ _44171;
  wire _59508 = _59506 ^ _59507;
  wire _59509 = uncoded_block[727] ^ uncoded_block[738];
  wire _59510 = _1988 ^ _59509;
  wire _59511 = uncoded_block[748] ^ uncoded_block[755];
  wire _59512 = _23870 ^ _59511;
  wire _59513 = _59510 ^ _59512;
  wire _59514 = _59508 ^ _59513;
  wire _59515 = _4298 ^ _2006;
  wire _59516 = uncoded_block[766] ^ uncoded_block[780];
  wire _59517 = _59516 ^ _3570;
  wire _59518 = _59515 ^ _59517;
  wire _59519 = uncoded_block[791] ^ uncoded_block[806];
  wire _59520 = _4311 ^ _59519;
  wire _59521 = _1238 ^ _57408;
  wire _59522 = _59520 ^ _59521;
  wire _59523 = _59518 ^ _59522;
  wire _59524 = _59514 ^ _59523;
  wire _59525 = _52500 ^ _10490;
  wire _59526 = uncoded_block[841] ^ uncoded_block[847];
  wire _59527 = _4336 ^ _59526;
  wire _59528 = _59525 ^ _59527;
  wire _59529 = _1262 ^ _57922;
  wire _59530 = uncoded_block[890] ^ uncoded_block[897];
  wire _59531 = _43820 ^ _59530;
  wire _59532 = _59529 ^ _59531;
  wire _59533 = _59528 ^ _59532;
  wire _59534 = _3617 ^ _10508;
  wire _59535 = _59534 ^ _37717;
  wire _59536 = uncoded_block[922] ^ uncoded_block[939];
  wire _59537 = _3629 ^ _59536;
  wire _59538 = _13263 ^ _9975;
  wire _59539 = _59537 ^ _59538;
  wire _59540 = _59535 ^ _59539;
  wire _59541 = _59533 ^ _59540;
  wire _59542 = _59524 ^ _59541;
  wire _59543 = _59504 ^ _59542;
  wire _59544 = _59472 ^ _59543;
  wire _59545 = uncoded_block[959] ^ uncoded_block[973];
  wire _59546 = _57120 ^ _59545;
  wire _59547 = _43842 ^ _7689;
  wire _59548 = _59546 ^ _59547;
  wire _59549 = _1318 ^ _38123;
  wire _59550 = uncoded_block[1003] ^ uncoded_block[1017];
  wire _59551 = _2111 ^ _59550;
  wire _59552 = _59549 ^ _59551;
  wire _59553 = _59548 ^ _59552;
  wire _59554 = _7108 ^ _498;
  wire _59555 = uncoded_block[1042] ^ uncoded_block[1048];
  wire _59556 = _9459 ^ _59555;
  wire _59557 = _59554 ^ _59556;
  wire _59558 = _10564 ^ _1360;
  wire _59559 = _10566 ^ _5826;
  wire _59560 = _59558 ^ _59559;
  wire _59561 = _59557 ^ _59560;
  wire _59562 = _59553 ^ _59561;
  wire _59563 = _34934 ^ _20251;
  wire _59564 = uncoded_block[1089] ^ uncoded_block[1094];
  wire _59565 = _42054 ^ _59564;
  wire _59566 = _59563 ^ _59565;
  wire _59567 = uncoded_block[1106] ^ uncoded_block[1115];
  wire _59568 = _4444 ^ _59567;
  wire _59569 = uncoded_block[1132] ^ uncoded_block[1138];
  wire _59570 = _7736 ^ _59569;
  wire _59571 = _59568 ^ _59570;
  wire _59572 = _59566 ^ _59571;
  wire _59573 = uncoded_block[1149] ^ uncoded_block[1155];
  wire _59574 = _25790 ^ _59573;
  wire _59575 = _43875 ^ _3740;
  wire _59576 = _59574 ^ _59575;
  wire _59577 = _10608 ^ _35354;
  wire _59578 = uncoded_block[1190] ^ uncoded_block[1197];
  wire _59579 = _59578 ^ _17400;
  wire _59580 = _59577 ^ _59579;
  wire _59581 = _59576 ^ _59580;
  wire _59582 = _59572 ^ _59581;
  wire _59583 = _59562 ^ _59582;
  wire _59584 = _6529 ^ _1427;
  wire _59585 = _1432 ^ _13355;
  wire _59586 = _59584 ^ _59585;
  wire _59587 = uncoded_block[1232] ^ uncoded_block[1248];
  wire _59588 = uncoded_block[1255] ^ uncoded_block[1262];
  wire _59589 = _59587 ^ _59588;
  wire _59590 = _7770 ^ _59589;
  wire _59591 = _59586 ^ _59590;
  wire _59592 = uncoded_block[1274] ^ uncoded_block[1289];
  wire _59593 = _6550 ^ _59592;
  wire _59594 = uncoded_block[1305] ^ uncoded_block[1317];
  wire _59595 = _55370 ^ _59594;
  wire _59596 = _59593 ^ _59595;
  wire _59597 = _47945 ^ _44316;
  wire _59598 = uncoded_block[1340] ^ uncoded_block[1357];
  wire _59599 = _5259 ^ _59598;
  wire _59600 = _59597 ^ _59599;
  wire _59601 = _59596 ^ _59600;
  wire _59602 = _59591 ^ _59601;
  wire _59603 = _2283 ^ _54880;
  wire _59604 = _36191 ^ _59603;
  wire _59605 = uncoded_block[1373] ^ uncoded_block[1380];
  wire _59606 = uncoded_block[1386] ^ uncoded_block[1392];
  wire _59607 = _59605 ^ _59606;
  wire _59608 = _5955 ^ _3846;
  wire _59609 = _59607 ^ _59608;
  wire _59610 = _59604 ^ _59609;
  wire _59611 = _2300 ^ _1523;
  wire _59612 = uncoded_block[1414] ^ uncoded_block[1419];
  wire _59613 = _59612 ^ _29095;
  wire _59614 = _59611 ^ _59613;
  wire _59615 = uncoded_block[1430] ^ uncoded_block[1436];
  wire _59616 = _59615 ^ _26763;
  wire _59617 = uncoded_block[1455] ^ uncoded_block[1462];
  wire _59618 = _59617 ^ _14989;
  wire _59619 = _59616 ^ _59618;
  wire _59620 = _59614 ^ _59619;
  wire _59621 = _59610 ^ _59620;
  wire _59622 = _59602 ^ _59621;
  wire _59623 = _59583 ^ _59622;
  wire _59624 = uncoded_block[1494] ^ uncoded_block[1499];
  wire _59625 = _49448 ^ _59624;
  wire _59626 = uncoded_block[1508] ^ uncoded_block[1516];
  wire _59627 = _11813 ^ _59626;
  wire _59628 = _59625 ^ _59627;
  wire _59629 = _754 ^ _11270;
  wire _59630 = _5344 ^ _3905;
  wire _59631 = _59629 ^ _59630;
  wire _59632 = _59628 ^ _59631;
  wire _59633 = uncoded_block[1540] ^ uncoded_block[1545];
  wire _59634 = uncoded_block[1546] ^ uncoded_block[1554];
  wire _59635 = _59633 ^ _59634;
  wire _59636 = uncoded_block[1568] ^ uncoded_block[1578];
  wire _59637 = _13991 ^ _59636;
  wire _59638 = _59635 ^ _59637;
  wire _59639 = _784 ^ _56938;
  wire _59640 = _6673 ^ _8499;
  wire _59641 = _59639 ^ _59640;
  wire _59642 = _59638 ^ _59641;
  wire _59643 = _59632 ^ _59642;
  wire _59644 = _1624 ^ _2396;
  wire _59645 = _3937 ^ _804;
  wire _59646 = _59644 ^ _59645;
  wire _59647 = _59392 ^ _6048;
  wire _59648 = _59647 ^ _43237;
  wire _59649 = _59646 ^ _59648;
  wire _59650 = uncoded_block[1652] ^ uncoded_block[1660];
  wire _59651 = _59650 ^ _22761;
  wire _59652 = uncoded_block[1667] ^ uncoded_block[1678];
  wire _59653 = _59652 ^ _23671;
  wire _59654 = _59651 ^ _59653;
  wire _59655 = _6705 ^ _6066;
  wire _59656 = _1669 ^ _35477;
  wire _59657 = _59655 ^ _59656;
  wire _59658 = _59654 ^ _59657;
  wire _59659 = _59649 ^ _59658;
  wire _59660 = _59643 ^ _59659;
  wire _59661 = _16064 ^ uncoded_block[1718];
  wire _59662 = _59660 ^ _59661;
  wire _59663 = _59623 ^ _59662;
  wire _59664 = _59544 ^ _59663;
  wire _59665 = _10787 ^ _55821;
  wire _59666 = _17060 ^ _25941;
  wire _59667 = _59665 ^ _59666;
  wire _59668 = _58050 ^ _7966;
  wire _59669 = _33467 ^ _19019;
  wire _59670 = _59668 ^ _59669;
  wire _59671 = _59667 ^ _59670;
  wire _59672 = _2487 ^ _4741;
  wire _59673 = _6116 ^ _13011;
  wire _59674 = _59672 ^ _59673;
  wire _59675 = _6128 ^ _42875;
  wire _59676 = _64 ^ _6138;
  wire _59677 = _59675 ^ _59676;
  wire _59678 = _59674 ^ _59677;
  wire _59679 = _59671 ^ _59678;
  wire _59680 = _4047 ^ _10835;
  wire _59681 = uncoded_block[163] ^ uncoded_block[170];
  wire _59682 = uncoded_block[177] ^ uncoded_block[186];
  wire _59683 = _59681 ^ _59682;
  wire _59684 = _2529 ^ _9744;
  wire _59685 = _59683 ^ _59684;
  wire _59686 = _59680 ^ _59685;
  wire _59687 = _95 ^ _30963;
  wire _59688 = uncoded_block[212] ^ uncoded_block[218];
  wire _59689 = _59688 ^ _4076;
  wire _59690 = _59687 ^ _59689;
  wire _59691 = uncoded_block[231] ^ uncoded_block[235];
  wire _59692 = _11945 ^ _59691;
  wire _59693 = _4084 ^ _14116;
  wire _59694 = _59692 ^ _59693;
  wire _59695 = _59690 ^ _59694;
  wire _59696 = _59686 ^ _59695;
  wire _59697 = _59679 ^ _59696;
  wire _59698 = _31834 ^ _26441;
  wire _59699 = _18600 ^ _10303;
  wire _59700 = _59698 ^ _59699;
  wire _59701 = _5515 ^ _29238;
  wire _59702 = uncoded_block[302] ^ uncoded_block[309];
  wire _59703 = _2573 ^ _59702;
  wire _59704 = _59701 ^ _59703;
  wire _59705 = _59700 ^ _59704;
  wire _59706 = uncoded_block[320] ^ uncoded_block[325];
  wire _59707 = _59706 ^ _13081;
  wire _59708 = _1017 ^ _37186;
  wire _59709 = _59707 ^ _59708;
  wire _59710 = uncoded_block[352] ^ uncoded_block[375];
  wire _59711 = _8652 ^ _59710;
  wire _59712 = uncoded_block[394] ^ uncoded_block[399];
  wire _59713 = _59712 ^ _6244;
  wire _59714 = _59711 ^ _59713;
  wire _59715 = _59709 ^ _59714;
  wire _59716 = _59705 ^ _59715;
  wire _59717 = uncoded_block[412] ^ uncoded_block[421];
  wire _59718 = _59717 ^ _24248;
  wire _59719 = _14689 ^ _1067;
  wire _59720 = _59718 ^ _59719;
  wire _59721 = _9275 ^ _4177;
  wire _59722 = uncoded_block[460] ^ uncoded_block[467];
  wire _59723 = _59722 ^ _3418;
  wire _59724 = _59721 ^ _59723;
  wire _59725 = _59720 ^ _59724;
  wire _59726 = uncoded_block[475] ^ uncoded_block[483];
  wire _59727 = _59726 ^ _8694;
  wire _59728 = uncoded_block[488] ^ uncoded_block[493];
  wire _59729 = _59728 ^ _4195;
  wire _59730 = _59727 ^ _59729;
  wire _59731 = _6921 ^ _231;
  wire _59732 = uncoded_block[519] ^ uncoded_block[525];
  wire _59733 = _8705 ^ _59732;
  wire _59734 = _59731 ^ _59733;
  wire _59735 = _59730 ^ _59734;
  wire _59736 = _59725 ^ _59735;
  wire _59737 = _59716 ^ _59736;
  wire _59738 = _59697 ^ _59737;
  wire _59739 = _1900 ^ _16215;
  wire _59740 = uncoded_block[535] ^ uncoded_block[544];
  wire _59741 = _59740 ^ _35996;
  wire _59742 = _59739 ^ _59741;
  wire _59743 = _24284 ^ _31490;
  wire _59744 = uncoded_block[575] ^ uncoded_block[580];
  wire _59745 = uncoded_block[584] ^ uncoded_block[595];
  wire _59746 = _59744 ^ _59745;
  wire _59747 = _59743 ^ _59746;
  wire _59748 = _59742 ^ _59747;
  wire _59749 = _274 ^ _20626;
  wire _59750 = _8745 ^ _17238;
  wire _59751 = _59749 ^ _59750;
  wire _59752 = uncoded_block[638] ^ uncoded_block[642];
  wire _59753 = _59752 ^ _10425;
  wire _59754 = _59753 ^ _43396;
  wire _59755 = _59751 ^ _59754;
  wire _59756 = _59748 ^ _59755;
  wire _59757 = _51249 ^ _19185;
  wire _59758 = _8179 ^ _1972;
  wire _59759 = _59757 ^ _59758;
  wire _59760 = _325 ^ _12092;
  wire _59761 = _14766 ^ _14255;
  wire _59762 = _59760 ^ _59761;
  wire _59763 = _59759 ^ _59762;
  wire _59764 = uncoded_block[720] ^ uncoded_block[726];
  wire _59765 = _8190 ^ _59764;
  wire _59766 = _1995 ^ _20156;
  wire _59767 = _59765 ^ _59766;
  wire _59768 = uncoded_block[743] ^ uncoded_block[747];
  wire _59769 = _59768 ^ _4298;
  wire _59770 = _24796 ^ _7616;
  wire _59771 = _59769 ^ _59770;
  wire _59772 = _59767 ^ _59771;
  wire _59773 = _59763 ^ _59772;
  wire _59774 = _59756 ^ _59773;
  wire _59775 = _8213 ^ _9384;
  wire _59776 = uncoded_block[783] ^ uncoded_block[789];
  wire _59777 = _59776 ^ _5723;
  wire _59778 = _59775 ^ _59777;
  wire _59779 = _5042 ^ _7634;
  wire _59780 = _41215 ^ _59779;
  wire _59781 = _59778 ^ _59780;
  wire _59782 = uncoded_block[833] ^ uncoded_block[842];
  wire _59783 = _59782 ^ _1257;
  wire _59784 = uncoded_block[852] ^ uncoded_block[860];
  wire _59785 = _14814 ^ _59784;
  wire _59786 = _59783 ^ _59785;
  wire _59787 = _9416 ^ _44603;
  wire _59788 = _5750 ^ _59787;
  wire _59789 = _59786 ^ _59788;
  wire _59790 = _59781 ^ _59789;
  wire _59791 = _58199 ^ _2070;
  wire _59792 = _27463 ^ _3629;
  wire _59793 = _59791 ^ _59792;
  wire _59794 = _2073 ^ _29379;
  wire _59795 = _9971 ^ _29387;
  wire _59796 = _59794 ^ _59795;
  wire _59797 = _59793 ^ _59796;
  wire _59798 = _10531 ^ _19268;
  wire _59799 = _32425 ^ _34906;
  wire _59800 = _59798 ^ _59799;
  wire _59801 = uncoded_block[1004] ^ uncoded_block[1010];
  wire _59802 = _2111 ^ _59801;
  wire _59803 = _48631 ^ _59802;
  wire _59804 = _59800 ^ _59803;
  wire _59805 = _59797 ^ _59804;
  wire _59806 = _59790 ^ _59805;
  wire _59807 = _59774 ^ _59806;
  wire _59808 = _59738 ^ _59807;
  wire _59809 = _8296 ^ _2894;
  wire _59810 = uncoded_block[1022] ^ uncoded_block[1033];
  wire _59811 = _59810 ^ _6474;
  wire _59812 = _59809 ^ _59811;
  wire _59813 = _6478 ^ _1356;
  wire _59814 = _8311 ^ _522;
  wire _59815 = _59813 ^ _59814;
  wire _59816 = _59812 ^ _59815;
  wire _59817 = uncoded_block[1065] ^ uncoded_block[1072];
  wire _59818 = _59817 ^ _29859;
  wire _59819 = _5163 ^ _17369;
  wire _59820 = _59818 ^ _59819;
  wire _59821 = _15405 ^ _19795;
  wire _59822 = uncoded_block[1125] ^ uncoded_block[1133];
  wire _59823 = _59822 ^ _564;
  wire _59824 = _59821 ^ _59823;
  wire _59825 = _59820 ^ _59824;
  wire _59826 = _59816 ^ _59825;
  wire _59827 = _2188 ^ _49385;
  wire _59828 = _55071 ^ _59827;
  wire _59829 = uncoded_block[1182] ^ uncoded_block[1196];
  wire _59830 = _5872 ^ _59829;
  wire _59831 = _8951 ^ _6529;
  wire _59832 = _59830 ^ _59831;
  wire _59833 = _59828 ^ _59832;
  wire _59834 = _23544 ^ _54471;
  wire _59835 = uncoded_block[1225] ^ uncoded_block[1235];
  wire _59836 = _59835 ^ _2989;
  wire _59837 = _59834 ^ _59836;
  wire _59838 = uncoded_block[1238] ^ uncoded_block[1244];
  wire _59839 = _59838 ^ _2232;
  wire _59840 = uncoded_block[1249] ^ uncoded_block[1260];
  wire _59841 = _59840 ^ _34563;
  wire _59842 = _59839 ^ _59841;
  wire _59843 = _59837 ^ _59842;
  wire _59844 = _59833 ^ _59843;
  wire _59845 = _59826 ^ _59844;
  wire _59846 = uncoded_block[1268] ^ uncoded_block[1274];
  wire _59847 = _59846 ^ _1463;
  wire _59848 = uncoded_block[1278] ^ uncoded_block[1296];
  wire _59849 = _59848 ^ _20812;
  wire _59850 = _59847 ^ _59849;
  wire _59851 = _3807 ^ _2261;
  wire _59852 = uncoded_block[1317] ^ uncoded_block[1323];
  wire _59853 = _59852 ^ _16435;
  wire _59854 = _59851 ^ _59853;
  wire _59855 = _59850 ^ _59854;
  wire _59856 = _9564 ^ _13401;
  wire _59857 = _5260 ^ _59856;
  wire _59858 = _50644 ^ _7821;
  wire _59859 = uncoded_block[1366] ^ uncoded_block[1381];
  wire _59860 = uncoded_block[1382] ^ uncoded_block[1390];
  wire _59861 = _59859 ^ _59860;
  wire _59862 = _59858 ^ _59861;
  wire _59863 = _59857 ^ _59862;
  wire _59864 = _59855 ^ _59863;
  wire _59865 = _21774 ^ _2296;
  wire _59866 = _59865 ^ _7836;
  wire _59867 = uncoded_block[1416] ^ uncoded_block[1424];
  wire _59868 = _1523 ^ _59867;
  wire _59869 = _7844 ^ _47970;
  wire _59870 = _59868 ^ _59869;
  wire _59871 = _59866 ^ _59870;
  wire _59872 = uncoded_block[1436] ^ uncoded_block[1447];
  wire _59873 = uncoded_block[1450] ^ uncoded_block[1454];
  wire _59874 = _59872 ^ _59873;
  wire _59875 = _14985 ^ _20855;
  wire _59876 = _59874 ^ _59875;
  wire _59877 = _14989 ^ _5990;
  wire _59878 = _6631 ^ _44357;
  wire _59879 = _59877 ^ _59878;
  wire _59880 = _59876 ^ _59879;
  wire _59881 = _59871 ^ _59880;
  wire _59882 = _59864 ^ _59881;
  wire _59883 = _59845 ^ _59882;
  wire _59884 = _18931 ^ _7875;
  wire _59885 = _9055 ^ _4620;
  wire _59886 = _59884 ^ _59885;
  wire _59887 = uncoded_block[1523] ^ uncoded_block[1529];
  wire _59888 = _59887 ^ _11820;
  wire _59889 = uncoded_block[1536] ^ uncoded_block[1544];
  wire _59890 = _59889 ^ _18492;
  wire _59891 = _59888 ^ _59890;
  wire _59892 = _59886 ^ _59891;
  wire _59893 = _16501 ^ _4644;
  wire _59894 = _10163 ^ _784;
  wire _59895 = _59893 ^ _59894;
  wire _59896 = uncoded_block[1593] ^ uncoded_block[1599];
  wire _59897 = _5371 ^ _59896;
  wire _59898 = _9088 ^ _42166;
  wire _59899 = _59897 ^ _59898;
  wire _59900 = _59895 ^ _59899;
  wire _59901 = _59892 ^ _59900;
  wire _59902 = _47634 ^ _10185;
  wire _59903 = uncoded_block[1627] ^ uncoded_block[1635];
  wire _59904 = _59903 ^ _51456;
  wire _59905 = _59902 ^ _59904;
  wire _59906 = _815 ^ _9661;
  wire _59907 = uncoded_block[1660] ^ uncoded_block[1667];
  wire _59908 = _9106 ^ _59907;
  wire _59909 = _59906 ^ _59908;
  wire _59910 = _59905 ^ _59909;
  wire _59911 = uncoded_block[1675] ^ uncoded_block[1698];
  wire _59912 = _2422 ^ _59911;
  wire _59913 = _8536 ^ _4703;
  wire _59914 = _59912 ^ _59913;
  wire _59915 = _59914 ^ uncoded_block[1722];
  wire _59916 = _59910 ^ _59915;
  wire _59917 = _59901 ^ _59916;
  wire _59918 = _59883 ^ _59917;
  wire _59919 = _59808 ^ _59918;
  wire _59920 = uncoded_block[11] ^ uncoded_block[18];
  wire _59921 = _19959 ^ _59920;
  wire _59922 = _15076 ^ _11343;
  wire _59923 = _59921 ^ _59922;
  wire _59924 = uncoded_block[27] ^ uncoded_block[60];
  wire _59925 = uncoded_block[63] ^ uncoded_block[68];
  wire _59926 = _59924 ^ _59925;
  wire _59927 = _11904 ^ _11363;
  wire _59928 = _59926 ^ _59927;
  wire _59929 = _59923 ^ _59928;
  wire _59930 = uncoded_block[105] ^ uncoded_block[115];
  wire _59931 = _59930 ^ _33056;
  wire _59932 = _10821 ^ _2504;
  wire _59933 = _59931 ^ _59932;
  wire _59934 = _3265 ^ _3272;
  wire _59935 = uncoded_block[164] ^ uncoded_block[177];
  wire _59936 = _59935 ^ _9195;
  wire _59937 = _59934 ^ _59936;
  wire _59938 = _59933 ^ _59937;
  wire _59939 = _59929 ^ _59938;
  wire _59940 = uncoded_block[189] ^ uncoded_block[199];
  wire _59941 = _59940 ^ _98;
  wire _59942 = uncoded_block[219] ^ uncoded_block[229];
  wire _59943 = _959 ^ _59942;
  wire _59944 = _59941 ^ _59943;
  wire _59945 = uncoded_block[238] ^ uncoded_block[251];
  wire _59946 = _59945 ^ _14639;
  wire _59947 = uncoded_block[277] ^ uncoded_block[287];
  wire _59948 = uncoded_block[288] ^ uncoded_block[296];
  wire _59949 = _59947 ^ _59948;
  wire _59950 = _59946 ^ _59949;
  wire _59951 = _59944 ^ _59950;
  wire _59952 = _29656 ^ _22866;
  wire _59953 = _145 ^ _9780;
  wire _59954 = _59952 ^ _59953;
  wire _59955 = uncoded_block[328] ^ uncoded_block[337];
  wire _59956 = _59955 ^ _2593;
  wire _59957 = _16158 ^ _4844;
  wire _59958 = _59956 ^ _59957;
  wire _59959 = _59954 ^ _59958;
  wire _59960 = _59951 ^ _59959;
  wire _59961 = _59939 ^ _59960;
  wire _59962 = uncoded_block[351] ^ uncoded_block[367];
  wire _59963 = uncoded_block[368] ^ uncoded_block[382];
  wire _59964 = _59962 ^ _59963;
  wire _59965 = uncoded_block[385] ^ uncoded_block[399];
  wire _59966 = _59965 ^ _10344;
  wire _59967 = _59964 ^ _59966;
  wire _59968 = uncoded_block[418] ^ uncoded_block[425];
  wire _59969 = _59968 ^ _21974;
  wire _59970 = _31453 ^ _59969;
  wire _59971 = _59967 ^ _59970;
  wire _59972 = _26491 ^ _32709;
  wire _59973 = _30155 ^ _6906;
  wire _59974 = _59972 ^ _59973;
  wire _59975 = uncoded_block[508] ^ uncoded_block[523];
  wire _59976 = _59975 ^ _15230;
  wire _59977 = _25168 ^ _59976;
  wire _59978 = _59974 ^ _59977;
  wire _59979 = _59971 ^ _59978;
  wire _59980 = _52785 ^ _1909;
  wire _59981 = _1122 ^ _31907;
  wire _59982 = _59980 ^ _59981;
  wire _59983 = uncoded_block[572] ^ uncoded_block[579];
  wire _59984 = _59983 ^ _3475;
  wire _59985 = _59984 ^ _32743;
  wire _59986 = _59982 ^ _59985;
  wire _59987 = uncoded_block[593] ^ uncoded_block[600];
  wire _59988 = uncoded_block[610] ^ uncoded_block[617];
  wire _59989 = _59987 ^ _59988;
  wire _59990 = uncoded_block[625] ^ uncoded_block[633];
  wire _59991 = _59990 ^ _55587;
  wire _59992 = _59989 ^ _59991;
  wire _59993 = _31929 ^ _1164;
  wire _59994 = _13188 ^ _3521;
  wire _59995 = _59993 ^ _59994;
  wire _59996 = _59992 ^ _59995;
  wire _59997 = _59986 ^ _59996;
  wire _59998 = _59979 ^ _59997;
  wire _59999 = _59961 ^ _59998;
  wire _60000 = uncoded_block[680] ^ uncoded_block[689];
  wire _60001 = _60000 ^ _2754;
  wire _60002 = uncoded_block[698] ^ uncoded_block[708];
  wire _60003 = _4987 ^ _60002;
  wire _60004 = _60001 ^ _60003;
  wire _60005 = uncoded_block[710] ^ uncoded_block[719];
  wire _60006 = _60005 ^ _8200;
  wire _60007 = uncoded_block[746] ^ uncoded_block[751];
  wire _60008 = _41193 ^ _60007;
  wire _60009 = _60006 ^ _60008;
  wire _60010 = _60004 ^ _60009;
  wire _60011 = uncoded_block[790] ^ uncoded_block[796];
  wire _60012 = _364 ^ _60011;
  wire _60013 = _16791 ^ _10485;
  wire _60014 = _60012 ^ _60013;
  wire _60015 = uncoded_block[839] ^ uncoded_block[843];
  wire _60016 = _2808 ^ _60015;
  wire _60017 = _60016 ^ _37309;
  wire _60018 = _60014 ^ _60017;
  wire _60019 = _60010 ^ _60018;
  wire _60020 = uncoded_block[858] ^ uncoded_block[873];
  wire _60021 = uncoded_block[883] ^ uncoded_block[893];
  wire _60022 = _60020 ^ _60021;
  wire _60023 = uncoded_block[898] ^ uncoded_block[907];
  wire _60024 = uncoded_block[909] ^ uncoded_block[917];
  wire _60025 = _60023 ^ _60024;
  wire _60026 = _60022 ^ _60025;
  wire _60027 = _15350 ^ _12169;
  wire _60028 = uncoded_block[939] ^ uncoded_block[950];
  wire _60029 = _60028 ^ _5105;
  wire _60030 = _60027 ^ _60029;
  wire _60031 = _60026 ^ _60030;
  wire _60032 = _12180 ^ _11091;
  wire _60033 = uncoded_block[980] ^ uncoded_block[985];
  wire _60034 = uncoded_block[986] ^ uncoded_block[994];
  wire _60035 = _60033 ^ _60034;
  wire _60036 = _60032 ^ _60035;
  wire _60037 = uncoded_block[998] ^ uncoded_block[1011];
  wire _60038 = _60037 ^ _8868;
  wire _60039 = _35708 ^ _2898;
  wire _60040 = _60038 ^ _60039;
  wire _60041 = _60036 ^ _60040;
  wire _60042 = _60031 ^ _60041;
  wire _60043 = _60019 ^ _60042;
  wire _60044 = uncoded_block[1042] ^ uncoded_block[1062];
  wire _60045 = _60044 ^ _15395;
  wire _60046 = _26661 ^ _9478;
  wire _60047 = _60045 ^ _60046;
  wire _60048 = uncoded_block[1113] ^ uncoded_block[1121];
  wire _60049 = _60048 ^ _2942;
  wire _60050 = _40138 ^ _60049;
  wire _60051 = _60047 ^ _60050;
  wire _60052 = _12791 ^ _15896;
  wire _60053 = uncoded_block[1147] ^ uncoded_block[1165];
  wire _60054 = _45022 ^ _60053;
  wire _60055 = _60052 ^ _60054;
  wire _60056 = uncoded_block[1184] ^ uncoded_block[1192];
  wire _60057 = _60056 ^ _8951;
  wire _60058 = _14902 ^ _60057;
  wire _60059 = _60055 ^ _60058;
  wire _60060 = _60051 ^ _60059;
  wire _60061 = uncoded_block[1209] ^ uncoded_block[1226];
  wire _60062 = _11722 ^ _60061;
  wire _60063 = uncoded_block[1227] ^ uncoded_block[1245];
  wire _60064 = _60063 ^ _2998;
  wire _60065 = _60062 ^ _60064;
  wire _60066 = _4514 ^ _9532;
  wire _60067 = uncoded_block[1284] ^ uncoded_block[1294];
  wire _60068 = _60067 ^ _7799;
  wire _60069 = _60066 ^ _60068;
  wire _60070 = _60065 ^ _60069;
  wire _60071 = uncoded_block[1316] ^ uncoded_block[1321];
  wire _60072 = _60071 ^ _34996;
  wire _60073 = _657 ^ _23576;
  wire _60074 = _60072 ^ _60073;
  wire _60075 = _3823 ^ _23148;
  wire _60076 = uncoded_block[1366] ^ uncoded_block[1376];
  wire _60077 = uncoded_block[1377] ^ uncoded_block[1385];
  wire _60078 = _60076 ^ _60077;
  wire _60079 = _60075 ^ _60078;
  wire _60080 = _60074 ^ _60079;
  wire _60081 = _60070 ^ _60080;
  wire _60082 = _60060 ^ _60081;
  wire _60083 = _60043 ^ _60082;
  wire _60084 = _59999 ^ _60083;
  wire _60085 = uncoded_block[1387] ^ uncoded_block[1394];
  wire _60086 = _60085 ^ _3846;
  wire _60087 = uncoded_block[1408] ^ uncoded_block[1433];
  wire _60088 = _2300 ^ _60087;
  wire _60089 = _60086 ^ _60088;
  wire _60090 = _24521 ^ _716;
  wire _60091 = uncoded_block[1458] ^ uncoded_block[1471];
  wire _60092 = _20852 ^ _60091;
  wire _60093 = _60090 ^ _60092;
  wire _60094 = _60089 ^ _60093;
  wire _60095 = uncoded_block[1487] ^ uncoded_block[1494];
  wire _60096 = _5316 ^ _60095;
  wire _60097 = uncoded_block[1501] ^ uncoded_block[1523];
  wire _60098 = uncoded_block[1527] ^ uncoded_block[1534];
  wire _60099 = _60097 ^ _60098;
  wire _60100 = _60096 ^ _60099;
  wire _60101 = _10157 ^ _29986;
  wire _60102 = _782 ^ _1609;
  wire _60103 = _60101 ^ _60102;
  wire _60104 = _60100 ^ _60103;
  wire _60105 = _60094 ^ _60104;
  wire _60106 = uncoded_block[1594] ^ uncoded_block[1604];
  wire _60107 = uncoded_block[1605] ^ uncoded_block[1620];
  wire _60108 = _60106 ^ _60107;
  wire _60109 = _60108 ^ _39462;
  wire _60110 = uncoded_block[1639] ^ uncoded_block[1643];
  wire _60111 = uncoded_block[1644] ^ uncoded_block[1657];
  wire _60112 = _60110 ^ _60111;
  wire _60113 = _29569 ^ _17032;
  wire _60114 = _60112 ^ _60113;
  wire _60115 = _60109 ^ _60114;
  wire _60116 = uncoded_block[1672] ^ uncoded_block[1686];
  wire _60117 = uncoded_block[1695] ^ uncoded_block[1704];
  wire _60118 = _60116 ^ _60117;
  wire _60119 = _15063 ^ _54215;
  wire _60120 = _60118 ^ _60119;
  wire _60121 = _14552 ^ uncoded_block[1719];
  wire _60122 = _60120 ^ _60121;
  wire _60123 = _60115 ^ _60122;
  wire _60124 = _60105 ^ _60123;
  wire _60125 = _60084 ^ _60124;
  wire _60126 = uncoded_block[8] ^ uncoded_block[15];
  wire _60127 = _18539 ^ _60126;
  wire _60128 = _60127 ^ _55824;
  wire _60129 = _4001 ^ _874;
  wire _60130 = _3225 ^ _3227;
  wire _60131 = _60129 ^ _60130;
  wire _60132 = _60128 ^ _60131;
  wire _60133 = _2466 ^ _7965;
  wire _60134 = _12425 ^ _22795;
  wire _60135 = _60133 ^ _60134;
  wire _60136 = _4726 ^ _1703;
  wire _60137 = _2472 ^ _9705;
  wire _60138 = _60136 ^ _60137;
  wire _60139 = _60135 ^ _60138;
  wire _60140 = _60132 ^ _60139;
  wire _60141 = _50732 ^ _50011;
  wire _60142 = _14586 ^ _7981;
  wire _60143 = _4736 ^ _60142;
  wire _60144 = _60141 ^ _60143;
  wire _60145 = _20952 ^ _47;
  wire _60146 = _4745 ^ _4031;
  wire _60147 = _60145 ^ _60146;
  wire _60148 = _19028 ^ _19523;
  wire _60149 = _60147 ^ _60148;
  wire _60150 = _60144 ^ _60149;
  wire _60151 = _60140 ^ _60150;
  wire _60152 = _2499 ^ _43281;
  wire _60153 = _8581 ^ _4760;
  wire _60154 = _22358 ^ _60153;
  wire _60155 = _60152 ^ _60154;
  wire _60156 = _7999 ^ _55477;
  wire _60157 = _9186 ^ _23281;
  wire _60158 = _60156 ^ _60157;
  wire _60159 = _16604 ^ _5473;
  wire _60160 = _25532 ^ _60159;
  wire _60161 = _60158 ^ _60160;
  wire _60162 = _60155 ^ _60161;
  wire _60163 = _15123 ^ _20979;
  wire _60164 = _18110 ^ _1759;
  wire _60165 = _60163 ^ _60164;
  wire _60166 = _18111 ^ _2531;
  wire _60167 = _18583 ^ _10849;
  wire _60168 = _60166 ^ _60167;
  wire _60169 = _60165 ^ _60168;
  wire _60170 = uncoded_block[211] ^ uncoded_block[214];
  wire _60171 = _58384 ^ _60170;
  wire _60172 = _39141 ^ _60171;
  wire _60173 = _5492 ^ _2545;
  wire _60174 = _21461 ^ _60173;
  wire _60175 = _60172 ^ _60174;
  wire _60176 = _60169 ^ _60175;
  wire _60177 = _60162 ^ _60176;
  wire _60178 = _60151 ^ _60177;
  wire _60179 = _4082 ^ _7424;
  wire _60180 = _7425 ^ _6179;
  wire _60181 = _16626 ^ _4800;
  wire _60182 = _60180 ^ _60181;
  wire _60183 = _60179 ^ _60182;
  wire _60184 = _20519 ^ _6189;
  wire _60185 = _21472 ^ _14124;
  wire _60186 = _6833 ^ _7445;
  wire _60187 = _60185 ^ _60186;
  wire _60188 = _60184 ^ _60187;
  wire _60189 = _60183 ^ _60188;
  wire _60190 = _3327 ^ _38762;
  wire _60191 = _11425 ^ _60190;
  wire _60192 = _13615 ^ _4824;
  wire _60193 = _12515 ^ _22866;
  wire _60194 = _60192 ^ _60193;
  wire _60195 = _60191 ^ _60194;
  wire _60196 = uncoded_block[328] ^ uncoded_block[333];
  wire _60197 = _21947 ^ _60196;
  wire _60198 = _21943 ^ _60197;
  wire _60199 = _15173 ^ _9242;
  wire _60200 = _60199 ^ _3356;
  wire _60201 = _60198 ^ _60200;
  wire _60202 = _60195 ^ _60201;
  wire _60203 = _60189 ^ _60202;
  wire _60204 = _3359 ^ _42277;
  wire _60205 = _20554 ^ _35170;
  wire _60206 = _60204 ^ _60205;
  wire _60207 = uncoded_block[371] ^ uncoded_block[374];
  wire _60208 = _60207 ^ _8079;
  wire _60209 = _1836 ^ _60208;
  wire _60210 = _60206 ^ _60209;
  wire _60211 = _46607 ^ _10907;
  wire _60212 = _47736 ^ _60211;
  wire _60213 = _15696 ^ _183;
  wire _60214 = _184 ^ _11473;
  wire _60215 = _60213 ^ _60214;
  wire _60216 = _60212 ^ _60215;
  wire _60217 = _60210 ^ _60216;
  wire _60218 = _8092 ^ _6249;
  wire _60219 = _60218 ^ _4165;
  wire _60220 = _2633 ^ _1062;
  wire _60221 = _34771 ^ _13117;
  wire _60222 = _60220 ^ _60221;
  wire _60223 = _60219 ^ _60222;
  wire _60224 = _34379 ^ _54677;
  wire _60225 = _5590 ^ _1085;
  wire _60226 = _36805 ^ _60225;
  wire _60227 = _60224 ^ _60226;
  wire _60228 = _60223 ^ _60227;
  wire _60229 = _60217 ^ _60228;
  wire _60230 = _60203 ^ _60229;
  wire _60231 = _60178 ^ _60230;
  wire _60232 = _12028 ^ _4897;
  wire _60233 = _5600 ^ _14183;
  wire _60234 = _60232 ^ _60233;
  wire _60235 = _33992 ^ _39994;
  wire _60236 = _60234 ^ _60235;
  wire _60237 = _43360 ^ _46252;
  wire _60238 = _1108 ^ _9301;
  wire _60239 = _6290 ^ _16215;
  wire _60240 = _60238 ^ _60239;
  wire _60241 = _60237 ^ _60240;
  wire _60242 = _60236 ^ _60241;
  wire _60243 = _3451 ^ _25173;
  wire _60244 = _60243 ^ _26520;
  wire _60245 = _25182 ^ _9319;
  wire _60246 = _9320 ^ _18682;
  wire _60247 = _60245 ^ _60246;
  wire _60248 = _60244 ^ _60247;
  wire _60249 = _1931 ^ _4229;
  wire _60250 = _4225 ^ _60249;
  wire _60251 = _2696 ^ _4233;
  wire _60252 = _2700 ^ _17721;
  wire _60253 = _60251 ^ _60252;
  wire _60254 = _60250 ^ _60253;
  wire _60255 = _60248 ^ _60254;
  wire _60256 = _60242 ^ _60255;
  wire _60257 = _5648 ^ _33608;
  wire _60258 = _6960 ^ _2719;
  wire _60259 = _60258 ^ _51240;
  wire _60260 = _60257 ^ _60259;
  wire _60261 = uncoded_block[643] ^ uncoded_block[647];
  wire _60262 = _29741 ^ _60261;
  wire _60263 = _25206 ^ _4975;
  wire _60264 = _60262 ^ _60263;
  wire _60265 = _40030 ^ _13726;
  wire _60266 = _311 ^ _15775;
  wire _60267 = _60265 ^ _60266;
  wire _60268 = _60264 ^ _60267;
  wire _60269 = _60260 ^ _60268;
  wire _60270 = uncoded_block[679] ^ uncoded_block[684];
  wire _60271 = _13731 ^ _60270;
  wire _60272 = _60271 ^ _29755;
  wire _60273 = uncoded_block[705] ^ uncoded_block[710];
  wire _60274 = _45691 ^ _60273;
  wire _60275 = _330 ^ _60274;
  wire _60276 = _60272 ^ _60275;
  wire _60277 = _49778 ^ _13745;
  wire _60278 = uncoded_block[732] ^ uncoded_block[740];
  wire _60279 = _4283 ^ _60278;
  wire _60280 = _7006 ^ _5702;
  wire _60281 = _60279 ^ _60280;
  wire _60282 = _60277 ^ _60281;
  wire _60283 = _60276 ^ _60282;
  wire _60284 = _60269 ^ _60283;
  wire _60285 = _60256 ^ _60284;
  wire _60286 = _5013 ^ _2777;
  wire _60287 = _60286 ^ _9913;
  wire _60288 = _26579 ^ _5709;
  wire _60289 = _60288 ^ _18745;
  wire _60290 = _60287 ^ _60289;
  wire _60291 = _3562 ^ _34862;
  wire _60292 = _60291 ^ _25237;
  wire _60293 = _15806 ^ _36054;
  wire _60294 = _60292 ^ _60293;
  wire _60295 = _60290 ^ _60294;
  wire _60296 = _48591 ^ _31114;
  wire _60297 = _4325 ^ _45332;
  wire _60298 = _55991 ^ _1249;
  wire _60299 = _60297 ^ _60298;
  wire _60300 = _60296 ^ _60299;
  wire _60301 = _47836 ^ _14812;
  wire _60302 = _19233 ^ _60301;
  wire _60303 = _2044 ^ _29368;
  wire _60304 = _60303 ^ _22086;
  wire _60305 = _60302 ^ _60304;
  wire _60306 = _60300 ^ _60305;
  wire _60307 = _60295 ^ _60306;
  wire _60308 = _6416 ^ _41628;
  wire _60309 = _14303 ^ _60308;
  wire _60310 = _55042 ^ _7660;
  wire _60311 = _11060 ^ _14829;
  wire _60312 = _60310 ^ _60311;
  wire _60313 = _60309 ^ _60312;
  wire _60314 = _46035 ^ _49819;
  wire _60315 = _7665 ^ _42399;
  wire _60316 = _60314 ^ _60315;
  wire _60317 = _5772 ^ _448;
  wire _60318 = _60317 ^ _454;
  wire _60319 = _60316 ^ _60318;
  wire _60320 = _60313 ^ _60319;
  wire _60321 = _2865 ^ _13266;
  wire _60322 = _60321 ^ _42018;
  wire _60323 = _11643 ^ _12180;
  wire _60324 = _11649 ^ _5790;
  wire _60325 = _60323 ^ _60324;
  wire _60326 = _60322 ^ _60325;
  wire _60327 = _55311 ^ _34908;
  wire _60328 = _2883 ^ _22584;
  wire _60329 = _60328 ^ _58555;
  wire _60330 = _60327 ^ _60329;
  wire _60331 = _60326 ^ _60330;
  wire _60332 = _60320 ^ _60331;
  wire _60333 = _60307 ^ _60332;
  wire _60334 = _60285 ^ _60333;
  wire _60335 = _60231 ^ _60334;
  wire _60336 = _13283 ^ _9996;
  wire _60337 = _60336 ^ _6464;
  wire _60338 = _53228 ^ _3675;
  wire _60339 = _60338 ^ _48639;
  wire _60340 = _60337 ^ _60339;
  wire _60341 = _48641 ^ _59337;
  wire _60342 = _5147 ^ _8311;
  wire _60343 = _60341 ^ _60342;
  wire _60344 = _6483 ^ _42044;
  wire _60345 = _60344 ^ _42429;
  wire _60346 = _60343 ^ _60345;
  wire _60347 = _60340 ^ _60346;
  wire _60348 = _9478 ^ _20251;
  wire _60349 = _20753 ^ _13311;
  wire _60350 = _60348 ^ _60349;
  wire _60351 = _10021 ^ _29014;
  wire _60352 = uncoded_block[1100] ^ uncoded_block[1104];
  wire _60353 = _1380 ^ _60352;
  wire _60354 = _60351 ^ _60353;
  wire _60355 = _60350 ^ _60354;
  wire _60356 = _8917 ^ _3713;
  wire _60357 = _34532 ^ _60356;
  wire _60358 = _11147 ^ _2944;
  wire _60359 = _4459 ^ _18371;
  wire _60360 = _60358 ^ _60359;
  wire _60361 = _60357 ^ _60360;
  wire _60362 = _60355 ^ _60361;
  wire _60363 = _60347 ^ _60362;
  wire _60364 = _13866 ^ _14380;
  wire _60365 = uncoded_block[1140] ^ uncoded_block[1144];
  wire _60366 = _10593 ^ _60365;
  wire _60367 = _60364 ^ _60366;
  wire _60368 = _38557 ^ _27105;
  wire _60369 = _29026 ^ _60368;
  wire _60370 = _60367 ^ _60369;
  wire _60371 = _3736 ^ _2967;
  wire _60372 = _34961 ^ _35354;
  wire _60373 = _60371 ^ _60372;
  wire _60374 = _596 ^ _1421;
  wire _60375 = _19340 ^ _60374;
  wire _60376 = _60373 ^ _60375;
  wire _60377 = _60370 ^ _60376;
  wire _60378 = _44674 ^ _18395;
  wire _60379 = _17901 ^ _60378;
  wire _60380 = _4502 ^ _54853;
  wire _60381 = _23106 ^ _60380;
  wire _60382 = _60379 ^ _60381;
  wire _60383 = _38977 ^ _27560;
  wire _60384 = uncoded_block[1246] ^ uncoded_block[1252];
  wire _60385 = _60384 ^ _6546;
  wire _60386 = _5234 ^ _9532;
  wire _60387 = _60385 ^ _60386;
  wire _60388 = _60383 ^ _60387;
  wire _60389 = _60382 ^ _60388;
  wire _60390 = _60377 ^ _60389;
  wire _60391 = _60363 ^ _60390;
  wire _60392 = _1464 ^ _7794;
  wire _60393 = _7186 ^ _4530;
  wire _60394 = _60392 ^ _60393;
  wire _60395 = _13915 ^ _1479;
  wire _60396 = _60395 ^ _22667;
  wire _60397 = _58620 ^ _1489;
  wire _60398 = _8413 ^ _13399;
  wire _60399 = _60397 ^ _60398;
  wire _60400 = _60396 ^ _60399;
  wire _60401 = _60394 ^ _60400;
  wire _60402 = _1497 ^ _7815;
  wire _60403 = _18434 ^ _16942;
  wire _60404 = _60402 ^ _60403;
  wire _60405 = _5940 ^ _676;
  wire _60406 = _3828 ^ _7823;
  wire _60407 = _60405 ^ _60406;
  wire _60408 = _60404 ^ _60407;
  wire _60409 = _5284 ^ _7219;
  wire _60410 = _58634 ^ _18444;
  wire _60411 = _60409 ^ _60410;
  wire _60412 = _47205 ^ _6600;
  wire _60413 = _16954 ^ _5957;
  wire _60414 = _60412 ^ _60413;
  wire _60415 = _60411 ^ _60414;
  wire _60416 = _60408 ^ _60415;
  wire _60417 = _60401 ^ _60416;
  wire _60418 = _9022 ^ _32948;
  wire _60419 = _2313 ^ _9595;
  wire _60420 = _60418 ^ _60419;
  wire _60421 = _36629 ^ _60420;
  wire _60422 = _5304 ^ _716;
  wire _60423 = _60422 ^ _11248;
  wire _60424 = _11249 ^ _23614;
  wire _60425 = _4603 ^ _2344;
  wire _60426 = _60424 ^ _60425;
  wire _60427 = _60423 ^ _60426;
  wire _60428 = _60421 ^ _60427;
  wire _60429 = _19887 ^ _5990;
  wire _60430 = _12896 ^ _2352;
  wire _60431 = _60429 ^ _60430;
  wire _60432 = _747 ^ _11813;
  wire _60433 = _60432 ^ _23628;
  wire _60434 = _60431 ^ _60433;
  wire _60435 = _36655 ^ _44364;
  wire _60436 = uncoded_block[1535] ^ uncoded_block[1544];
  wire _60437 = _3905 ^ _60436;
  wire _60438 = _60435 ^ _60437;
  wire _60439 = _767 ^ _769;
  wire _60440 = _22731 ^ _1597;
  wire _60441 = _60439 ^ _60440;
  wire _60442 = _60438 ^ _60441;
  wire _60443 = _60434 ^ _60442;
  wire _60444 = _60428 ^ _60443;
  wire _60445 = _60417 ^ _60444;
  wire _60446 = _60391 ^ _60445;
  wire _60447 = _56614 ^ _4648;
  wire _60448 = _32158 ^ _60447;
  wire _60449 = _6663 ^ _40243;
  wire _60450 = _60449 ^ _17014;
  wire _60451 = _60448 ^ _60450;
  wire _60452 = _27968 ^ _2396;
  wire _60453 = _14520 ^ _9647;
  wire _60454 = _60452 ^ _60453;
  wire _60455 = _27649 ^ _5388;
  wire _60456 = _9659 ^ _7309;
  wire _60457 = _60455 ^ _60456;
  wire _60458 = _60454 ^ _60457;
  wire _60459 = _60451 ^ _60458;
  wire _60460 = _32178 ^ _820;
  wire _60461 = _33856 ^ _60460;
  wire _60462 = _19466 ^ _25476;
  wire _60463 = _27979 ^ _60462;
  wire _60464 = _60461 ^ _60463;
  wire _60465 = _3186 ^ _17040;
  wire _60466 = _17037 ^ _60465;
  wire _60467 = _59238 ^ _840;
  wire _60468 = _60467 ^ _42840;
  wire _60469 = _60466 ^ _60468;
  wire _60470 = _60464 ^ _60469;
  wire _60471 = _60459 ^ _60470;
  wire _60472 = uncoded_block[1704] ^ uncoded_block[1709];
  wire _60473 = _60472 ^ _55813;
  wire _60474 = _60473 ^ _39873;
  wire _60475 = _60471 ^ _60474;
  wire _60476 = _60446 ^ _60475;
  wire _60477 = _60335 ^ _60476;
  wire _60478 = uncoded_block[10] ^ uncoded_block[19];
  wire _60479 = _41026 ^ _60478;
  wire _60480 = uncoded_block[38] ^ uncoded_block[46];
  wire _60481 = uncoded_block[64] ^ uncoded_block[76];
  wire _60482 = _60480 ^ _60481;
  wire _60483 = _60479 ^ _60482;
  wire _60484 = uncoded_block[99] ^ uncoded_block[110];
  wire _60485 = _41044 ^ _60484;
  wire _60486 = uncoded_block[116] ^ uncoded_block[125];
  wire _60487 = uncoded_block[126] ^ uncoded_block[133];
  wire _60488 = _60486 ^ _60487;
  wire _60489 = _60485 ^ _60488;
  wire _60490 = _60483 ^ _60489;
  wire _60491 = uncoded_block[176] ^ uncoded_block[184];
  wire _60492 = _22819 ^ _60491;
  wire _60493 = uncoded_block[198] ^ uncoded_block[214];
  wire _60494 = uncoded_block[228] ^ uncoded_block[251];
  wire _60495 = _60493 ^ _60494;
  wire _60496 = _60492 ^ _60495;
  wire _60497 = _17628 ^ _7438;
  wire _60498 = _33522 ^ _30106;
  wire _60499 = _60497 ^ _60498;
  wire _60500 = _60496 ^ _60499;
  wire _60501 = _60490 ^ _60500;
  wire _60502 = uncoded_block[311] ^ uncoded_block[322];
  wire _60503 = uncoded_block[334] ^ uncoded_block[350];
  wire _60504 = _60502 ^ _60503;
  wire _60505 = uncoded_block[356] ^ uncoded_block[368];
  wire _60506 = _60505 ^ _35563;
  wire _60507 = _60504 ^ _60506;
  wire _60508 = uncoded_block[404] ^ uncoded_block[420];
  wire _60509 = _17668 ^ _60508;
  wire _60510 = uncoded_block[422] ^ uncoded_block[429];
  wire _60511 = uncoded_block[450] ^ uncoded_block[469];
  wire _60512 = _60510 ^ _60511;
  wire _60513 = _60509 ^ _60512;
  wire _60514 = _60507 ^ _60513;
  wire _60515 = uncoded_block[476] ^ uncoded_block[496];
  wire _60516 = _60515 ^ _21992;
  wire _60517 = uncoded_block[522] ^ uncoded_block[540];
  wire _60518 = _60517 ^ _1126;
  wire _60519 = _60516 ^ _60518;
  wire _60520 = uncoded_block[584] ^ uncoded_block[601];
  wire _60521 = _60520 ^ _15758;
  wire _60522 = uncoded_block[621] ^ uncoded_block[635];
  wire _60523 = uncoded_block[654] ^ uncoded_block[664];
  wire _60524 = _60522 ^ _60523;
  wire _60525 = _60521 ^ _60524;
  wire _60526 = _60519 ^ _60525;
  wire _60527 = _60514 ^ _60526;
  wire _60528 = _60501 ^ _60527;
  wire _60529 = _14240 ^ _23412;
  wire _60530 = uncoded_block[686] ^ uncoded_block[726];
  wire _60531 = uncoded_block[729] ^ uncoded_block[746];
  wire _60532 = _60530 ^ _60531;
  wire _60533 = _60529 ^ _60532;
  wire _60534 = uncoded_block[750] ^ uncoded_block[762];
  wire _60535 = uncoded_block[768] ^ uncoded_block[784];
  wire _60536 = _60534 ^ _60535;
  wire _60537 = _55619 ^ _24804;
  wire _60538 = _60536 ^ _60537;
  wire _60539 = _60533 ^ _60538;
  wire _60540 = uncoded_block[817] ^ uncoded_block[834];
  wire _60541 = uncoded_block[835] ^ uncoded_block[860];
  wire _60542 = _60540 ^ _60541;
  wire _60543 = uncoded_block[878] ^ uncoded_block[893];
  wire _60544 = _17304 ^ _60543;
  wire _60545 = _60542 ^ _60544;
  wire _60546 = _5761 ^ _12165;
  wire _60547 = uncoded_block[925] ^ uncoded_block[947];
  wire _60548 = uncoded_block[949] ^ uncoded_block[968];
  wire _60549 = _60547 ^ _60548;
  wire _60550 = _60546 ^ _60549;
  wire _60551 = _60545 ^ _60550;
  wire _60552 = _60539 ^ _60551;
  wire _60553 = uncoded_block[984] ^ uncoded_block[989];
  wire _60554 = uncoded_block[993] ^ uncoded_block[1012];
  wire _60555 = _60553 ^ _60554;
  wire _60556 = uncoded_block[1035] ^ uncoded_block[1049];
  wire _60557 = _35710 ^ _60556;
  wire _60558 = _60555 ^ _60557;
  wire _60559 = uncoded_block[1052] ^ uncoded_block[1067];
  wire _60560 = _60559 ^ _22149;
  wire _60561 = uncoded_block[1107] ^ uncoded_block[1114];
  wire _60562 = _36955 ^ _60561;
  wire _60563 = _60560 ^ _60562;
  wire _60564 = _60558 ^ _60563;
  wire _60565 = uncoded_block[1127] ^ uncoded_block[1140];
  wire _60566 = _60565 ^ _4466;
  wire _60567 = uncoded_block[1158] ^ uncoded_block[1169];
  wire _60568 = uncoded_block[1175] ^ uncoded_block[1200];
  wire _60569 = _60567 ^ _60568;
  wire _60570 = _60566 ^ _60569;
  wire _60571 = uncoded_block[1218] ^ uncoded_block[1238];
  wire _60572 = _2207 ^ _60571;
  wire _60573 = uncoded_block[1252] ^ uncoded_block[1260];
  wire _60574 = _32903 ^ _60573;
  wire _60575 = _60572 ^ _60574;
  wire _60576 = _60570 ^ _60575;
  wire _60577 = _60564 ^ _60576;
  wire _60578 = _60552 ^ _60577;
  wire _60579 = _60528 ^ _60578;
  wire _60580 = uncoded_block[1270] ^ uncoded_block[1280];
  wire _60581 = uncoded_block[1283] ^ uncoded_block[1290];
  wire _60582 = _60580 ^ _60581;
  wire _60583 = uncoded_block[1301] ^ uncoded_block[1346];
  wire _60584 = _60583 ^ _54498;
  wire _60585 = _60582 ^ _60584;
  wire _60586 = uncoded_block[1389] ^ uncoded_block[1395];
  wire _60587 = _27160 ^ _60586;
  wire _60588 = uncoded_block[1406] ^ uncoded_block[1413];
  wire _60589 = uncoded_block[1416] ^ uncoded_block[1433];
  wire _60590 = _60588 ^ _60589;
  wire _60591 = _60587 ^ _60590;
  wire _60592 = _60585 ^ _60591;
  wire _60593 = uncoded_block[1455] ^ uncoded_block[1464];
  wire _60594 = _1541 ^ _60593;
  wire _60595 = uncoded_block[1526] ^ uncoded_block[1536];
  wire _60596 = uncoded_block[1539] ^ uncoded_block[1549];
  wire _60597 = _60595 ^ _60596;
  wire _60598 = _60594 ^ _60597;
  wire _60599 = uncoded_block[1564] ^ uncoded_block[1574];
  wire _60600 = _57554 ^ _60599;
  wire _60601 = uncoded_block[1592] ^ uncoded_block[1602];
  wire _60602 = _60601 ^ _22746;
  wire _60603 = _60600 ^ _60602;
  wire _60604 = _60598 ^ _60603;
  wire _60605 = _60592 ^ _60604;
  wire _60606 = _59392 ^ _12947;
  wire _60607 = uncoded_block[1636] ^ uncoded_block[1649];
  wire _60608 = _60607 ^ _24578;
  wire _60609 = _60606 ^ _60608;
  wire _60610 = uncoded_block[1657] ^ uncoded_block[1695];
  wire _60611 = _60610 ^ uncoded_block[1706];
  wire _60612 = _60609 ^ _60611;
  wire _60613 = _60605 ^ _60612;
  wire _60614 = _60579 ^ _60613;
  wire _60615 = uncoded_block[4] ^ uncoded_block[22];
  wire _60616 = uncoded_block[45] ^ uncoded_block[54];
  wire _60617 = _60615 ^ _60616;
  wire _60618 = _35 ^ _7377;
  wire _60619 = _60617 ^ _60618;
  wire _60620 = uncoded_block[141] ^ uncoded_block[161];
  wire _60621 = _22819 ^ _60620;
  wire _60622 = uncoded_block[169] ^ uncoded_block[185];
  wire _60623 = _60622 ^ _20500;
  wire _60624 = _60621 ^ _60623;
  wire _60625 = _60619 ^ _60624;
  wire _60626 = uncoded_block[204] ^ uncoded_block[209];
  wire _60627 = uncoded_block[226] ^ uncoded_block[239];
  wire _60628 = _60626 ^ _60627;
  wire _60629 = uncoded_block[264] ^ uncoded_block[300];
  wire _60630 = _5505 ^ _60629;
  wire _60631 = _60628 ^ _60630;
  wire _60632 = uncoded_block[302] ^ uncoded_block[315];
  wire _60633 = uncoded_block[321] ^ uncoded_block[328];
  wire _60634 = _60632 ^ _60633;
  wire _60635 = uncoded_block[350] ^ uncoded_block[372];
  wire _60636 = uncoded_block[374] ^ uncoded_block[387];
  wire _60637 = _60635 ^ _60636;
  wire _60638 = _60634 ^ _60637;
  wire _60639 = _60631 ^ _60638;
  wire _60640 = _60625 ^ _60639;
  wire _60641 = uncoded_block[388] ^ uncoded_block[406];
  wire _60642 = _60641 ^ _48499;
  wire _60643 = uncoded_block[448] ^ uncoded_block[454];
  wire _60644 = _10352 ^ _60643;
  wire _60645 = _60642 ^ _60644;
  wire _60646 = uncoded_block[473] ^ uncoded_block[481];
  wire _60647 = uncoded_block[485] ^ uncoded_block[512];
  wire _60648 = _60646 ^ _60647;
  wire _60649 = uncoded_block[513] ^ uncoded_block[532];
  wire _60650 = uncoded_block[537] ^ uncoded_block[554];
  wire _60651 = _60649 ^ _60650;
  wire _60652 = _60648 ^ _60651;
  wire _60653 = _60645 ^ _60652;
  wire _60654 = uncoded_block[582] ^ uncoded_block[597];
  wire _60655 = _15239 ^ _60654;
  wire _60656 = uncoded_block[609] ^ uncoded_block[618];
  wire _60657 = uncoded_block[628] ^ uncoded_block[642];
  wire _60658 = _60656 ^ _60657;
  wire _60659 = _60655 ^ _60658;
  wire _60660 = uncoded_block[647] ^ uncoded_block[654];
  wire _60661 = uncoded_block[678] ^ uncoded_block[688];
  wire _60662 = _60660 ^ _60661;
  wire _60663 = uncoded_block[715] ^ uncoded_block[723];
  wire _60664 = _46294 ^ _60663;
  wire _60665 = _60662 ^ _60664;
  wire _60666 = _60659 ^ _60665;
  wire _60667 = _60653 ^ _60666;
  wire _60668 = _60640 ^ _60667;
  wire _60669 = uncoded_block[748] ^ uncoded_block[760];
  wire _60670 = _60669 ^ _6382;
  wire _60671 = uncoded_block[815] ^ uncoded_block[820];
  wire _60672 = _59776 ^ _60671;
  wire _60673 = _60670 ^ _60672;
  wire _60674 = uncoded_block[829] ^ uncoded_block[840];
  wire _60675 = uncoded_block[856] ^ uncoded_block[863];
  wire _60676 = _60674 ^ _60675;
  wire _60677 = uncoded_block[864] ^ uncoded_block[883];
  wire _60678 = _60677 ^ _9960;
  wire _60679 = _60676 ^ _60678;
  wire _60680 = _60673 ^ _60679;
  wire _60681 = uncoded_block[929] ^ uncoded_block[946];
  wire _60682 = _3631 ^ _60681;
  wire _60683 = uncoded_block[972] ^ uncoded_block[992];
  wire _60684 = uncoded_block[1015] ^ uncoded_block[1024];
  wire _60685 = _60683 ^ _60684;
  wire _60686 = _60682 ^ _60685;
  wire _60687 = uncoded_block[1027] ^ uncoded_block[1035];
  wire _60688 = uncoded_block[1039] ^ uncoded_block[1061];
  wire _60689 = _60687 ^ _60688;
  wire _60690 = uncoded_block[1092] ^ uncoded_block[1111];
  wire _60691 = _10569 ^ _60690;
  wire _60692 = _60689 ^ _60691;
  wire _60693 = _60686 ^ _60692;
  wire _60694 = _60680 ^ _60693;
  wire _60695 = uncoded_block[1134] ^ uncoded_block[1139];
  wire _60696 = _46066 ^ _60695;
  wire _60697 = uncoded_block[1158] ^ uncoded_block[1184];
  wire _60698 = uncoded_block[1187] ^ uncoded_block[1194];
  wire _60699 = _60697 ^ _60698;
  wire _60700 = _60696 ^ _60699;
  wire _60701 = uncoded_block[1205] ^ uncoded_block[1210];
  wire _60702 = uncoded_block[1241] ^ uncoded_block[1255];
  wire _60703 = _60701 ^ _60702;
  wire _60704 = uncoded_block[1295] ^ uncoded_block[1311];
  wire _60705 = _52951 ^ _60704;
  wire _60706 = _60703 ^ _60705;
  wire _60707 = _60700 ^ _60706;
  wire _60708 = uncoded_block[1334] ^ uncoded_block[1344];
  wire _60709 = _35389 ^ _60708;
  wire _60710 = uncoded_block[1345] ^ uncoded_block[1356];
  wire _60711 = uncoded_block[1365] ^ uncoded_block[1380];
  wire _60712 = _60710 ^ _60711;
  wire _60713 = _60709 ^ _60712;
  wire _60714 = uncoded_block[1420] ^ uncoded_block[1446];
  wire _60715 = _6596 ^ _60714;
  wire _60716 = uncoded_block[1448] ^ uncoded_block[1469];
  wire _60717 = uncoded_block[1486] ^ uncoded_block[1524];
  wire _60718 = _60716 ^ _60717;
  wire _60719 = _60715 ^ _60718;
  wire _60720 = _60713 ^ _60719;
  wire _60721 = _60707 ^ _60720;
  wire _60722 = _60694 ^ _60721;
  wire _60723 = _60668 ^ _60722;
  wire _60724 = _6647 ^ _9634;
  wire _60725 = uncoded_block[1576] ^ uncoded_block[1605];
  wire _60726 = uncoded_block[1610] ^ uncoded_block[1613];
  wire _60727 = _60725 ^ _60726;
  wire _60728 = _60724 ^ _60727;
  wire _60729 = uncoded_block[1630] ^ uncoded_block[1639];
  wire _60730 = uncoded_block[1647] ^ uncoded_block[1654];
  wire _60731 = _60729 ^ _60730;
  wire _60732 = _5398 ^ _6705;
  wire _60733 = _60731 ^ _60732;
  wire _60734 = _60728 ^ _60733;
  wire _60735 = _47273 ^ uncoded_block[1709];
  wire _60736 = _60734 ^ _60735;
  wire _60737 = _60723 ^ _60736;
  wire _60738 = uncoded_block[7] ^ uncoded_block[21];
  wire _60739 = _21861 ^ _60738;
  wire _60740 = uncoded_block[28] ^ uncoded_block[44];
  wire _60741 = _13539 ^ _60740;
  wire _60742 = _60739 ^ _60741;
  wire _60743 = _10234 ^ _4015;
  wire _60744 = uncoded_block[86] ^ uncoded_block[98];
  wire _60745 = _12438 ^ _60744;
  wire _60746 = _60743 ^ _60745;
  wire _60747 = _60742 ^ _60746;
  wire _60748 = uncoded_block[99] ^ uncoded_block[104];
  wire _60749 = uncoded_block[124] ^ uncoded_block[137];
  wire _60750 = _60748 ^ _60749;
  wire _60751 = uncoded_block[154] ^ uncoded_block[162];
  wire _60752 = _18100 ^ _60751;
  wire _60753 = _60750 ^ _60752;
  wire _60754 = uncoded_block[169] ^ uncoded_block[180];
  wire _60755 = _60754 ^ _944;
  wire _60756 = uncoded_block[186] ^ uncoded_block[196];
  wire _60757 = _60756 ^ _25983;
  wire _60758 = _60755 ^ _60757;
  wire _60759 = _60753 ^ _60758;
  wire _60760 = _60747 ^ _60759;
  wire _60761 = uncoded_block[205] ^ uncoded_block[213];
  wire _60762 = uncoded_block[215] ^ uncoded_block[225];
  wire _60763 = _60761 ^ _60762;
  wire _60764 = uncoded_block[227] ^ uncoded_block[233];
  wire _60765 = uncoded_block[234] ^ uncoded_block[242];
  wire _60766 = _60764 ^ _60765;
  wire _60767 = _60763 ^ _60766;
  wire _60768 = uncoded_block[244] ^ uncoded_block[251];
  wire _60769 = _60768 ^ _10864;
  wire _60770 = uncoded_block[267] ^ uncoded_block[281];
  wire _60771 = _60770 ^ _7446;
  wire _60772 = _60769 ^ _60771;
  wire _60773 = _60767 ^ _60772;
  wire _60774 = uncoded_block[295] ^ uncoded_block[300];
  wire _60775 = _60774 ^ _8052;
  wire _60776 = _1008 ^ _59955;
  wire _60777 = _60775 ^ _60776;
  wire _60778 = uncoded_block[352] ^ uncoded_block[369];
  wire _60779 = _5541 ^ _60778;
  wire _60780 = uncoded_block[382] ^ uncoded_block[387];
  wire _60781 = _16664 ^ _60780;
  wire _60782 = _60779 ^ _60781;
  wire _60783 = _60777 ^ _60782;
  wire _60784 = _60773 ^ _60783;
  wire _60785 = _60760 ^ _60784;
  wire _60786 = _18633 ^ _10340;
  wire _60787 = uncoded_block[401] ^ uncoded_block[412];
  wire _60788 = _60787 ^ _14689;
  wire _60789 = _60786 ^ _60788;
  wire _60790 = uncoded_block[468] ^ uncoded_block[476];
  wire _60791 = _4169 ^ _60790;
  wire _60792 = _1086 ^ _7515;
  wire _60793 = _60791 ^ _60792;
  wire _60794 = _60789 ^ _60793;
  wire _60795 = _6919 ^ _21536;
  wire _60796 = _10376 ^ _2681;
  wire _60797 = _60795 ^ _60796;
  wire _60798 = uncoded_block[526] ^ uncoded_block[543];
  wire _60799 = uncoded_block[571] ^ uncoded_block[577];
  wire _60800 = _60798 ^ _60799;
  wire _60801 = uncoded_block[583] ^ uncoded_block[592];
  wire _60802 = _60801 ^ _1142;
  wire _60803 = _60800 ^ _60802;
  wire _60804 = _60797 ^ _60803;
  wire _60805 = _60794 ^ _60804;
  wire _60806 = uncoded_block[619] ^ uncoded_block[625];
  wire _60807 = _2715 ^ _60806;
  wire _60808 = uncoded_block[627] ^ uncoded_block[642];
  wire _60809 = _60808 ^ _1960;
  wire _60810 = _60807 ^ _60809;
  wire _60811 = uncoded_block[653] ^ uncoded_block[661];
  wire _60812 = _60811 ^ _21113;
  wire _60813 = _4265 ^ _1971;
  wire _60814 = _60812 ^ _60813;
  wire _60815 = _60810 ^ _60814;
  wire _60816 = uncoded_block[693] ^ uncoded_block[700];
  wire _60817 = _60816 ^ _18721;
  wire _60818 = uncoded_block[708] ^ uncoded_block[716];
  wire _60819 = uncoded_block[733] ^ uncoded_block[745];
  wire _60820 = _60818 ^ _60819;
  wire _60821 = _60817 ^ _60820;
  wire _60822 = uncoded_block[761] ^ uncoded_block[773];
  wire _60823 = _60822 ^ _4309;
  wire _60824 = _31539 ^ _60823;
  wire _60825 = _60821 ^ _60824;
  wire _60826 = _60815 ^ _60825;
  wire _60827 = _60805 ^ _60826;
  wire _60828 = _60785 ^ _60827;
  wire _60829 = uncoded_block[796] ^ uncoded_block[802];
  wire _60830 = _2798 ^ _60829;
  wire _60831 = uncoded_block[816] ^ uncoded_block[824];
  wire _60832 = _4322 ^ _60831;
  wire _60833 = _60830 ^ _60832;
  wire _60834 = uncoded_block[846] ^ uncoded_block[858];
  wire _60835 = _15324 ^ _60834;
  wire _60836 = uncoded_block[871] ^ uncoded_block[879];
  wire _60837 = _5069 ^ _60836;
  wire _60838 = _60835 ^ _60837;
  wire _60839 = _60833 ^ _60838;
  wire _60840 = _421 ^ _4358;
  wire _60841 = uncoded_block[915] ^ uncoded_block[921];
  wire _60842 = _9961 ^ _60841;
  wire _60843 = _60840 ^ _60842;
  wire _60844 = uncoded_block[927] ^ uncoded_block[940];
  wire _60845 = uncoded_block[948] ^ uncoded_block[956];
  wire _60846 = _60844 ^ _60845;
  wire _60847 = _59545 ^ _12733;
  wire _60848 = _60846 ^ _60847;
  wire _60849 = _60843 ^ _60848;
  wire _60850 = _60839 ^ _60849;
  wire _60851 = _35704 ^ _8296;
  wire _60852 = uncoded_block[1028] ^ uncoded_block[1034];
  wire _60853 = _5134 ^ _60852;
  wire _60854 = _60851 ^ _60853;
  wire _60855 = _27085 ^ _28256;
  wire _60856 = uncoded_block[1060] ^ uncoded_block[1069];
  wire _60857 = _60856 ^ _6486;
  wire _60858 = _60855 ^ _60857;
  wire _60859 = _60854 ^ _60858;
  wire _60860 = uncoded_block[1100] ^ uncoded_block[1113];
  wire _60861 = _5166 ^ _60860;
  wire _60862 = uncoded_block[1121] ^ uncoded_block[1127];
  wire _60863 = uncoded_block[1130] ^ uncoded_block[1148];
  wire _60864 = _60862 ^ _60863;
  wire _60865 = _60861 ^ _60864;
  wire _60866 = uncoded_block[1186] ^ uncoded_block[1193];
  wire _60867 = _17890 ^ _60866;
  wire _60868 = _44274 ^ _60867;
  wire _60869 = _60865 ^ _60868;
  wire _60870 = _60859 ^ _60869;
  wire _60871 = _60850 ^ _60870;
  wire _60872 = _40903 ^ _2981;
  wire _60873 = _2985 ^ _45037;
  wire _60874 = _60872 ^ _60873;
  wire _60875 = uncoded_block[1264] ^ uncoded_block[1269];
  wire _60876 = _621 ^ _60875;
  wire _60877 = uncoded_block[1271] ^ uncoded_block[1277];
  wire _60878 = _60877 ^ _22657;
  wire _60879 = _60876 ^ _60878;
  wire _60880 = _60874 ^ _60879;
  wire _60881 = uncoded_block[1297] ^ uncoded_block[1302];
  wire _60882 = _4529 ^ _60881;
  wire _60883 = uncoded_block[1315] ^ uncoded_block[1321];
  wire _60884 = _14430 ^ _60883;
  wire _60885 = _60882 ^ _60884;
  wire _60886 = _6578 ^ _9564;
  wire _60887 = uncoded_block[1346] ^ uncoded_block[1352];
  wire _60888 = _60887 ^ _5940;
  wire _60889 = _60886 ^ _60888;
  wire _60890 = _60885 ^ _60889;
  wire _60891 = _60880 ^ _60890;
  wire _60892 = uncoded_block[1373] ^ uncoded_block[1379];
  wire _60893 = _12300 ^ _60892;
  wire _60894 = _688 ^ _5955;
  wire _60895 = _60893 ^ _60894;
  wire _60896 = uncoded_block[1399] ^ uncoded_block[1415];
  wire _60897 = uncoded_block[1417] ^ uncoded_block[1431];
  wire _60898 = _60896 ^ _60897;
  wire _60899 = uncoded_block[1435] ^ uncoded_block[1458];
  wire _60900 = uncoded_block[1462] ^ uncoded_block[1473];
  wire _60901 = _60899 ^ _60900;
  wire _60902 = _60898 ^ _60901;
  wire _60903 = _60895 ^ _60902;
  wire _60904 = uncoded_block[1476] ^ uncoded_block[1492];
  wire _60905 = _60904 ^ _6643;
  wire _60906 = _56921 ^ _5350;
  wire _60907 = _60905 ^ _60906;
  wire _60908 = uncoded_block[1543] ^ uncoded_block[1554];
  wire _60909 = _60908 ^ _4640;
  wire _60910 = _58314 ^ _46487;
  wire _60911 = _60909 ^ _60910;
  wire _60912 = _60907 ^ _60911;
  wire _60913 = _60903 ^ _60912;
  wire _60914 = _60891 ^ _60913;
  wire _60915 = _60871 ^ _60914;
  wire _60916 = _60828 ^ _60915;
  wire _60917 = uncoded_block[1593] ^ uncoded_block[1598];
  wire _60918 = _60917 ^ _4660;
  wire _60919 = uncoded_block[1625] ^ uncoded_block[1631];
  wire _60920 = _36256 ^ _60919;
  wire _60921 = _60918 ^ _60920;
  wire _60922 = uncoded_block[1642] ^ uncoded_block[1666];
  wire _60923 = _3948 ^ _60922;
  wire _60924 = uncoded_block[1667] ^ uncoded_block[1675];
  wire _60925 = _60924 ^ _39083;
  wire _60926 = _60923 ^ _60925;
  wire _60927 = _60921 ^ _60926;
  wire _60928 = _50710 ^ uncoded_block[1718];
  wire _60929 = _60927 ^ _60928;
  wire _60930 = _60916 ^ _60929;
  wire _60931 = uncoded_block[4] ^ uncoded_block[18];
  wire _60932 = _60931 ^ _28752;
  wire _60933 = uncoded_block[47] ^ uncoded_block[69];
  wire _60934 = _60933 ^ _10246;
  wire _60935 = _60932 ^ _60934;
  wire _60936 = _44430 ^ _57813;
  wire _60937 = uncoded_block[140] ^ uncoded_block[148];
  wire _60938 = _2498 ^ _60937;
  wire _60939 = _60936 ^ _60938;
  wire _60940 = _60935 ^ _60939;
  wire _60941 = uncoded_block[166] ^ uncoded_block[173];
  wire _60942 = uncoded_block[178] ^ uncoded_block[183];
  wire _60943 = _60941 ^ _60942;
  wire _60944 = uncoded_block[215] ^ uncoded_block[228];
  wire _60945 = _4780 ^ _60944;
  wire _60946 = _60943 ^ _60945;
  wire _60947 = uncoded_block[256] ^ uncoded_block[267];
  wire _60948 = _6182 ^ _60947;
  wire _60949 = uncoded_block[271] ^ uncoded_block[295];
  wire _60950 = _60949 ^ _28067;
  wire _60951 = _60948 ^ _60950;
  wire _60952 = _60946 ^ _60951;
  wire _60953 = _60940 ^ _60952;
  wire _60954 = uncoded_block[327] ^ uncoded_block[349];
  wire _60955 = _3341 ^ _60954;
  wire _60956 = _2602 ^ _57854;
  wire _60957 = _60955 ^ _60956;
  wire _60958 = uncoded_block[387] ^ uncoded_block[399];
  wire _60959 = uncoded_block[415] ^ uncoded_block[422];
  wire _60960 = _60958 ^ _60959;
  wire _60961 = uncoded_block[447] ^ uncoded_block[457];
  wire _60962 = _12015 ^ _60961;
  wire _60963 = _60960 ^ _60962;
  wire _60964 = _60957 ^ _60963;
  wire _60965 = uncoded_block[460] ^ uncoded_block[484];
  wire _60966 = uncoded_block[492] ^ uncoded_block[499];
  wire _60967 = _60965 ^ _60966;
  wire _60968 = uncoded_block[501] ^ uncoded_block[508];
  wire _60969 = uncoded_block[513] ^ uncoded_block[525];
  wire _60970 = _60968 ^ _60969;
  wire _60971 = _60967 ^ _60970;
  wire _60972 = uncoded_block[526] ^ uncoded_block[541];
  wire _60973 = uncoded_block[552] ^ uncoded_block[568];
  wire _60974 = _60972 ^ _60973;
  wire _60975 = _6945 ^ _16727;
  wire _60976 = _60974 ^ _60975;
  wire _60977 = _60971 ^ _60976;
  wire _60978 = _60964 ^ _60977;
  wire _60979 = _60953 ^ _60978;
  wire _60980 = uncoded_block[599] ^ uncoded_block[625];
  wire _60981 = uncoded_block[651] ^ uncoded_block[659];
  wire _60982 = _60980 ^ _60981;
  wire _60983 = uncoded_block[666] ^ uncoded_block[675];
  wire _60984 = _60983 ^ _60661;
  wire _60985 = _60982 ^ _60984;
  wire _60986 = uncoded_block[711] ^ uncoded_block[739];
  wire _60987 = _60986 ^ _5699;
  wire _60988 = uncoded_block[754] ^ uncoded_block[765];
  wire _60989 = _60988 ^ _4308;
  wire _60990 = _60987 ^ _60989;
  wire _60991 = _60985 ^ _60990;
  wire _60992 = uncoded_block[789] ^ uncoded_block[802];
  wire _60993 = _2794 ^ _60992;
  wire _60994 = uncoded_block[818] ^ uncoded_block[840];
  wire _60995 = _60994 ^ _25710;
  wire _60996 = _60993 ^ _60995;
  wire _60997 = uncoded_block[859] ^ uncoded_block[891];
  wire _60998 = _21631 ^ _60997;
  wire _60999 = uncoded_block[895] ^ uncoded_block[902];
  wire _61000 = uncoded_block[924] ^ uncoded_block[941];
  wire _61001 = _60999 ^ _61000;
  wire _61002 = _60998 ^ _61001;
  wire _61003 = _60996 ^ _61002;
  wire _61004 = _60991 ^ _61003;
  wire _61005 = uncoded_block[950] ^ uncoded_block[983];
  wire _61006 = uncoded_block[985] ^ uncoded_block[997];
  wire _61007 = _61005 ^ _61006;
  wire _61008 = uncoded_block[1004] ^ uncoded_block[1017];
  wire _61009 = _61008 ^ _48257;
  wire _61010 = _61007 ^ _61009;
  wire _61011 = _37755 ^ _59142;
  wire _61012 = _13316 ^ _15407;
  wire _61013 = _61011 ^ _61012;
  wire _61014 = _61010 ^ _61013;
  wire _61015 = uncoded_block[1140] ^ uncoded_block[1146];
  wire _61016 = _61015 ^ _22627;
  wire _61017 = uncoded_block[1172] ^ uncoded_block[1193];
  wire _61018 = uncoded_block[1195] ^ uncoded_block[1220];
  wire _61019 = _61017 ^ _61018;
  wire _61020 = _61016 ^ _61019;
  wire _61021 = uncoded_block[1241] ^ uncoded_block[1249];
  wire _61022 = _14921 ^ _61021;
  wire _61023 = uncoded_block[1258] ^ uncoded_block[1270];
  wire _61024 = uncoded_block[1289] ^ uncoded_block[1301];
  wire _61025 = _61023 ^ _61024;
  wire _61026 = _61022 ^ _61025;
  wire _61027 = _61020 ^ _61026;
  wire _61028 = _61014 ^ _61027;
  wire _61029 = _61004 ^ _61028;
  wire _61030 = _60979 ^ _61029;
  wire _61031 = uncoded_block[1317] ^ uncoded_block[1335];
  wire _61032 = _648 ^ _61031;
  wire _61033 = uncoded_block[1348] ^ uncoded_block[1359];
  wire _61034 = uncoded_block[1372] ^ uncoded_block[1381];
  wire _61035 = _61033 ^ _61034;
  wire _61036 = _61032 ^ _61035;
  wire _61037 = uncoded_block[1404] ^ uncoded_block[1417];
  wire _61038 = _61037 ^ _1526;
  wire _61039 = _21323 ^ _4590;
  wire _61040 = _61038 ^ _61039;
  wire _61041 = _61036 ^ _61040;
  wire _61042 = uncoded_block[1447] ^ uncoded_block[1457];
  wire _61043 = uncoded_block[1475] ^ uncoded_block[1483];
  wire _61044 = _61042 ^ _61043;
  wire _61045 = uncoded_block[1488] ^ uncoded_block[1509];
  wire _61046 = _27184 ^ _61045;
  wire _61047 = _61044 ^ _61046;
  wire _61048 = uncoded_block[1511] ^ uncoded_block[1519];
  wire _61049 = uncoded_block[1527] ^ uncoded_block[1535];
  wire _61050 = _61048 ^ _61049;
  wire _61051 = uncoded_block[1594] ^ uncoded_block[1602];
  wire _61052 = uncoded_block[1610] ^ uncoded_block[1627];
  wire _61053 = _61051 ^ _61052;
  wire _61054 = _61050 ^ _61053;
  wire _61055 = _61047 ^ _61054;
  wire _61056 = _61041 ^ _61055;
  wire _61057 = uncoded_block[1629] ^ uncoded_block[1637];
  wire _61058 = uncoded_block[1656] ^ uncoded_block[1670];
  wire _61059 = _61057 ^ _61058;
  wire _61060 = _6059 ^ _33862;
  wire _61061 = _61059 ^ _61060;
  wire _61062 = _7935 ^ _6072;
  wire _61063 = _61062 ^ uncoded_block[1722];
  wire _61064 = _61061 ^ _61063;
  wire _61065 = _61056 ^ _61064;
  wire _61066 = _61030 ^ _61065;
  wire _61067 = uncoded_block[12] ^ uncoded_block[24];
  wire _61068 = _3993 ^ _61067;
  wire _61069 = _19965 ^ _19006;
  wire _61070 = _61068 ^ _61069;
  wire _61071 = _12428 ^ _28757;
  wire _61072 = _6742 ^ _42215;
  wire _61073 = _61071 ^ _61072;
  wire _61074 = _61070 ^ _61073;
  wire _61075 = _901 ^ _58993;
  wire _61076 = _51123 ^ _57813;
  wire _61077 = _61075 ^ _61076;
  wire _61078 = uncoded_block[131] ^ uncoded_block[138];
  wire _61079 = _61078 ^ _42602;
  wire _61080 = _57816 ^ _61079;
  wire _61081 = _61077 ^ _61080;
  wire _61082 = _61074 ^ _61081;
  wire _61083 = _6785 ^ _14092;
  wire _61084 = _61083 ^ _57827;
  wire _61085 = _963 ^ _33088;
  wire _61086 = _57830 ^ _61085;
  wire _61087 = _61084 ^ _61086;
  wire _61088 = uncoded_block[246] ^ uncoded_block[251];
  wire _61089 = uncoded_block[254] ^ uncoded_block[262];
  wire _61090 = _61088 ^ _61089;
  wire _61091 = _14122 ^ _43681;
  wire _61092 = _61090 ^ _61091;
  wire _61093 = uncoded_block[284] ^ uncoded_block[294];
  wire _61094 = _61093 ^ _4110;
  wire _61095 = uncoded_block[299] ^ uncoded_block[305];
  wire _61096 = _61095 ^ _146;
  wire _61097 = _61094 ^ _61096;
  wire _61098 = _61092 ^ _61097;
  wire _61099 = _61087 ^ _61098;
  wire _61100 = _61082 ^ _61099;
  wire _61101 = uncoded_block[317] ^ uncoded_block[323];
  wire _61102 = _61101 ^ _5534;
  wire _61103 = _8646 ^ _4129;
  wire _61104 = _61102 ^ _61103;
  wire _61105 = uncoded_block[347] ^ uncoded_block[356];
  wire _61106 = _61105 ^ _57853;
  wire _61107 = _57854 ^ _12005;
  wire _61108 = _61106 ^ _61107;
  wire _61109 = _61104 ^ _61108;
  wire _61110 = _1847 ^ _37991;
  wire _61111 = _13650 ^ _59046;
  wire _61112 = _61110 ^ _61111;
  wire _61113 = _23349 ^ _13662;
  wire _61114 = uncoded_block[466] ^ uncoded_block[484];
  wire _61115 = uncoded_block[486] ^ uncoded_block[497];
  wire _61116 = _61114 ^ _61115;
  wire _61117 = _61113 ^ _61116;
  wire _61118 = _61112 ^ _61117;
  wire _61119 = _61109 ^ _61118;
  wire _61120 = _4905 ^ _15725;
  wire _61121 = _27369 ^ _57876;
  wire _61122 = _61120 ^ _61121;
  wire _61123 = _20602 ^ _57878;
  wire _61124 = _5628 ^ _25631;
  wire _61125 = _61123 ^ _61124;
  wire _61126 = _61122 ^ _61125;
  wire _61127 = _39617 ^ _4941;
  wire _61128 = _55572 ^ _18222;
  wire _61129 = _61127 ^ _61128;
  wire _61130 = uncoded_block[591] ^ uncoded_block[598];
  wire _61131 = _61130 ^ _274;
  wire _61132 = _56482 ^ _57666;
  wire _61133 = _61131 ^ _61132;
  wire _61134 = _61129 ^ _61133;
  wire _61135 = _61126 ^ _61134;
  wire _61136 = _61119 ^ _61135;
  wire _61137 = _61100 ^ _61136;
  wire _61138 = uncoded_block[638] ^ uncoded_block[645];
  wire _61139 = _61138 ^ _19177;
  wire _61140 = _4261 ^ _9886;
  wire _61141 = _61139 ^ _61140;
  wire _61142 = uncoded_block[700] ^ uncoded_block[707];
  wire _61143 = _2755 ^ _61142;
  wire _61144 = _57899 ^ _61143;
  wire _61145 = _61141 ^ _61144;
  wire _61146 = _340 ^ _4287;
  wire _61147 = _61146 ^ _59766;
  wire _61148 = uncoded_block[745] ^ uncoded_block[751];
  wire _61149 = _61148 ^ _7015;
  wire _61150 = uncoded_block[758] ^ uncoded_block[768];
  wire _61151 = _61150 ^ _57912;
  wire _61152 = _61149 ^ _61151;
  wire _61153 = _61147 ^ _61152;
  wire _61154 = _61145 ^ _61153;
  wire _61155 = uncoded_block[789] ^ uncoded_block[796];
  wire _61156 = _61155 ^ _2801;
  wire _61157 = _3582 ^ _18288;
  wire _61158 = _61156 ^ _61157;
  wire _61159 = _1256 ^ _2821;
  wire _61160 = uncoded_block[858] ^ uncoded_block[867];
  wire _61161 = _61160 ^ _15826;
  wire _61162 = _61159 ^ _61161;
  wire _61163 = _61158 ^ _61162;
  wire _61164 = _35678 ^ _5085;
  wire _61165 = _6425 ^ _16313;
  wire _61166 = _61164 ^ _61165;
  wire _61167 = uncoded_block[924] ^ uncoded_block[931];
  wire _61168 = _41238 ^ _61167;
  wire _61169 = uncoded_block[950] ^ uncoded_block[957];
  wire _61170 = _2083 ^ _61169;
  wire _61171 = _61168 ^ _61170;
  wire _61172 = _61166 ^ _61171;
  wire _61173 = _61163 ^ _61172;
  wire _61174 = _61154 ^ _61173;
  wire _61175 = uncoded_block[963] ^ uncoded_block[968];
  wire _61176 = _61175 ^ _37341;
  wire _61177 = uncoded_block[980] ^ uncoded_block[997];
  wire _61178 = _5114 ^ _61177;
  wire _61179 = _61176 ^ _61178;
  wire _61180 = uncoded_block[999] ^ uncoded_block[1009];
  wire _61181 = _61180 ^ _1338;
  wire _61182 = _48255 ^ _6478;
  wire _61183 = _61181 ^ _61182;
  wire _61184 = _61179 ^ _61183;
  wire _61185 = uncoded_block[1057] ^ uncoded_block[1067];
  wire _61186 = _4430 ^ _61185;
  wire _61187 = uncoded_block[1070] ^ uncoded_block[1078];
  wire _61188 = _61187 ^ _14366;
  wire _61189 = _61186 ^ _61188;
  wire _61190 = _57955 ^ _57959;
  wire _61191 = _61189 ^ _61190;
  wire _61192 = _61184 ^ _61191;
  wire _61193 = uncoded_block[1133] ^ uncoded_block[1146];
  wire _61194 = _61193 ^ _1401;
  wire _61195 = _19330 ^ _49385;
  wire _61196 = _61194 ^ _61195;
  wire _61197 = uncoded_block[1178] ^ uncoded_block[1192];
  wire _61198 = _27111 ^ _61197;
  wire _61199 = uncoded_block[1193] ^ uncoded_block[1214];
  wire _61200 = _61199 ^ _27912;
  wire _61201 = _61198 ^ _61200;
  wire _61202 = _61196 ^ _61201;
  wire _61203 = uncoded_block[1297] ^ uncoded_block[1308];
  wire _61204 = _40925 ^ _61203;
  wire _61205 = _30800 ^ _5926;
  wire _61206 = _61204 ^ _61205;
  wire _61207 = _57976 ^ _61206;
  wire _61208 = _61202 ^ _61207;
  wire _61209 = _61192 ^ _61208;
  wire _61210 = _61174 ^ _61209;
  wire _61211 = _61137 ^ _61210;
  wire _61212 = _3029 ^ _5256;
  wire _61213 = _61212 ^ _57989;
  wire _61214 = uncoded_block[1348] ^ uncoded_block[1353];
  wire _61215 = _61214 ^ _673;
  wire _61216 = _3045 ^ _57994;
  wire _61217 = _61215 ^ _61216;
  wire _61218 = _61213 ^ _61217;
  wire _61219 = uncoded_block[1387] ^ uncoded_block[1398];
  wire _61220 = _11781 ^ _61219;
  wire _61221 = _10678 ^ _32942;
  wire _61222 = _61220 ^ _61221;
  wire _61223 = _8443 ^ _712;
  wire _61224 = _54518 ^ _719;
  wire _61225 = _61223 ^ _61224;
  wire _61226 = _61222 ^ _61225;
  wire _61227 = _61218 ^ _61226;
  wire _61228 = _9037 ^ _19411;
  wire _61229 = _16479 ^ _58943;
  wire _61230 = _61228 ^ _61229;
  wire _61231 = _11264 ^ _15002;
  wire _61232 = _26321 ^ _23194;
  wire _61233 = _61231 ^ _61232;
  wire _61234 = _61230 ^ _61233;
  wire _61235 = _44372 ^ _16025;
  wire _61236 = _58019 ^ _61235;
  wire _61237 = _42829 ^ _813;
  wire _61238 = uncoded_block[1651] ^ uncoded_block[1662];
  wire _61239 = _36263 ^ _61238;
  wire _61240 = _61237 ^ _61239;
  wire _61241 = _61236 ^ _61240;
  wire _61242 = _61234 ^ _61241;
  wire _61243 = _61227 ^ _61242;
  wire _61244 = _22303 ^ _58034;
  wire _61245 = _61244 ^ _58038;
  wire _61246 = _11327 ^ _21400;
  wire _61247 = _22316 ^ uncoded_block[1721];
  wire _61248 = _61246 ^ _61247;
  wire _61249 = _61245 ^ _61248;
  wire _61250 = _61243 ^ _61249;
  wire _61251 = _61211 ^ _61250;
  wire _61252 = uncoded_block[3] ^ uncoded_block[19];
  wire _61253 = _61252 ^ _18549;
  wire _61254 = uncoded_block[53] ^ uncoded_block[61];
  wire _61255 = _3230 ^ _61254;
  wire _61256 = _61253 ^ _61255;
  wire _61257 = _16089 ^ _6122;
  wire _61258 = uncoded_block[128] ^ uncoded_block[146];
  wire _61259 = _10821 ^ _61258;
  wire _61260 = _61257 ^ _61259;
  wire _61261 = _61256 ^ _61260;
  wire _61262 = uncoded_block[167] ^ uncoded_block[174];
  wire _61263 = _61262 ^ _4773;
  wire _61264 = _6800 ^ _11943;
  wire _61265 = _61263 ^ _61264;
  wire _61266 = uncoded_block[225] ^ uncoded_block[243];
  wire _61267 = _61266 ^ _30548;
  wire _61268 = uncoded_block[275] ^ uncoded_block[280];
  wire _61269 = _61268 ^ _994;
  wire _61270 = _61267 ^ _61269;
  wire _61271 = _61265 ^ _61270;
  wire _61272 = _61261 ^ _61271;
  wire _61273 = uncoded_block[307] ^ uncoded_block[332];
  wire _61274 = _24216 ^ _61273;
  wire _61275 = _61274 ^ _22875;
  wire _61276 = uncoded_block[348] ^ uncoded_block[384];
  wire _61277 = uncoded_block[385] ^ uncoded_block[393];
  wire _61278 = _61276 ^ _61277;
  wire _61279 = uncoded_block[408] ^ uncoded_block[432];
  wire _61280 = _61279 ^ _10352;
  wire _61281 = _61278 ^ _61280;
  wire _61282 = _61275 ^ _61281;
  wire _61283 = _25601 ^ _26495;
  wire _61284 = uncoded_block[466] ^ uncoded_block[481];
  wire _61285 = _8105 ^ _61284;
  wire _61286 = _61283 ^ _61285;
  wire _61287 = uncoded_block[501] ^ uncoded_block[509];
  wire _61288 = _61287 ^ _20598;
  wire _61289 = uncoded_block[533] ^ uncoded_block[541];
  wire _61290 = uncoded_block[550] ^ uncoded_block[557];
  wire _61291 = _61289 ^ _61290;
  wire _61292 = _61288 ^ _61291;
  wire _61293 = _61286 ^ _61292;
  wire _61294 = _61282 ^ _61293;
  wire _61295 = _61272 ^ _61294;
  wire _61296 = uncoded_block[578] ^ uncoded_block[585];
  wire _61297 = _6942 ^ _61296;
  wire _61298 = uncoded_block[588] ^ uncoded_block[611];
  wire _61299 = uncoded_block[612] ^ uncoded_block[619];
  wire _61300 = _61298 ^ _61299;
  wire _61301 = _61297 ^ _61300;
  wire _61302 = _4255 ^ _296;
  wire _61303 = _60523 ^ _36442;
  wire _61304 = _61302 ^ _61303;
  wire _61305 = _61301 ^ _61304;
  wire _61306 = uncoded_block[680] ^ uncoded_block[699];
  wire _61307 = _61306 ^ _4996;
  wire _61308 = uncoded_block[714] ^ uncoded_block[731];
  wire _61309 = _61308 ^ _3549;
  wire _61310 = _61307 ^ _61309;
  wire _61311 = uncoded_block[746] ^ uncoded_block[779];
  wire _61312 = uncoded_block[783] ^ uncoded_block[794];
  wire _61313 = _61311 ^ _61312;
  wire _61314 = uncoded_block[810] ^ uncoded_block[822];
  wire _61315 = _389 ^ _61314;
  wire _61316 = _61313 ^ _61315;
  wire _61317 = _61310 ^ _61316;
  wire _61318 = _61305 ^ _61317;
  wire _61319 = uncoded_block[839] ^ uncoded_block[857];
  wire _61320 = _1253 ^ _61319;
  wire _61321 = uncoded_block[877] ^ uncoded_block[889];
  wire _61322 = _2828 ^ _61321;
  wire _61323 = _61320 ^ _61322;
  wire _61324 = _56807 ^ _2843;
  wire _61325 = uncoded_block[958] ^ uncoded_block[974];
  wire _61326 = _7665 ^ _61325;
  wire _61327 = _61324 ^ _61326;
  wire _61328 = _61323 ^ _61327;
  wire _61329 = _2882 ^ _4402;
  wire _61330 = uncoded_block[1001] ^ uncoded_block[1008];
  wire _61331 = uncoded_block[1015] ^ uncoded_block[1036];
  wire _61332 = _61330 ^ _61331;
  wire _61333 = _61329 ^ _61332;
  wire _61334 = uncoded_block[1041] ^ uncoded_block[1049];
  wire _61335 = _61334 ^ _519;
  wire _61336 = uncoded_block[1061] ^ uncoded_block[1072];
  wire _61337 = uncoded_block[1086] ^ uncoded_block[1097];
  wire _61338 = _61336 ^ _61337;
  wire _61339 = _61335 ^ _61338;
  wire _61340 = _61333 ^ _61339;
  wire _61341 = _61328 ^ _61340;
  wire _61342 = _61318 ^ _61341;
  wire _61343 = _61295 ^ _61342;
  wire _61344 = uncoded_block[1100] ^ uncoded_block[1122];
  wire _61345 = _543 ^ _61344;
  wire _61346 = uncoded_block[1143] ^ uncoded_block[1152];
  wire _61347 = _61346 ^ _6507;
  wire _61348 = _61345 ^ _61347;
  wire _61349 = _43884 ^ _3742;
  wire _61350 = _9508 ^ _620;
  wire _61351 = _61349 ^ _61350;
  wire _61352 = _61348 ^ _61351;
  wire _61353 = uncoded_block[1268] ^ uncoded_block[1276];
  wire _61354 = _61353 ^ _1465;
  wire _61355 = _26263 ^ _61354;
  wire _61356 = uncoded_block[1286] ^ uncoded_block[1304];
  wire _61357 = uncoded_block[1313] ^ uncoded_block[1330];
  wire _61358 = _61356 ^ _61357;
  wire _61359 = uncoded_block[1344] ^ uncoded_block[1357];
  wire _61360 = uncoded_block[1365] ^ uncoded_block[1370];
  wire _61361 = _61359 ^ _61360;
  wire _61362 = _61358 ^ _61361;
  wire _61363 = _61355 ^ _61362;
  wire _61364 = _61352 ^ _61363;
  wire _61365 = uncoded_block[1371] ^ uncoded_block[1382];
  wire _61366 = uncoded_block[1383] ^ uncoded_block[1413];
  wire _61367 = _61365 ^ _61366;
  wire _61368 = _55746 ^ _2311;
  wire _61369 = _61367 ^ _61368;
  wire _61370 = uncoded_block[1448] ^ uncoded_block[1455];
  wire _61371 = _2319 ^ _61370;
  wire _61372 = uncoded_block[1460] ^ uncoded_block[1475];
  wire _61373 = _61372 ^ _1558;
  wire _61374 = _61371 ^ _61373;
  wire _61375 = _61369 ^ _61374;
  wire _61376 = uncoded_block[1485] ^ uncoded_block[1510];
  wire _61377 = _61376 ^ _26321;
  wire _61378 = uncoded_block[1527] ^ uncoded_block[1537];
  wire _61379 = _61378 ^ _1589;
  wire _61380 = _61377 ^ _61379;
  wire _61381 = uncoded_block[1547] ^ uncoded_block[1578];
  wire _61382 = _61381 ^ _2383;
  wire _61383 = uncoded_block[1605] ^ uncoded_block[1623];
  wire _61384 = uncoded_block[1635] ^ uncoded_block[1653];
  wire _61385 = _61383 ^ _61384;
  wire _61386 = _61382 ^ _61385;
  wire _61387 = _61380 ^ _61386;
  wire _61388 = _61375 ^ _61387;
  wire _61389 = _61364 ^ _61388;
  wire _61390 = _12960 ^ _17040;
  wire _61391 = uncoded_block[1698] ^ uncoded_block[1707];
  wire _61392 = _42191 ^ _61391;
  wire _61393 = _61390 ^ _61392;
  wire _61394 = _61393 ^ uncoded_block[1715];
  wire _61395 = _61389 ^ _61394;
  wire _61396 = _61343 ^ _61395;
  wire _61397 = uncoded_block[0] ^ uncoded_block[18];
  wire _61398 = _61397 ^ _2458;
  wire _61399 = uncoded_block[31] ^ uncoded_block[42];
  wire _61400 = _3224 ^ _61399;
  wire _61401 = _61398 ^ _61400;
  wire _61402 = uncoded_block[43] ^ uncoded_block[52];
  wire _61403 = _61402 ^ _6106;
  wire _61404 = _6107 ^ _6750;
  wire _61405 = _61403 ^ _61404;
  wire _61406 = _61401 ^ _61405;
  wire _61407 = uncoded_block[85] ^ uncoded_block[96];
  wire _61408 = _61407 ^ _59416;
  wire _61409 = _54 ^ _4042;
  wire _61410 = _61408 ^ _61409;
  wire _61411 = uncoded_block[147] ^ uncoded_block[153];
  wire _61412 = _7999 ^ _61411;
  wire _61413 = _46182 ^ _938;
  wire _61414 = _61412 ^ _61413;
  wire _61415 = _61410 ^ _61414;
  wire _61416 = _61406 ^ _61415;
  wire _61417 = _14092 ^ _4776;
  wire _61418 = uncoded_block[216] ^ uncoded_block[223];
  wire _61419 = _6805 ^ _61418;
  wire _61420 = _61417 ^ _61419;
  wire _61421 = uncoded_block[226] ^ uncoded_block[234];
  wire _61422 = _61421 ^ _57002;
  wire _61423 = uncoded_block[260] ^ uncoded_block[272];
  wire _61424 = _23746 ^ _61423;
  wire _61425 = _61422 ^ _61424;
  wire _61426 = _61420 ^ _61425;
  wire _61427 = uncoded_block[286] ^ uncoded_block[294];
  wire _61428 = _10303 ^ _61427;
  wire _61429 = _61428 ^ _24681;
  wire _61430 = uncoded_block[334] ^ uncoded_block[347];
  wire _61431 = _3341 ^ _61430;
  wire _61432 = _2601 ^ _13093;
  wire _61433 = _61431 ^ _61432;
  wire _61434 = _61429 ^ _61433;
  wire _61435 = _61426 ^ _61434;
  wire _61436 = _61416 ^ _61435;
  wire _61437 = uncoded_block[373] ^ uncoded_block[385];
  wire _61438 = _61437 ^ _7487;
  wire _61439 = _11476 ^ _14690;
  wire _61440 = _61438 ^ _61439;
  wire _61441 = uncoded_block[468] ^ uncoded_block[484];
  wire _61442 = uncoded_block[487] ^ uncoded_block[494];
  wire _61443 = _61441 ^ _61442;
  wire _61444 = _59465 ^ _61443;
  wire _61445 = _61440 ^ _61444;
  wire _61446 = _1887 ^ _13152;
  wire _61447 = _61446 ^ _37241;
  wire _61448 = uncoded_block[578] ^ uncoded_block[590];
  wire _61449 = _13697 ^ _61448;
  wire _61450 = _8138 ^ _61449;
  wire _61451 = _61447 ^ _61450;
  wire _61452 = _61445 ^ _61451;
  wire _61453 = _8148 ^ _59489;
  wire _61454 = uncoded_block[607] ^ uncoded_block[615];
  wire _61455 = _61454 ^ _31924;
  wire _61456 = _61453 ^ _61455;
  wire _61457 = uncoded_block[636] ^ uncoded_block[644];
  wire _61458 = _36847 ^ _61457;
  wire _61459 = uncoded_block[676] ^ uncoded_block[682];
  wire _61460 = _17745 ^ _61459;
  wire _61461 = _61458 ^ _61460;
  wire _61462 = _61456 ^ _61461;
  wire _61463 = uncoded_block[710] ^ uncoded_block[721];
  wire _61464 = _61463 ^ _4283;
  wire _61465 = _59760 ^ _61464;
  wire _61466 = _23870 ^ _10464;
  wire _61467 = uncoded_block[753] ^ uncoded_block[757];
  wire _61468 = uncoded_block[758] ^ uncoded_block[780];
  wire _61469 = _61467 ^ _61468;
  wire _61470 = _61466 ^ _61469;
  wire _61471 = _61465 ^ _61470;
  wire _61472 = _61462 ^ _61471;
  wire _61473 = _61452 ^ _61472;
  wire _61474 = _61436 ^ _61473;
  wire _61475 = uncoded_block[783] ^ uncoded_block[796];
  wire _61476 = _61475 ^ _16791;
  wire _61477 = uncoded_block[829] ^ uncoded_block[841];
  wire _61478 = _57408 ^ _61477;
  wire _61479 = _61476 ^ _61478;
  wire _61480 = uncoded_block[850] ^ uncoded_block[858];
  wire _61481 = _61480 ^ _57922;
  wire _61482 = uncoded_block[886] ^ uncoded_block[896];
  wire _61483 = _4347 ^ _61482;
  wire _61484 = _61481 ^ _61483;
  wire _61485 = _61479 ^ _61484;
  wire _61486 = _20704 ^ _10508;
  wire _61487 = _19251 ^ _24832;
  wire _61488 = _61486 ^ _61487;
  wire _61489 = _1300 ^ _57120;
  wire _61490 = uncoded_block[966] ^ uncoded_block[973];
  wire _61491 = _61490 ^ _5118;
  wire _61492 = _61489 ^ _61491;
  wire _61493 = _61488 ^ _61492;
  wire _61494 = _61485 ^ _61493;
  wire _61495 = uncoded_block[1001] ^ uncoded_block[1017];
  wire _61496 = _12737 ^ _61495;
  wire _61497 = _7108 ^ _10564;
  wire _61498 = _61496 ^ _61497;
  wire _61499 = _23062 ^ _13307;
  wire _61500 = uncoded_block[1085] ^ uncoded_block[1089];
  wire _61501 = _530 ^ _61500;
  wire _61502 = _61499 ^ _61501;
  wire _61503 = _61498 ^ _61502;
  wire _61504 = uncoded_block[1102] ^ uncoded_block[1106];
  wire _61505 = _61504 ^ _57147;
  wire _61506 = uncoded_block[1122] ^ uncoded_block[1137];
  wire _61507 = _61506 ^ _565;
  wire _61508 = _61505 ^ _61507;
  wire _61509 = uncoded_block[1155] ^ uncoded_block[1176];
  wire _61510 = _61509 ^ _6519;
  wire _61511 = uncoded_block[1183] ^ uncoded_block[1197];
  wire _61512 = _61511 ^ _43135;
  wire _61513 = _61510 ^ _61512;
  wire _61514 = _61508 ^ _61513;
  wire _61515 = _61503 ^ _61514;
  wire _61516 = _61494 ^ _61515;
  wire _61517 = uncoded_block[1215] ^ uncoded_block[1221];
  wire _61518 = _23544 ^ _61517;
  wire _61519 = _61518 ^ _46798;
  wire _61520 = uncoded_block[1292] ^ uncoded_block[1305];
  wire _61521 = _12834 ^ _61520;
  wire _61522 = _59589 ^ _61521;
  wire _61523 = _61519 ^ _61522;
  wire _61524 = _3812 ^ _47945;
  wire _61525 = uncoded_block[1336] ^ uncoded_block[1358];
  wire _61526 = _61525 ^ _16444;
  wire _61527 = _61524 ^ _61526;
  wire _61528 = uncoded_block[1372] ^ uncoded_block[1380];
  wire _61529 = _21762 ^ _61528;
  wire _61530 = uncoded_block[1387] ^ uncoded_block[1403];
  wire _61531 = _6596 ^ _61530;
  wire _61532 = _61529 ^ _61531;
  wire _61533 = _61527 ^ _61532;
  wire _61534 = _61523 ^ _61533;
  wire _61535 = _13420 ^ _5962;
  wire _61536 = _9021 ^ _9025;
  wire _61537 = _61535 ^ _61536;
  wire _61538 = _26763 ^ _24528;
  wire _61539 = _39034 ^ _59624;
  wire _61540 = _61538 ^ _61539;
  wire _61541 = _61537 ^ _61540;
  wire _61542 = _11813 ^ _13973;
  wire _61543 = uncoded_block[1521] ^ uncoded_block[1529];
  wire _61544 = _61543 ^ _3905;
  wire _61545 = _61542 ^ _61544;
  wire _61546 = uncoded_block[1545] ^ uncoded_block[1568];
  wire _61547 = uncoded_block[1581] ^ uncoded_block[1587];
  wire _61548 = _61546 ^ _61547;
  wire _61549 = _61548 ^ _9643;
  wire _61550 = _61545 ^ _61549;
  wire _61551 = _61541 ^ _61550;
  wire _61552 = _61534 ^ _61551;
  wire _61553 = _61516 ^ _61552;
  wire _61554 = _61474 ^ _61553;
  wire _61555 = uncoded_block[1618] ^ uncoded_block[1630];
  wire _61556 = _3154 ^ _61555;
  wire _61557 = uncoded_block[1633] ^ uncoded_block[1648];
  wire _61558 = _61557 ^ _4677;
  wire _61559 = _61556 ^ _61558;
  wire _61560 = uncoded_block[1666] ^ uncoded_block[1684];
  wire _61561 = _22761 ^ _61560;
  wire _61562 = uncoded_block[1685] ^ uncoded_block[1694];
  wire _61563 = _61562 ^ _35477;
  wire _61564 = _61561 ^ _61563;
  wire _61565 = _61559 ^ _61564;
  wire _61566 = _61565 ^ uncoded_block[1706];
  wire _61567 = _61554 ^ _61566;
  wire _61568 = uncoded_block[9] ^ uncoded_block[28];
  wire _61569 = uncoded_block[30] ^ uncoded_block[36];
  wire _61570 = _61568 ^ _61569;
  wire _61571 = uncoded_block[41] ^ uncoded_block[55];
  wire _61572 = _61571 ^ _1703;
  wire _61573 = _61570 ^ _61572;
  wire _61574 = _7974 ^ _26393;
  wire _61575 = uncoded_block[89] ^ uncoded_block[103];
  wire _61576 = uncoded_block[106] ^ uncoded_block[112];
  wire _61577 = _61575 ^ _61576;
  wire _61578 = _61574 ^ _61577;
  wire _61579 = _61573 ^ _61578;
  wire _61580 = _3253 ^ _59257;
  wire _61581 = uncoded_block[129] ^ uncoded_block[136];
  wire _61582 = _61581 ^ _4043;
  wire _61583 = _61580 ^ _61582;
  wire _61584 = uncoded_block[154] ^ uncoded_block[171];
  wire _61585 = _61584 ^ _9738;
  wire _61586 = uncoded_block[188] ^ uncoded_block[199];
  wire _61587 = _11395 ^ _61586;
  wire _61588 = _61585 ^ _61587;
  wire _61589 = _61583 ^ _61588;
  wire _61590 = _61579 ^ _61589;
  wire _61591 = uncoded_block[201] ^ uncoded_block[206];
  wire _61592 = uncoded_block[218] ^ uncoded_block[236];
  wire _61593 = _61591 ^ _61592;
  wire _61594 = _2552 ^ _4085;
  wire _61595 = _61593 ^ _61594;
  wire _61596 = uncoded_block[246] ^ uncoded_block[268];
  wire _61597 = _61596 ^ _128;
  wire _61598 = uncoded_block[275] ^ uncoded_block[285];
  wire _61599 = _61598 ^ _61427;
  wire _61600 = _61597 ^ _61599;
  wire _61601 = _61595 ^ _61600;
  wire _61602 = uncoded_block[304] ^ uncoded_block[325];
  wire _61603 = _61602 ^ _4838;
  wire _61604 = uncoded_block[348] ^ uncoded_block[367];
  wire _61605 = _61604 ^ _4140;
  wire _61606 = _61603 ^ _61605;
  wire _61607 = _4858 ^ _12541;
  wire _61608 = _10340 ^ _13646;
  wire _61609 = _61607 ^ _61608;
  wire _61610 = _61606 ^ _61609;
  wire _61611 = _61601 ^ _61610;
  wire _61612 = _61590 ^ _61611;
  wire _61613 = uncoded_block[408] ^ uncoded_block[416];
  wire _61614 = _61613 ^ _24711;
  wire _61615 = uncoded_block[453] ^ uncoded_block[462];
  wire _61616 = _4882 ^ _61615;
  wire _61617 = _61614 ^ _61616;
  wire _61618 = uncoded_block[473] ^ uncoded_block[477];
  wire _61619 = _61618 ^ _16693;
  wire _61620 = uncoded_block[484] ^ uncoded_block[492];
  wire _61621 = uncoded_block[498] ^ uncoded_block[507];
  wire _61622 = _61620 ^ _61621;
  wire _61623 = _61619 ^ _61622;
  wire _61624 = _61617 ^ _61623;
  wire _61625 = uncoded_block[520] ^ uncoded_block[530];
  wire _61626 = _20594 ^ _61625;
  wire _61627 = _5628 ^ _4933;
  wire _61628 = _61626 ^ _61627;
  wire _61629 = uncoded_block[552] ^ uncoded_block[578];
  wire _61630 = _61629 ^ _14214;
  wire _61631 = _37253 ^ _9870;
  wire _61632 = _61630 ^ _61631;
  wire _61633 = _61628 ^ _61632;
  wire _61634 = _61624 ^ _61633;
  wire _61635 = uncoded_block[613] ^ uncoded_block[619];
  wire _61636 = _61635 ^ _43761;
  wire _61637 = uncoded_block[649] ^ uncoded_block[654];
  wire _61638 = _2727 ^ _61637;
  wire _61639 = _61636 ^ _61638;
  wire _61640 = _16747 ^ _51249;
  wire _61641 = uncoded_block[673] ^ uncoded_block[684];
  wire _61642 = uncoded_block[687] ^ uncoded_block[695];
  wire _61643 = _61641 ^ _61642;
  wire _61644 = _61640 ^ _61643;
  wire _61645 = _61639 ^ _61644;
  wire _61646 = uncoded_block[706] ^ uncoded_block[717];
  wire _61647 = _11562 ^ _61646;
  wire _61648 = uncoded_block[721] ^ uncoded_block[728];
  wire _61649 = _61648 ^ _26137;
  wire _61650 = _61647 ^ _61649;
  wire _61651 = uncoded_block[756] ^ uncoded_block[761];
  wire _61652 = _24331 ^ _61651;
  wire _61653 = _5020 ^ _31963;
  wire _61654 = _61652 ^ _61653;
  wire _61655 = _61650 ^ _61654;
  wire _61656 = _61645 ^ _61655;
  wire _61657 = _61634 ^ _61656;
  wire _61658 = _61612 ^ _61657;
  wire _61659 = _23442 ^ _18288;
  wire _61660 = _61659 ^ _32803;
  wire _61661 = uncoded_block[837] ^ uncoded_block[850];
  wire _61662 = uncoded_block[853] ^ uncoded_block[867];
  wire _61663 = _61661 ^ _61662;
  wire _61664 = uncoded_block[870] ^ uncoded_block[886];
  wire _61665 = _61664 ^ _28962;
  wire _61666 = _61663 ^ _61665;
  wire _61667 = _61660 ^ _61666;
  wire _61668 = uncoded_block[896] ^ uncoded_block[906];
  wire _61669 = uncoded_block[912] ^ uncoded_block[924];
  wire _61670 = _61668 ^ _61669;
  wire _61671 = uncoded_block[932] ^ uncoded_block[948];
  wire _61672 = uncoded_block[953] ^ uncoded_block[959];
  wire _61673 = _61671 ^ _61672;
  wire _61674 = _61670 ^ _61673;
  wire _61675 = uncoded_block[960] ^ uncoded_block[966];
  wire _61676 = uncoded_block[967] ^ uncoded_block[971];
  wire _61677 = _61675 ^ _61676;
  wire _61678 = uncoded_block[972] ^ uncoded_block[981];
  wire _61679 = uncoded_block[997] ^ uncoded_block[1007];
  wire _61680 = _61678 ^ _61679;
  wire _61681 = _61677 ^ _61680;
  wire _61682 = _61674 ^ _61681;
  wire _61683 = _61667 ^ _61682;
  wire _61684 = uncoded_block[1014] ^ uncoded_block[1023];
  wire _61685 = _61684 ^ _60852;
  wire _61686 = _19777 ^ _12762;
  wire _61687 = _61685 ^ _61686;
  wire _61688 = _1363 ^ _28260;
  wire _61689 = uncoded_block[1086] ^ uncoded_block[1093];
  wire _61690 = _29859 ^ _61689;
  wire _61691 = _61688 ^ _61690;
  wire _61692 = _61687 ^ _61691;
  wire _61693 = _14366 ^ _3713;
  wire _61694 = uncoded_block[1118] ^ uncoded_block[1126];
  wire _61695 = uncoded_block[1129] ^ uncoded_block[1145];
  wire _61696 = _61694 ^ _61695;
  wire _61697 = _61693 ^ _61696;
  wire _61698 = uncoded_block[1173] ^ uncoded_block[1179];
  wire _61699 = _9502 ^ _61698;
  wire _61700 = _4482 ^ _12808;
  wire _61701 = _61699 ^ _61700;
  wire _61702 = _61697 ^ _61701;
  wire _61703 = _61692 ^ _61702;
  wire _61704 = _61683 ^ _61703;
  wire _61705 = uncoded_block[1190] ^ uncoded_block[1207];
  wire _61706 = uncoded_block[1208] ^ uncoded_block[1219];
  wire _61707 = _61705 ^ _61706;
  wire _61708 = _2223 ^ _22188;
  wire _61709 = _61707 ^ _61708;
  wire _61710 = uncoded_block[1239] ^ uncoded_block[1255];
  wire _61711 = uncoded_block[1257] ^ uncoded_block[1262];
  wire _61712 = _61710 ^ _61711;
  wire _61713 = uncoded_block[1264] ^ uncoded_block[1272];
  wire _61714 = _61713 ^ _639;
  wire _61715 = _61712 ^ _61714;
  wire _61716 = _61709 ^ _61715;
  wire _61717 = _9545 ^ _39382;
  wire _61718 = _654 ^ _40932;
  wire _61719 = _61717 ^ _61718;
  wire _61720 = uncoded_block[1341] ^ uncoded_block[1351];
  wire _61721 = _61720 ^ _11773;
  wire _61722 = _61360 ^ _23589;
  wire _61723 = _61721 ^ _61722;
  wire _61724 = _61719 ^ _61723;
  wire _61725 = _61716 ^ _61724;
  wire _61726 = uncoded_block[1386] ^ uncoded_block[1398];
  wire _61727 = _61726 ^ _2297;
  wire _61728 = uncoded_block[1421] ^ uncoded_block[1428];
  wire _61729 = _23163 ^ _61728;
  wire _61730 = _61727 ^ _61729;
  wire _61731 = uncoded_block[1451] ^ uncoded_block[1460];
  wire _61732 = _24065 ^ _61731;
  wire _61733 = uncoded_block[1475] ^ uncoded_block[1491];
  wire _61734 = _18919 ^ _61733;
  wire _61735 = _61732 ^ _61734;
  wire _61736 = _61730 ^ _61735;
  wire _61737 = uncoded_block[1499] ^ uncoded_block[1513];
  wire _61738 = uncoded_block[1521] ^ uncoded_block[1546];
  wire _61739 = _61737 ^ _61738;
  wire _61740 = _6015 ^ _32985;
  wire _61741 = _61739 ^ _61740;
  wire _61742 = _9080 ^ _15537;
  wire _61743 = _8496 ^ _11849;
  wire _61744 = _61742 ^ _61743;
  wire _61745 = _61741 ^ _61744;
  wire _61746 = _61736 ^ _61745;
  wire _61747 = _61725 ^ _61746;
  wire _61748 = _61704 ^ _61747;
  wire _61749 = _61658 ^ _61748;
  wire _61750 = uncoded_block[1609] ^ uncoded_block[1616];
  wire _61751 = _61750 ^ _9095;
  wire _61752 = uncoded_block[1631] ^ uncoded_block[1643];
  wire _61753 = _61752 ^ _4678;
  wire _61754 = _61751 ^ _61753;
  wire _61755 = _46508 ^ _830;
  wire _61756 = _4698 ^ _54216;
  wire _61757 = _61755 ^ _61756;
  wire _61758 = _61754 ^ _61757;
  wire _61759 = _61758 ^ uncoded_block[1721];
  wire _61760 = _61749 ^ _61759;
  wire _61761 = _4712 ^ _22326;
  wire _61762 = uncoded_block[25] ^ uncoded_block[35];
  wire _61763 = _44790 ^ _61762;
  wire _61764 = _61761 ^ _61763;
  wire _61765 = uncoded_block[57] ^ uncoded_block[66];
  wire _61766 = _12429 ^ _61765;
  wire _61767 = _24155 ^ _61766;
  wire _61768 = _61764 ^ _61767;
  wire _61769 = uncoded_block[76] ^ uncoded_block[83];
  wire _61770 = _61769 ^ _4738;
  wire _61771 = uncoded_block[91] ^ uncoded_block[102];
  wire _61772 = _61771 ^ _50;
  wire _61773 = _61770 ^ _61772;
  wire _61774 = uncoded_block[136] ^ uncoded_block[144];
  wire _61775 = uncoded_block[146] ^ uncoded_block[153];
  wire _61776 = _61774 ^ _61775;
  wire _61777 = _54597 ^ _61776;
  wire _61778 = _61773 ^ _61777;
  wire _61779 = _61768 ^ _61778;
  wire _61780 = _39128 ^ _60941;
  wire _61781 = uncoded_block[174] ^ uncoded_block[184];
  wire _61782 = _61781 ^ _14616;
  wire _61783 = _61780 ^ _61782;
  wire _61784 = uncoded_block[203] ^ uncoded_block[210];
  wire _61785 = _2532 ^ _61784;
  wire _61786 = _56429 ^ _963;
  wire _61787 = _61785 ^ _61786;
  wire _61788 = _61783 ^ _61787;
  wire _61789 = _29642 ^ _20021;
  wire _61790 = _15656 ^ _4095;
  wire _61791 = _61789 ^ _61790;
  wire _61792 = uncoded_block[277] ^ uncoded_block[285];
  wire _61793 = _61792 ^ _15665;
  wire _61794 = uncoded_block[297] ^ uncoded_block[306];
  wire _61795 = _61794 ^ _4830;
  wire _61796 = _61793 ^ _61795;
  wire _61797 = _61791 ^ _61796;
  wire _61798 = _61788 ^ _61797;
  wire _61799 = _61779 ^ _61798;
  wire _61800 = _13625 ^ _30117;
  wire _61801 = uncoded_block[353] ^ uncoded_block[363];
  wire _61802 = _13629 ^ _61801;
  wire _61803 = _61800 ^ _61802;
  wire _61804 = _18160 ^ _173;
  wire _61805 = uncoded_block[381] ^ uncoded_block[396];
  wire _61806 = _20056 ^ _61805;
  wire _61807 = _61804 ^ _61806;
  wire _61808 = _61803 ^ _61807;
  wire _61809 = _2625 ^ _12545;
  wire _61810 = _40748 ^ _6894;
  wire _61811 = _61809 ^ _61810;
  wire _61812 = uncoded_block[431] ^ uncoded_block[439];
  wire _61813 = _61812 ^ _42300;
  wire _61814 = _56716 ^ _31024;
  wire _61815 = _61813 ^ _61814;
  wire _61816 = _61811 ^ _61815;
  wire _61817 = _61808 ^ _61816;
  wire _61818 = uncoded_block[504] ^ uncoded_block[511];
  wire _61819 = _61442 ^ _61818;
  wire _61820 = _8122 ^ _4922;
  wire _61821 = _61819 ^ _61820;
  wire _61822 = _3450 ^ _1115;
  wire _61823 = uncoded_block[565] ^ uncoded_block[577];
  wire _61824 = _9314 ^ _61823;
  wire _61825 = _61822 ^ _61824;
  wire _61826 = _61821 ^ _61825;
  wire _61827 = uncoded_block[583] ^ uncoded_block[591];
  wire _61828 = _61827 ^ _21565;
  wire _61829 = uncoded_block[612] ^ uncoded_block[624];
  wire _61830 = _41941 ^ _61829;
  wire _61831 = _61828 ^ _61830;
  wire _61832 = _8159 ^ _6331;
  wire _61833 = _26545 ^ _2729;
  wire _61834 = _61832 ^ _61833;
  wire _61835 = _61831 ^ _61834;
  wire _61836 = _61826 ^ _61835;
  wire _61837 = _61817 ^ _61836;
  wire _61838 = _61799 ^ _61837;
  wire _61839 = uncoded_block[650] ^ uncoded_block[666];
  wire _61840 = uncoded_block[671] ^ uncoded_block[684];
  wire _61841 = _61839 ^ _61840;
  wire _61842 = _3527 ^ _11557;
  wire _61843 = _61841 ^ _61842;
  wire _61844 = _7595 ^ _17266;
  wire _61845 = _30221 ^ _1988;
  wire _61846 = _61844 ^ _61845;
  wire _61847 = _61843 ^ _61846;
  wire _61848 = uncoded_block[741] ^ uncoded_block[753];
  wire _61849 = _1206 ^ _61848;
  wire _61850 = uncoded_block[767] ^ uncoded_block[774];
  wire _61851 = _359 ^ _61850;
  wire _61852 = _61849 ^ _61851;
  wire _61853 = uncoded_block[779] ^ uncoded_block[785];
  wire _61854 = _61853 ^ _31963;
  wire _61855 = _3574 ^ _26588;
  wire _61856 = _61854 ^ _61855;
  wire _61857 = _61852 ^ _61856;
  wire _61858 = _61847 ^ _61857;
  wire _61859 = uncoded_block[809] ^ uncoded_block[816];
  wire _61860 = uncoded_block[817] ^ uncoded_block[825];
  wire _61861 = _61859 ^ _61860;
  wire _61862 = uncoded_block[828] ^ uncoded_block[834];
  wire _61863 = _61862 ^ _401;
  wire _61864 = _61861 ^ _61863;
  wire _61865 = _11610 ^ _3600;
  wire _61866 = uncoded_block[866] ^ uncoded_block[872];
  wire _61867 = _23010 ^ _61866;
  wire _61868 = _61865 ^ _61867;
  wire _61869 = _61864 ^ _61868;
  wire _61870 = uncoded_block[880] ^ uncoded_block[886];
  wire _61871 = _61870 ^ _2061;
  wire _61872 = _13251 ^ _5761;
  wire _61873 = _61871 ^ _61872;
  wire _61874 = uncoded_block[915] ^ uncoded_block[924];
  wire _61875 = uncoded_block[925] ^ uncoded_block[933];
  wire _61876 = _61874 ^ _61875;
  wire _61877 = uncoded_block[937] ^ uncoded_block[944];
  wire _61878 = _61877 ^ _14329;
  wire _61879 = _61876 ^ _61878;
  wire _61880 = _61873 ^ _61879;
  wire _61881 = _61869 ^ _61880;
  wire _61882 = _61858 ^ _61881;
  wire _61883 = uncoded_block[968] ^ uncoded_block[977];
  wire _61884 = _61883 ^ _2100;
  wire _61885 = _4397 ^ _6457;
  wire _61886 = _61884 ^ _61885;
  wire _61887 = uncoded_block[1003] ^ uncoded_block[1016];
  wire _61888 = _61887 ^ _48635;
  wire _61889 = uncoded_block[1035] ^ uncoded_block[1043];
  wire _61890 = _39719 ^ _61889;
  wire _61891 = _61888 ^ _61890;
  wire _61892 = _61886 ^ _61891;
  wire _61893 = uncoded_block[1046] ^ uncoded_block[1054];
  wire _61894 = _61893 ^ _11122;
  wire _61895 = _15396 ^ _42736;
  wire _61896 = _61894 ^ _61895;
  wire _61897 = _30740 ^ _1378;
  wire _61898 = _549 ^ _8339;
  wire _61899 = _61897 ^ _61898;
  wire _61900 = _61896 ^ _61899;
  wire _61901 = _61892 ^ _61900;
  wire _61902 = uncoded_block[1122] ^ uncoded_block[1134];
  wire _61903 = _61902 ^ _9496;
  wire _61904 = _15420 ^ _3727;
  wire _61905 = _61903 ^ _61904;
  wire _61906 = _7749 ^ _2965;
  wire _61907 = uncoded_block[1190] ^ uncoded_block[1195];
  wire _61908 = uncoded_block[1197] ^ uncoded_block[1210];
  wire _61909 = _61907 ^ _61908;
  wire _61910 = _61906 ^ _61909;
  wire _61911 = _61905 ^ _61910;
  wire _61912 = _3762 ^ _49397;
  wire _61913 = uncoded_block[1221] ^ uncoded_block[1236];
  wire _61914 = _61913 ^ _5221;
  wire _61915 = _61912 ^ _61914;
  wire _61916 = _3784 ^ _2244;
  wire _61917 = _30789 ^ _23124;
  wire _61918 = _61916 ^ _61917;
  wire _61919 = _61915 ^ _61918;
  wire _61920 = _61911 ^ _61919;
  wire _61921 = _61901 ^ _61920;
  wire _61922 = _61882 ^ _61921;
  wire _61923 = _61838 ^ _61922;
  wire _61924 = _9545 ^ _6563;
  wire _61925 = uncoded_block[1298] ^ uncoded_block[1309];
  wire _61926 = uncoded_block[1319] ^ uncoded_block[1338];
  wire _61927 = _61925 ^ _61926;
  wire _61928 = _61924 ^ _61927;
  wire _61929 = _5262 ^ _32102;
  wire _61930 = uncoded_block[1355] ^ uncoded_block[1368];
  wire _61931 = _33363 ^ _61930;
  wire _61932 = _61929 ^ _61931;
  wire _61933 = _61928 ^ _61932;
  wire _61934 = _684 ^ _10108;
  wire _61935 = uncoded_block[1400] ^ uncoded_block[1408];
  wire _61936 = _38613 ^ _61935;
  wire _61937 = _61934 ^ _61936;
  wire _61938 = uncoded_block[1413] ^ uncoded_block[1424];
  wire _61939 = _61938 ^ _1531;
  wire _61940 = uncoded_block[1453] ^ uncoded_block[1458];
  wire _61941 = _35416 ^ _61940;
  wire _61942 = _61939 ^ _61941;
  wire _61943 = _61937 ^ _61942;
  wire _61944 = _61933 ^ _61943;
  wire _61945 = uncoded_block[1464] ^ uncoded_block[1471];
  wire _61946 = uncoded_block[1477] ^ uncoded_block[1485];
  wire _61947 = _61945 ^ _61946;
  wire _61948 = uncoded_block[1489] ^ uncoded_block[1494];
  wire _61949 = uncoded_block[1499] ^ uncoded_block[1504];
  wire _61950 = _61948 ^ _61949;
  wire _61951 = _61947 ^ _61950;
  wire _61952 = _3894 ^ _58945;
  wire _61953 = uncoded_block[1522] ^ uncoded_block[1529];
  wire _61954 = uncoded_block[1534] ^ uncoded_block[1547];
  wire _61955 = _61953 ^ _61954;
  wire _61956 = _61952 ^ _61955;
  wire _61957 = _61951 ^ _61956;
  wire _61958 = _3914 ^ _23640;
  wire _61959 = uncoded_block[1572] ^ uncoded_block[1578];
  wire _61960 = _1606 ^ _61959;
  wire _61961 = _61958 ^ _61960;
  wire _61962 = _20397 ^ _56938;
  wire _61963 = uncoded_block[1599] ^ uncoded_block[1611];
  wire _61964 = _3933 ^ _61963;
  wire _61965 = _61962 ^ _61964;
  wire _61966 = _61961 ^ _61965;
  wire _61967 = _61957 ^ _61966;
  wire _61968 = _61944 ^ _61967;
  wire _61969 = uncoded_block[1612] ^ uncoded_block[1617];
  wire _61970 = uncoded_block[1618] ^ uncoded_block[1625];
  wire _61971 = _61969 ^ _61970;
  wire _61972 = uncoded_block[1638] ^ uncoded_block[1645];
  wire _61973 = _3942 ^ _61972;
  wire _61974 = _61971 ^ _61973;
  wire _61975 = uncoded_block[1652] ^ uncoded_block[1662];
  wire _61976 = _14530 ^ _61975;
  wire _61977 = uncoded_block[1666] ^ uncoded_block[1676];
  wire _61978 = uncoded_block[1678] ^ uncoded_block[1687];
  wire _61979 = _61977 ^ _61978;
  wire _61980 = _61976 ^ _61979;
  wire _61981 = _61974 ^ _61980;
  wire _61982 = _12400 ^ _847;
  wire _61983 = _61982 ^ uncoded_block[1716];
  wire _61984 = _61981 ^ _61983;
  wire _61985 = _61968 ^ _61984;
  wire _61986 = _61923 ^ _61985;
  wire _61987 = uncoded_block[11] ^ uncoded_block[19];
  wire _61988 = uncoded_block[23] ^ uncoded_block[32];
  wire _61989 = _61987 ^ _61988;
  wire _61990 = _25948 ^ _2474;
  wire _61991 = _61989 ^ _61990;
  wire _61992 = uncoded_block[108] ^ uncoded_block[129];
  wire _61993 = _910 ^ _61992;
  wire _61994 = _9730 ^ _2511;
  wire _61995 = _61993 ^ _61994;
  wire _61996 = _61991 ^ _61995;
  wire _61997 = uncoded_block[159] ^ uncoded_block[178];
  wire _61998 = _61997 ^ _1763;
  wire _61999 = uncoded_block[198] ^ uncoded_block[215];
  wire _62000 = uncoded_block[220] ^ uncoded_block[244];
  wire _62001 = _61999 ^ _62000;
  wire _62002 = _61998 ^ _62001;
  wire _62003 = uncoded_block[258] ^ uncoded_block[289];
  wire _62004 = _62003 ^ _1807;
  wire _62005 = uncoded_block[322] ^ uncoded_block[335];
  wire _62006 = _12516 ^ _62005;
  wire _62007 = _62004 ^ _62006;
  wire _62008 = _62002 ^ _62007;
  wire _62009 = _61996 ^ _62008;
  wire _62010 = uncoded_block[341] ^ uncoded_block[348];
  wire _62011 = _62010 ^ _3369;
  wire _62012 = uncoded_block[375] ^ uncoded_block[391];
  wire _62013 = _62012 ^ _48868;
  wire _62014 = _62011 ^ _62013;
  wire _62015 = uncoded_block[419] ^ uncoded_block[429];
  wire _62016 = _62015 ^ _31459;
  wire _62017 = _19621 ^ _7504;
  wire _62018 = _62016 ^ _62017;
  wire _62019 = _62014 ^ _62018;
  wire _62020 = uncoded_block[464] ^ uncoded_block[486];
  wire _62021 = uncoded_block[506] ^ uncoded_block[514];
  wire _62022 = _62020 ^ _62021;
  wire _62023 = uncoded_block[515] ^ uncoded_block[534];
  wire _62024 = uncoded_block[555] ^ uncoded_block[564];
  wire _62025 = _62023 ^ _62024;
  wire _62026 = _62022 ^ _62025;
  wire _62027 = uncoded_block[579] ^ uncoded_block[591];
  wire _62028 = uncoded_block[593] ^ uncoded_block[610];
  wire _62029 = _62027 ^ _62028;
  wire _62030 = uncoded_block[626] ^ uncoded_block[634];
  wire _62031 = _13178 ^ _62030;
  wire _62032 = _62029 ^ _62031;
  wire _62033 = _62026 ^ _62032;
  wire _62034 = _62019 ^ _62033;
  wire _62035 = _62009 ^ _62034;
  wire _62036 = uncoded_block[661] ^ uncoded_block[674];
  wire _62037 = _16241 ^ _62036;
  wire _62038 = uncoded_block[691] ^ uncoded_block[703];
  wire _62039 = _62038 ^ _11004;
  wire _62040 = _62037 ^ _62039;
  wire _62041 = uncoded_block[724] ^ uncoded_block[735];
  wire _62042 = _9369 ^ _62041;
  wire _62043 = uncoded_block[746] ^ uncoded_block[762];
  wire _62044 = _62043 ^ _2783;
  wire _62045 = _62042 ^ _62044;
  wire _62046 = _62040 ^ _62045;
  wire _62047 = uncoded_block[784] ^ uncoded_block[795];
  wire _62048 = _62047 ^ _8793;
  wire _62049 = uncoded_block[807] ^ uncoded_block[817];
  wire _62050 = uncoded_block[841] ^ uncoded_block[852];
  wire _62051 = _62049 ^ _62050;
  wire _62052 = _62048 ^ _62051;
  wire _62053 = uncoded_block[858] ^ uncoded_block[874];
  wire _62054 = uncoded_block[884] ^ uncoded_block[893];
  wire _62055 = _62053 ^ _62054;
  wire _62056 = uncoded_block[903] ^ uncoded_block[920];
  wire _62057 = _1278 ^ _62056;
  wire _62058 = _62055 ^ _62057;
  wire _62059 = _62052 ^ _62058;
  wire _62060 = _62046 ^ _62059;
  wire _62061 = uncoded_block[940] ^ uncoded_block[957];
  wire _62062 = uncoded_block[973] ^ uncoded_block[981];
  wire _62063 = _62061 ^ _62062;
  wire _62064 = uncoded_block[986] ^ uncoded_block[1002];
  wire _62065 = _62064 ^ _2118;
  wire _62066 = _62063 ^ _62065;
  wire _62067 = uncoded_block[1028] ^ uncoded_block[1037];
  wire _62068 = uncoded_block[1041] ^ uncoded_block[1055];
  wire _62069 = _62067 ^ _62068;
  wire _62070 = uncoded_block[1075] ^ uncoded_block[1081];
  wire _62071 = _2922 ^ _62070;
  wire _62072 = _62069 ^ _62071;
  wire _62073 = _62066 ^ _62072;
  wire _62074 = uncoded_block[1087] ^ uncoded_block[1095];
  wire _62075 = _62074 ^ _5176;
  wire _62076 = uncoded_block[1130] ^ uncoded_block[1135];
  wire _62077 = _62076 ^ _1403;
  wire _62078 = _62075 ^ _62077;
  wire _62079 = _59351 ^ _49583;
  wire _62080 = uncoded_block[1209] ^ uncoded_block[1221];
  wire _62081 = uncoded_block[1227] ^ uncoded_block[1244];
  wire _62082 = _62080 ^ _62081;
  wire _62083 = _62079 ^ _62082;
  wire _62084 = _62078 ^ _62083;
  wire _62085 = _62073 ^ _62084;
  wire _62086 = _62060 ^ _62085;
  wire _62087 = _62035 ^ _62086;
  wire _62088 = uncoded_block[1247] ^ uncoded_block[1267];
  wire _62089 = uncoded_block[1274] ^ uncoded_block[1286];
  wire _62090 = _62088 ^ _62089;
  wire _62091 = uncoded_block[1296] ^ uncoded_block[1322];
  wire _62092 = _3801 ^ _62091;
  wire _62093 = _62090 ^ _62092;
  wire _62094 = uncoded_block[1326] ^ uncoded_block[1334];
  wire _62095 = _62094 ^ _4556;
  wire _62096 = _61214 ^ _1519;
  wire _62097 = _62095 ^ _62096;
  wire _62098 = _62093 ^ _62097;
  wire _62099 = uncoded_block[1409] ^ uncoded_block[1426];
  wire _62100 = uncoded_block[1445] ^ uncoded_block[1453];
  wire _62101 = _62099 ^ _62100;
  wire _62102 = uncoded_block[1461] ^ uncoded_block[1472];
  wire _62103 = _62102 ^ _735;
  wire _62104 = _62101 ^ _62103;
  wire _62105 = uncoded_block[1493] ^ uncoded_block[1497];
  wire _62106 = uncoded_block[1501] ^ uncoded_block[1518];
  wire _62107 = _62105 ^ _62106;
  wire _62108 = uncoded_block[1522] ^ uncoded_block[1551];
  wire _62109 = uncoded_block[1557] ^ uncoded_block[1570];
  wire _62110 = _62108 ^ _62109;
  wire _62111 = _62107 ^ _62110;
  wire _62112 = _62104 ^ _62111;
  wire _62113 = _62098 ^ _62112;
  wire _62114 = _13478 ^ _61547;
  wire _62115 = uncoded_block[1595] ^ uncoded_block[1611];
  wire _62116 = _62115 ^ _13494;
  wire _62117 = _62114 ^ _62116;
  wire _62118 = uncoded_block[1631] ^ uncoded_block[1644];
  wire _62119 = uncoded_block[1665] ^ uncoded_block[1677];
  wire _62120 = _62118 ^ _62119;
  wire _62121 = uncoded_block[1680] ^ uncoded_block[1687];
  wire _62122 = _62121 ^ _2435;
  wire _62123 = _62120 ^ _62122;
  wire _62124 = _62117 ^ _62123;
  wire _62125 = _62124 ^ uncoded_block[1722];
  wire _62126 = _62113 ^ _62125;
  wire _62127 = _62087 ^ _62126;
  wire _62128 = _56963 ^ _20937;
  wire _62129 = _58985 ^ _62128;
  wire _62130 = uncoded_block[41] ^ uncoded_block[48];
  wire _62131 = _879 ^ _62130;
  wire _62132 = _27252 ^ _5440;
  wire _62133 = _62131 ^ _62132;
  wire _62134 = _62129 ^ _62133;
  wire _62135 = _11904 ^ _28765;
  wire _62136 = uncoded_block[83] ^ uncoded_block[89];
  wire _62137 = uncoded_block[90] ^ uncoded_block[98];
  wire _62138 = _62136 ^ _62137;
  wire _62139 = _62135 ^ _62138;
  wire _62140 = uncoded_block[109] ^ uncoded_block[119];
  wire _62141 = _910 ^ _62140;
  wire _62142 = _23269 ^ _917;
  wire _62143 = _62141 ^ _62142;
  wire _62144 = _62139 ^ _62143;
  wire _62145 = _62134 ^ _62144;
  wire _62146 = _27274 ^ _30511;
  wire _62147 = uncoded_block[148] ^ uncoded_block[166];
  wire _62148 = _62147 ^ _23729;
  wire _62149 = _62146 ^ _62148;
  wire _62150 = _13032 ^ _1757;
  wire _62151 = _62150 ^ _59012;
  wire _62152 = _62149 ^ _62151;
  wire _62153 = _6158 ^ _11405;
  wire _62154 = _60170 ^ _17617;
  wire _62155 = _62153 ^ _62154;
  wire _62156 = uncoded_block[242] ^ uncoded_block[250];
  wire _62157 = _25104 ^ _62156;
  wire _62158 = _39537 ^ _26441;
  wire _62159 = _62157 ^ _62158;
  wire _62160 = _62155 ^ _62159;
  wire _62161 = _62152 ^ _62160;
  wire _62162 = _62145 ^ _62161;
  wire _62163 = uncoded_block[264] ^ uncoded_block[272];
  wire _62164 = _62163 ^ _3321;
  wire _62165 = _36768 ^ _1803;
  wire _62166 = _62164 ^ _62165;
  wire _62167 = _6837 ^ _13615;
  wire _62168 = _7453 ^ _20539;
  wire _62169 = _62167 ^ _62168;
  wire _62170 = _62166 ^ _62169;
  wire _62171 = uncoded_block[329] ^ uncoded_block[336];
  wire _62172 = _48476 ^ _62171;
  wire _62173 = _32687 ^ _5541;
  wire _62174 = _62172 ^ _62173;
  wire _62175 = uncoded_block[354] ^ uncoded_block[361];
  wire _62176 = _62175 ^ _17658;
  wire _62177 = _4141 ^ _59041;
  wire _62178 = _62176 ^ _62177;
  wire _62179 = _62174 ^ _62178;
  wire _62180 = _62170 ^ _62179;
  wire _62181 = _1847 ^ _10341;
  wire _62182 = _59044 ^ _59046;
  wire _62183 = _62181 ^ _62182;
  wire _62184 = _201 ^ _1067;
  wire _62185 = _9275 ^ _24254;
  wire _62186 = _62184 ^ _62185;
  wire _62187 = _62183 ^ _62186;
  wire _62188 = uncoded_block[502] ^ uncoded_block[517];
  wire _62189 = _21987 ^ _62188;
  wire _62190 = _62189 ^ _59065;
  wire _62191 = _59056 ^ _62190;
  wire _62192 = _62187 ^ _62191;
  wire _62193 = _62180 ^ _62192;
  wire _62194 = _62162 ^ _62193;
  wire _62195 = _55228 ^ _4934;
  wire _62196 = _59067 ^ _62195;
  wire _62197 = _32327 ^ _21087;
  wire _62198 = _4229 ^ _22012;
  wire _62199 = _62197 ^ _62198;
  wire _62200 = _62196 ^ _62199;
  wire _62201 = _34013 ^ _41941;
  wire _62202 = uncoded_block[617] ^ uncoded_block[634];
  wire _62203 = _59076 ^ _62202;
  wire _62204 = _62201 ^ _62203;
  wire _62205 = uncoded_block[640] ^ uncoded_block[648];
  wire _62206 = _5661 ^ _62205;
  wire _62207 = _302 ^ _41957;
  wire _62208 = _62206 ^ _62207;
  wire _62209 = _62204 ^ _62208;
  wire _62210 = _62200 ^ _62209;
  wire _62211 = _9885 ^ _17745;
  wire _62212 = uncoded_block[675] ^ uncoded_block[681];
  wire _62213 = _62212 ^ _15281;
  wire _62214 = _62211 ^ _62213;
  wire _62215 = uncoded_block[688] ^ uncoded_block[692];
  wire _62216 = uncoded_block[693] ^ uncoded_block[701];
  wire _62217 = _62215 ^ _62216;
  wire _62218 = uncoded_block[704] ^ uncoded_block[715];
  wire _62219 = uncoded_block[734] ^ uncoded_block[739];
  wire _62220 = _62218 ^ _62219;
  wire _62221 = _62217 ^ _62220;
  wire _62222 = _62214 ^ _62221;
  wire _62223 = uncoded_block[742] ^ uncoded_block[753];
  wire _62224 = uncoded_block[754] ^ uncoded_block[762];
  wire _62225 = _62223 ^ _62224;
  wire _62226 = _13215 ^ _18274;
  wire _62227 = _62225 ^ _62226;
  wire _62228 = _34059 ^ _3577;
  wire _62229 = _48582 ^ _62228;
  wire _62230 = _62227 ^ _62229;
  wire _62231 = _62222 ^ _62230;
  wire _62232 = _62210 ^ _62231;
  wire _62233 = uncoded_block[806] ^ uncoded_block[814];
  wire _62234 = _62233 ^ _57409;
  wire _62235 = _62234 ^ _57415;
  wire _62236 = _59105 ^ _16811;
  wire _62237 = uncoded_block[897] ^ uncoded_block[910];
  wire _62238 = _59108 ^ _62237;
  wire _62239 = _62236 ^ _62238;
  wire _62240 = _62235 ^ _62239;
  wire _62241 = uncoded_block[929] ^ uncoded_block[936];
  wire _62242 = _31995 ^ _62241;
  wire _62243 = _59115 ^ _62242;
  wire _62244 = _453 ^ _13266;
  wire _62245 = uncoded_block[951] ^ uncoded_block[956];
  wire _62246 = _62245 ^ _45753;
  wire _62247 = _62244 ^ _62246;
  wire _62248 = _62243 ^ _62247;
  wire _62249 = _62240 ^ _62248;
  wire _62250 = _1310 ^ _11648;
  wire _62251 = uncoded_block[983] ^ uncoded_block[993];
  wire _62252 = _13272 ^ _62251;
  wire _62253 = _62250 ^ _62252;
  wire _62254 = _484 ^ _52890;
  wire _62255 = uncoded_block[1019] ^ uncoded_block[1022];
  wire _62256 = _62255 ^ _35710;
  wire _62257 = _62254 ^ _62256;
  wire _62258 = _62253 ^ _62257;
  wire _62259 = _50575 ^ _6475;
  wire _62260 = uncoded_block[1049] ^ uncoded_block[1061];
  wire _62261 = _62260 ^ _8889;
  wire _62262 = _62259 ^ _62261;
  wire _62263 = _5156 ^ _9480;
  wire _62264 = _8906 ^ _1378;
  wire _62265 = _62263 ^ _62264;
  wire _62266 = _62262 ^ _62265;
  wire _62267 = _62258 ^ _62266;
  wire _62268 = _62249 ^ _62267;
  wire _62269 = _62232 ^ _62268;
  wire _62270 = _62194 ^ _62269;
  wire _62271 = _25318 ^ _20761;
  wire _62272 = _14882 ^ _3713;
  wire _62273 = _62271 ^ _62272;
  wire _62274 = _59148 ^ _59153;
  wire _62275 = _62273 ^ _62274;
  wire _62276 = _1407 ^ _10608;
  wire _62277 = _62276 ^ _59158;
  wire _62278 = _59159 ^ _608;
  wire _62279 = _2986 ^ _43141;
  wire _62280 = _62278 ^ _62279;
  wire _62281 = _62277 ^ _62280;
  wire _62282 = _62275 ^ _62281;
  wire _62283 = _10067 ^ _13365;
  wire _62284 = _3780 ^ _56573;
  wire _62285 = _62283 ^ _62284;
  wire _62286 = uncoded_block[1270] ^ uncoded_block[1278];
  wire _62287 = _5235 ^ _62286;
  wire _62288 = _23123 ^ _19365;
  wire _62289 = _62287 ^ _62288;
  wire _62290 = _62285 ^ _62289;
  wire _62291 = uncoded_block[1301] ^ uncoded_block[1310];
  wire _62292 = uncoded_block[1313] ^ uncoded_block[1327];
  wire _62293 = _62291 ^ _62292;
  wire _62294 = _56878 ^ _62293;
  wire _62295 = _59179 ^ _11771;
  wire _62296 = _10097 ^ _13407;
  wire _62297 = _62295 ^ _62296;
  wire _62298 = _62294 ^ _62297;
  wire _62299 = _62290 ^ _62298;
  wire _62300 = _62282 ^ _62299;
  wire _62301 = _7219 ^ _19864;
  wire _62302 = _59188 ^ _62301;
  wire _62303 = _4572 ^ _40588;
  wire _62304 = _3069 ^ _6607;
  wire _62305 = _62303 ^ _62304;
  wire _62306 = _62302 ^ _62305;
  wire _62307 = _31274 ^ _21323;
  wire _62308 = _15982 ^ _45085;
  wire _62309 = _62307 ^ _62308;
  wire _62310 = _59201 ^ _36213;
  wire _62311 = uncoded_block[1469] ^ uncoded_block[1475];
  wire _62312 = _9602 ^ _62311;
  wire _62313 = _62310 ^ _62312;
  wire _62314 = _62309 ^ _62313;
  wire _62315 = _62306 ^ _62314;
  wire _62316 = uncoded_block[1480] ^ uncoded_block[1490];
  wire _62317 = _9610 ^ _62316;
  wire _62318 = _11260 ^ _9618;
  wire _62319 = _62317 ^ _62318;
  wire _62320 = _2356 ^ _12352;
  wire _62321 = _11272 ^ _39050;
  wire _62322 = _62320 ^ _62321;
  wire _62323 = _62319 ^ _62322;
  wire _62324 = _1587 ^ _57216;
  wire _62325 = uncoded_block[1562] ^ uncoded_block[1580];
  wire _62326 = _3914 ^ _62325;
  wire _62327 = _62324 ^ _62326;
  wire _62328 = _16515 ^ _11292;
  wire _62329 = _14517 ^ _42166;
  wire _62330 = _62328 ^ _62329;
  wire _62331 = _62327 ^ _62330;
  wire _62332 = _62323 ^ _62331;
  wire _62333 = _62315 ^ _62332;
  wire _62334 = _62300 ^ _62333;
  wire _62335 = _29997 ^ _6046;
  wire _62336 = _18511 ^ _16529;
  wire _62337 = _62335 ^ _62336;
  wire _62338 = _12383 ^ _3953;
  wire _62339 = _820 ^ _25476;
  wire _62340 = _62338 ^ _62339;
  wire _62341 = _62337 ^ _62340;
  wire _62342 = uncoded_block[1672] ^ uncoded_block[1679];
  wire _62343 = _62342 ^ _11327;
  wire _62344 = uncoded_block[1708] ^ uncoded_block[1718];
  wire _62345 = _3976 ^ _62344;
  wire _62346 = _62343 ^ _62345;
  wire _62347 = _62346 ^ uncoded_block[1722];
  wire _62348 = _62341 ^ _62347;
  wire _62349 = _62334 ^ _62348;
  wire _62350 = _62270 ^ _62349;
  wire _62351 = uncoded_block[6] ^ uncoded_block[14];
  wire _62352 = uncoded_block[67] ^ uncoded_block[82];
  wire _62353 = _62351 ^ _62352;
  wire _62354 = uncoded_block[86] ^ uncoded_block[105];
  wire _62355 = uncoded_block[122] ^ uncoded_block[128];
  wire _62356 = _62354 ^ _62355;
  wire _62357 = _62353 ^ _62356;
  wire _62358 = uncoded_block[133] ^ uncoded_block[153];
  wire _62359 = _62358 ^ _3281;
  wire _62360 = uncoded_block[230] ^ uncoded_block[250];
  wire _62361 = _59688 ^ _62360;
  wire _62362 = _62359 ^ _62361;
  wire _62363 = _62357 ^ _62362;
  wire _62364 = uncoded_block[252] ^ uncoded_block[267];
  wire _62365 = uncoded_block[287] ^ uncoded_block[298];
  wire _62366 = _62364 ^ _62365;
  wire _62367 = uncoded_block[317] ^ uncoded_block[321];
  wire _62368 = uncoded_block[346] ^ uncoded_block[371];
  wire _62369 = _62367 ^ _62368;
  wire _62370 = _62366 ^ _62369;
  wire _62371 = _50446 ^ _26042;
  wire _62372 = _4874 ^ _4890;
  wire _62373 = _62371 ^ _62372;
  wire _62374 = _62370 ^ _62373;
  wire _62375 = _62363 ^ _62374;
  wire _62376 = uncoded_block[487] ^ uncoded_block[498];
  wire _62377 = uncoded_block[506] ^ uncoded_block[527];
  wire _62378 = _62376 ^ _62377;
  wire _62379 = uncoded_block[589] ^ uncoded_block[599];
  wire _62380 = _4925 ^ _62379;
  wire _62381 = _62378 ^ _62380;
  wire _62382 = uncoded_block[605] ^ uncoded_block[612];
  wire _62383 = uncoded_block[628] ^ uncoded_block[640];
  wire _62384 = _62382 ^ _62383;
  wire _62385 = uncoded_block[678] ^ uncoded_block[693];
  wire _62386 = _8755 ^ _62385;
  wire _62387 = _62384 ^ _62386;
  wire _62388 = _62381 ^ _62387;
  wire _62389 = uncoded_block[703] ^ uncoded_block[750];
  wire _62390 = _62389 ^ _14270;
  wire _62391 = uncoded_block[774] ^ uncoded_block[787];
  wire _62392 = _62391 ^ _8228;
  wire _62393 = _62390 ^ _62392;
  wire _62394 = uncoded_block[825] ^ uncoded_block[832];
  wire _62395 = uncoded_block[842] ^ uncoded_block[866];
  wire _62396 = _62394 ^ _62395;
  wire _62397 = uncoded_block[882] ^ uncoded_block[917];
  wire _62398 = uncoded_block[935] ^ uncoded_block[939];
  wire _62399 = _62397 ^ _62398;
  wire _62400 = _62396 ^ _62399;
  wire _62401 = _62393 ^ _62400;
  wire _62402 = _62388 ^ _62401;
  wire _62403 = _62375 ^ _62402;
  wire _62404 = uncoded_block[970] ^ uncoded_block[979];
  wire _62405 = _1300 ^ _62404;
  wire _62406 = uncoded_block[997] ^ uncoded_block[1013];
  wire _62407 = _62406 ^ _61889;
  wire _62408 = _62405 ^ _62407;
  wire _62409 = uncoded_block[1080] ^ uncoded_block[1088];
  wire _62410 = _34122 ^ _62409;
  wire _62411 = _13327 ^ _8933;
  wire _62412 = _62410 ^ _62411;
  wire _62413 = _62408 ^ _62412;
  wire _62414 = uncoded_block[1185] ^ uncoded_block[1191];
  wire _62415 = _62414 ^ _57969;
  wire _62416 = uncoded_block[1220] ^ uncoded_block[1236];
  wire _62417 = uncoded_block[1251] ^ uncoded_block[1267];
  wire _62418 = _62416 ^ _62417;
  wire _62419 = _62415 ^ _62418;
  wire _62420 = uncoded_block[1274] ^ uncoded_block[1283];
  wire _62421 = uncoded_block[1303] ^ uncoded_block[1312];
  wire _62422 = _62420 ^ _62421;
  wire _62423 = uncoded_block[1315] ^ uncoded_block[1337];
  wire _62424 = uncoded_block[1344] ^ uncoded_block[1376];
  wire _62425 = _62423 ^ _62424;
  wire _62426 = _62422 ^ _62425;
  wire _62427 = _62419 ^ _62426;
  wire _62428 = _62413 ^ _62427;
  wire _62429 = uncoded_block[1384] ^ uncoded_block[1395];
  wire _62430 = uncoded_block[1400] ^ uncoded_block[1432];
  wire _62431 = _62429 ^ _62430;
  wire _62432 = uncoded_block[1444] ^ uncoded_block[1452];
  wire _62433 = uncoded_block[1454] ^ uncoded_block[1470];
  wire _62434 = _62432 ^ _62433;
  wire _62435 = _62431 ^ _62434;
  wire _62436 = uncoded_block[1480] ^ uncoded_block[1489];
  wire _62437 = uncoded_block[1498] ^ uncoded_block[1533];
  wire _62438 = _62436 ^ _62437;
  wire _62439 = uncoded_block[1561] ^ uncoded_block[1576];
  wire _62440 = uncoded_block[1580] ^ uncoded_block[1594];
  wire _62441 = _62439 ^ _62440;
  wire _62442 = _62438 ^ _62441;
  wire _62443 = _62435 ^ _62442;
  wire _62444 = uncoded_block[1611] ^ uncoded_block[1631];
  wire _62445 = uncoded_block[1638] ^ uncoded_block[1651];
  wire _62446 = _62444 ^ _62445;
  wire _62447 = uncoded_block[1671] ^ uncoded_block[1702];
  wire _62448 = _53353 ^ _62447;
  wire _62449 = _62446 ^ _62448;
  wire _62450 = _62449 ^ uncoded_block[1714];
  wire _62451 = _62443 ^ _62450;
  wire _62452 = _62428 ^ _62451;
  wire _62453 = _62403 ^ _62452;
  wire _62454 = uncoded_block[3] ^ uncoded_block[21];
  wire _62455 = _62454 ^ _11343;
  wire _62456 = uncoded_block[28] ^ uncoded_block[38];
  wire _62457 = uncoded_block[48] ^ uncoded_block[63];
  wire _62458 = _62456 ^ _62457;
  wire _62459 = _62455 ^ _62458;
  wire _62460 = uncoded_block[70] ^ uncoded_block[89];
  wire _62461 = uncoded_block[94] ^ uncoded_block[102];
  wire _62462 = _62460 ^ _62461;
  wire _62463 = uncoded_block[116] ^ uncoded_block[134];
  wire _62464 = uncoded_block[144] ^ uncoded_block[152];
  wire _62465 = _62463 ^ _62464;
  wire _62466 = _62462 ^ _62465;
  wire _62467 = _62459 ^ _62466;
  wire _62468 = uncoded_block[169] ^ uncoded_block[181];
  wire _62469 = _62468 ^ _17106;
  wire _62470 = uncoded_block[196] ^ uncoded_block[204];
  wire _62471 = _39921 ^ _62470;
  wire _62472 = _62469 ^ _62471;
  wire _62473 = uncoded_block[235] ^ uncoded_block[254];
  wire _62474 = _41482 ^ _62473;
  wire _62475 = uncoded_block[267] ^ uncoded_block[282];
  wire _62476 = _62475 ^ _35159;
  wire _62477 = _62474 ^ _62476;
  wire _62478 = _62472 ^ _62477;
  wire _62479 = _62467 ^ _62478;
  wire _62480 = _9779 ^ _19583;
  wire _62481 = uncoded_block[352] ^ uncoded_block[377];
  wire _62482 = uncoded_block[380] ^ uncoded_block[387];
  wire _62483 = _62481 ^ _62482;
  wire _62484 = _62480 ^ _62483;
  wire _62485 = uncoded_block[389] ^ uncoded_block[401];
  wire _62486 = _62485 ^ _4163;
  wire _62487 = uncoded_block[431] ^ uncoded_block[436];
  wire _62488 = uncoded_block[437] ^ uncoded_block[443];
  wire _62489 = _62487 ^ _62488;
  wire _62490 = _62486 ^ _62489;
  wire _62491 = _62484 ^ _62490;
  wire _62492 = uncoded_block[448] ^ uncoded_block[460];
  wire _62493 = _62492 ^ _5590;
  wire _62494 = uncoded_block[482] ^ uncoded_block[488];
  wire _62495 = uncoded_block[503] ^ uncoded_block[513];
  wire _62496 = _62494 ^ _62495;
  wire _62497 = _62493 ^ _62496;
  wire _62498 = uncoded_block[528] ^ uncoded_block[543];
  wire _62499 = _28503 ^ _62498;
  wire _62500 = uncoded_block[547] ^ uncoded_block[556];
  wire _62501 = _62500 ^ _19153;
  wire _62502 = _62499 ^ _62501;
  wire _62503 = _62497 ^ _62502;
  wire _62504 = _62491 ^ _62503;
  wire _62505 = _62479 ^ _62504;
  wire _62506 = uncoded_block[572] ^ uncoded_block[598];
  wire _62507 = _62506 ^ _8739;
  wire _62508 = uncoded_block[612] ^ uncoded_block[618];
  wire _62509 = _62508 ^ _20125;
  wire _62510 = _62507 ^ _62509;
  wire _62511 = uncoded_block[647] ^ uncoded_block[678];
  wire _62512 = _40023 ^ _62511;
  wire _62513 = uncoded_block[708] ^ uncoded_block[715];
  wire _62514 = _6360 ^ _62513;
  wire _62515 = _62512 ^ _62514;
  wire _62516 = _62510 ^ _62515;
  wire _62517 = _1195 ^ _34442;
  wire _62518 = uncoded_block[770] ^ uncoded_block[777];
  wire _62519 = _7002 ^ _62518;
  wire _62520 = _62517 ^ _62519;
  wire _62521 = _6388 ^ _5035;
  wire _62522 = _11030 ^ _35666;
  wire _62523 = _62521 ^ _62522;
  wire _62524 = _62520 ^ _62523;
  wire _62525 = _62516 ^ _62524;
  wire _62526 = uncoded_block[868] ^ uncoded_block[874];
  wire _62527 = _9949 ^ _62526;
  wire _62528 = uncoded_block[886] ^ uncoded_block[899];
  wire _62529 = _9954 ^ _62528;
  wire _62530 = _62527 ^ _62529;
  wire _62531 = uncoded_block[904] ^ uncoded_block[932];
  wire _62532 = uncoded_block[949] ^ uncoded_block[960];
  wire _62533 = _62531 ^ _62532;
  wire _62534 = _11649 ^ _3659;
  wire _62535 = _62533 ^ _62534;
  wire _62536 = _62530 ^ _62535;
  wire _62537 = uncoded_block[995] ^ uncoded_block[1029];
  wire _62538 = _62537 ^ _26653;
  wire _62539 = uncoded_block[1042] ^ uncoded_block[1051];
  wire _62540 = _62539 ^ _11116;
  wire _62541 = _62538 ^ _62540;
  wire _62542 = _13849 ^ _23969;
  wire _62543 = uncoded_block[1086] ^ uncoded_block[1098];
  wire _62544 = uncoded_block[1100] ^ uncoded_block[1119];
  wire _62545 = _62543 ^ _62544;
  wire _62546 = _62542 ^ _62545;
  wire _62547 = _62541 ^ _62546;
  wire _62548 = _62536 ^ _62547;
  wire _62549 = _62525 ^ _62548;
  wire _62550 = _62505 ^ _62549;
  wire _62551 = uncoded_block[1141] ^ uncoded_block[1145];
  wire _62552 = _57152 ^ _62551;
  wire _62553 = uncoded_block[1159] ^ uncoded_block[1171];
  wire _62554 = _62553 ^ _2967;
  wire _62555 = _62552 ^ _62554;
  wire _62556 = uncoded_block[1176] ^ uncoded_block[1189];
  wire _62557 = _62556 ^ _61907;
  wire _62558 = uncoded_block[1236] ^ uncoded_block[1249];
  wire _62559 = _8958 ^ _62558;
  wire _62560 = _62557 ^ _62559;
  wire _62561 = _62555 ^ _62560;
  wire _62562 = uncoded_block[1250] ^ uncoded_block[1260];
  wire _62563 = uncoded_block[1262] ^ uncoded_block[1269];
  wire _62564 = _62562 ^ _62563;
  wire _62565 = uncoded_block[1297] ^ uncoded_block[1307];
  wire _62566 = _62565 ^ _14430;
  wire _62567 = _62564 ^ _62566;
  wire _62568 = uncoded_block[1315] ^ uncoded_block[1319];
  wire _62569 = uncoded_block[1332] ^ uncoded_block[1355];
  wire _62570 = _62568 ^ _62569;
  wire _62571 = uncoded_block[1358] ^ uncoded_block[1368];
  wire _62572 = uncoded_block[1375] ^ uncoded_block[1384];
  wire _62573 = _62571 ^ _62572;
  wire _62574 = _62570 ^ _62573;
  wire _62575 = _62567 ^ _62574;
  wire _62576 = _62561 ^ _62575;
  wire _62577 = uncoded_block[1385] ^ uncoded_block[1392];
  wire _62578 = uncoded_block[1406] ^ uncoded_block[1415];
  wire _62579 = _62577 ^ _62578;
  wire _62580 = uncoded_block[1433] ^ uncoded_block[1444];
  wire _62581 = _62580 ^ _3868;
  wire _62582 = _62579 ^ _62581;
  wire _62583 = uncoded_block[1458] ^ uncoded_block[1476];
  wire _62584 = uncoded_block[1477] ^ uncoded_block[1487];
  wire _62585 = _62583 ^ _62584;
  wire _62586 = uncoded_block[1493] ^ uncoded_block[1507];
  wire _62587 = uncoded_block[1512] ^ uncoded_block[1528];
  wire _62588 = _62586 ^ _62587;
  wire _62589 = _62585 ^ _62588;
  wire _62590 = _62582 ^ _62589;
  wire _62591 = _58669 ^ _57216;
  wire _62592 = uncoded_block[1552] ^ uncoded_block[1566];
  wire _62593 = _62592 ^ _2379;
  wire _62594 = _62591 ^ _62593;
  wire _62595 = uncoded_block[1616] ^ uncoded_block[1621];
  wire _62596 = _56621 ^ _62595;
  wire _62597 = uncoded_block[1631] ^ uncoded_block[1657];
  wire _62598 = _13494 ^ _62597;
  wire _62599 = _62596 ^ _62598;
  wire _62600 = _62594 ^ _62599;
  wire _62601 = _62590 ^ _62600;
  wire _62602 = _62576 ^ _62601;
  wire _62603 = uncoded_block[1665] ^ uncoded_block[1672];
  wire _62604 = _62603 ^ _19475;
  wire _62605 = uncoded_block[1690] ^ uncoded_block[1696];
  wire _62606 = _62605 ^ _847;
  wire _62607 = _62604 ^ _62606;
  wire _62608 = _62607 ^ uncoded_block[1710];
  wire _62609 = _62602 ^ _62608;
  wire _62610 = _62550 ^ _62609;
  wire _62611 = uncoded_block[2] ^ uncoded_block[9];
  wire _62612 = uncoded_block[10] ^ uncoded_block[22];
  wire _62613 = _62611 ^ _62612;
  wire _62614 = _62613 ^ _55452;
  wire _62615 = uncoded_block[40] ^ uncoded_block[51];
  wire _62616 = uncoded_block[56] ^ uncoded_block[69];
  wire _62617 = _62615 ^ _62616;
  wire _62618 = _19511 ^ _6750;
  wire _62619 = _62617 ^ _62618;
  wire _62620 = _62614 ^ _62619;
  wire _62621 = uncoded_block[84] ^ uncoded_block[93];
  wire _62622 = uncoded_block[98] ^ uncoded_block[107];
  wire _62623 = _62621 ^ _62622;
  wire _62624 = uncoded_block[127] ^ uncoded_block[155];
  wire _62625 = _54 ^ _62624;
  wire _62626 = _62623 ^ _62625;
  wire _62627 = _73 ^ _1751;
  wire _62628 = uncoded_block[174] ^ uncoded_block[185];
  wire _62629 = _938 ^ _62628;
  wire _62630 = _62627 ^ _62629;
  wire _62631 = _62626 ^ _62630;
  wire _62632 = _62620 ^ _62631;
  wire _62633 = uncoded_block[203] ^ uncoded_block[212];
  wire _62634 = _22368 ^ _62633;
  wire _62635 = _62634 ^ _19554;
  wire _62636 = _4791 ^ _3311;
  wire _62637 = uncoded_block[257] ^ uncoded_block[264];
  wire _62638 = _62637 ^ _56436;
  wire _62639 = _62636 ^ _62638;
  wire _62640 = _62635 ^ _62639;
  wire _62641 = _5513 ^ _49687;
  wire _62642 = uncoded_block[297] ^ uncoded_block[302];
  wire _62643 = _62642 ^ _1002;
  wire _62644 = _62641 ^ _62643;
  wire _62645 = _4123 ^ _1819;
  wire _62646 = _8646 ^ _1826;
  wire _62647 = _62645 ^ _62646;
  wire _62648 = _62644 ^ _62647;
  wire _62649 = _62640 ^ _62648;
  wire _62650 = _62632 ^ _62649;
  wire _62651 = uncoded_block[360] ^ uncoded_block[372];
  wire _62652 = _2602 ^ _62651;
  wire _62653 = uncoded_block[375] ^ uncoded_block[388];
  wire _62654 = _62653 ^ _1046;
  wire _62655 = _62652 ^ _62654;
  wire _62656 = uncoded_block[402] ^ uncoded_block[410];
  wire _62657 = uncoded_block[425] ^ uncoded_block[444];
  wire _62658 = _62656 ^ _62657;
  wire _62659 = _9275 ^ _209;
  wire _62660 = _62658 ^ _62659;
  wire _62661 = _62655 ^ _62660;
  wire _62662 = _5584 ^ _15207;
  wire _62663 = uncoded_block[468] ^ uncoded_block[481];
  wire _62664 = _62663 ^ _4902;
  wire _62665 = _62662 ^ _62664;
  wire _62666 = _6921 ^ _3439;
  wire _62667 = _4921 ^ _3450;
  wire _62668 = _62666 ^ _62667;
  wire _62669 = _62665 ^ _62668;
  wire _62670 = _62661 ^ _62669;
  wire _62671 = _1906 ^ _48151;
  wire _62672 = uncoded_block[556] ^ uncoded_block[560];
  wire _62673 = uncoded_block[561] ^ uncoded_block[568];
  wire _62674 = _62672 ^ _62673;
  wire _62675 = _62671 ^ _62674;
  wire _62676 = uncoded_block[569] ^ uncoded_block[578];
  wire _62677 = uncoded_block[580] ^ uncoded_block[588];
  wire _62678 = _62676 ^ _62677;
  wire _62679 = _4234 ^ _59489;
  wire _62680 = _62678 ^ _62679;
  wire _62681 = _62675 ^ _62680;
  wire _62682 = uncoded_block[623] ^ uncoded_block[630];
  wire _62683 = _4960 ^ _62682;
  wire _62684 = _1161 ^ _4972;
  wire _62685 = _62683 ^ _62684;
  wire _62686 = uncoded_block[651] ^ uncoded_block[658];
  wire _62687 = _62686 ^ _4261;
  wire _62688 = uncoded_block[670] ^ uncoded_block[675];
  wire _62689 = _62688 ^ _8177;
  wire _62690 = _62687 ^ _62689;
  wire _62691 = _62685 ^ _62690;
  wire _62692 = _62681 ^ _62691;
  wire _62693 = _62670 ^ _62692;
  wire _62694 = _62650 ^ _62693;
  wire _62695 = uncoded_block[688] ^ uncoded_block[695];
  wire _62696 = uncoded_block[696] ^ uncoded_block[706];
  wire _62697 = _62695 ^ _62696;
  wire _62698 = uncoded_block[723] ^ uncoded_block[735];
  wire _62699 = _23863 ^ _62698;
  wire _62700 = _62697 ^ _62699;
  wire _62701 = _11009 ^ _13752;
  wire _62702 = _16775 ^ _2003;
  wire _62703 = _62701 ^ _62702;
  wire _62704 = _62700 ^ _62703;
  wire _62705 = uncoded_block[763] ^ uncoded_block[778];
  wire _62706 = _62705 ^ _2794;
  wire _62707 = uncoded_block[790] ^ uncoded_block[813];
  wire _62708 = _1224 ^ _62707;
  wire _62709 = _62706 ^ _62708;
  wire _62710 = _60831 ^ _17797;
  wire _62711 = _2036 ^ _11609;
  wire _62712 = _62710 ^ _62711;
  wire _62713 = _62709 ^ _62712;
  wire _62714 = _62704 ^ _62713;
  wire _62715 = _46711 ^ _8812;
  wire _62716 = uncoded_block[868] ^ uncoded_block[887];
  wire _62717 = _17804 ^ _62716;
  wire _62718 = _62715 ^ _62717;
  wire _62719 = uncoded_block[926] ^ uncoded_block[934];
  wire _62720 = _54408 ^ _62719;
  wire _62721 = _22105 ^ _460;
  wire _62722 = _62720 ^ _62721;
  wire _62723 = _62718 ^ _62722;
  wire _62724 = uncoded_block[964] ^ uncoded_block[968];
  wire _62725 = _19748 ^ _62724;
  wire _62726 = _8283 ^ _5114;
  wire _62727 = _62725 ^ _62726;
  wire _62728 = _47490 ^ _1330;
  wire _62729 = uncoded_block[1039] ^ uncoded_block[1053];
  wire _62730 = _34925 ^ _62729;
  wire _62731 = _62728 ^ _62730;
  wire _62732 = _62727 ^ _62731;
  wire _62733 = _62723 ^ _62732;
  wire _62734 = _62714 ^ _62733;
  wire _62735 = uncoded_block[1061] ^ uncoded_block[1082];
  wire _62736 = _62735 ^ _27515;
  wire _62737 = uncoded_block[1099] ^ uncoded_block[1106];
  wire _62738 = _62737 ^ _11147;
  wire _62739 = _62736 ^ _62738;
  wire _62740 = _4459 ^ _9496;
  wire _62741 = uncoded_block[1141] ^ uncoded_block[1148];
  wire _62742 = _62741 ^ _11157;
  wire _62743 = _62740 ^ _62742;
  wire _62744 = _62739 ^ _62743;
  wire _62745 = _6511 ^ _18382;
  wire _62746 = _61698 ^ _590;
  wire _62747 = _62745 ^ _62746;
  wire _62748 = uncoded_block[1185] ^ uncoded_block[1190];
  wire _62749 = _62748 ^ _4488;
  wire _62750 = _2979 ^ _23105;
  wire _62751 = _62749 ^ _62750;
  wire _62752 = _62747 ^ _62751;
  wire _62753 = _62744 ^ _62752;
  wire _62754 = _6532 ^ _5219;
  wire _62755 = uncoded_block[1254] ^ uncoded_block[1260];
  wire _62756 = _62755 ^ _30361;
  wire _62757 = _62754 ^ _62756;
  wire _62758 = uncoded_block[1266] ^ uncoded_block[1282];
  wire _62759 = _62758 ^ _4529;
  wire _62760 = uncoded_block[1294] ^ uncoded_block[1305];
  wire _62761 = _8399 ^ _62760;
  wire _62762 = _62759 ^ _62761;
  wire _62763 = _62757 ^ _62762;
  wire _62764 = uncoded_block[1311] ^ uncoded_block[1329];
  wire _62765 = uncoded_block[1333] ^ uncoded_block[1340];
  wire _62766 = _62764 ^ _62765;
  wire _62767 = uncoded_block[1348] ^ uncoded_block[1364];
  wire _62768 = _12854 ^ _62767;
  wire _62769 = _62766 ^ _62768;
  wire _62770 = uncoded_block[1366] ^ uncoded_block[1371];
  wire _62771 = uncoded_block[1375] ^ uncoded_block[1381];
  wire _62772 = _62770 ^ _62771;
  wire _62773 = uncoded_block[1388] ^ uncoded_block[1395];
  wire _62774 = _12307 ^ _62773;
  wire _62775 = _62772 ^ _62774;
  wire _62776 = _62769 ^ _62775;
  wire _62777 = _62763 ^ _62776;
  wire _62778 = _62753 ^ _62777;
  wire _62779 = _62734 ^ _62778;
  wire _62780 = _62694 ^ _62779;
  wire _62781 = uncoded_block[1413] ^ uncoded_block[1420];
  wire _62782 = _4578 ^ _62781;
  wire _62783 = _62782 ^ _23166;
  wire _62784 = _13951 ^ _20355;
  wire _62785 = uncoded_block[1458] ^ uncoded_block[1473];
  wire _62786 = _44727 ^ _62785;
  wire _62787 = _62784 ^ _62786;
  wire _62788 = _62783 ^ _62787;
  wire _62789 = uncoded_block[1475] ^ uncoded_block[1486];
  wire _62790 = _62789 ^ _60095;
  wire _62791 = _25430 ^ _3112;
  wire _62792 = _62790 ^ _62791;
  wire _62793 = _56921 ^ _6651;
  wire _62794 = _3918 ^ _1615;
  wire _62795 = _62793 ^ _62794;
  wire _62796 = _62792 ^ _62795;
  wire _62797 = _62788 ^ _62796;
  wire _62798 = _30875 ^ _11294;
  wire _62799 = uncoded_block[1606] ^ uncoded_block[1617];
  wire _62800 = uncoded_block[1619] ^ uncoded_block[1627];
  wire _62801 = _62799 ^ _62800;
  wire _62802 = _62798 ^ _62801;
  wire _62803 = uncoded_block[1630] ^ uncoded_block[1637];
  wire _62804 = _1636 ^ _62803;
  wire _62805 = uncoded_block[1643] ^ uncoded_block[1653];
  wire _62806 = _62805 ^ _10760;
  wire _62807 = _62804 ^ _62806;
  wire _62808 = _62802 ^ _62807;
  wire _62809 = uncoded_block[1667] ^ uncoded_block[1695];
  wire _62810 = _62809 ^ _20920;
  wire _62811 = _45907 ^ _62810;
  wire _62812 = _55812 ^ uncoded_block[1717];
  wire _62813 = _62811 ^ _62812;
  wire _62814 = _62808 ^ _62813;
  wire _62815 = _62797 ^ _62814;
  wire _62816 = _62780 ^ _62815;
  wire _62817 = _10787 ^ _61987;
  wire _62818 = _25941 ^ _58050;
  wire _62819 = _62817 ^ _62818;
  wire _62820 = _7966 ^ _34689;
  wire _62821 = uncoded_block[82] ^ uncoded_block[88];
  wire _62822 = _28765 ^ _62821;
  wire _62823 = _62820 ^ _62822;
  wire _62824 = _62819 ^ _62823;
  wire _62825 = _57271 ^ _6116;
  wire _62826 = uncoded_block[106] ^ uncoded_block[117];
  wire _62827 = uncoded_block[119] ^ uncoded_block[131];
  wire _62828 = _62826 ^ _62827;
  wire _62829 = _62825 ^ _62828;
  wire _62830 = _25075 ^ _15620;
  wire _62831 = _24178 ^ _53600;
  wire _62832 = _62830 ^ _62831;
  wire _62833 = _62829 ^ _62832;
  wire _62834 = _62824 ^ _62833;
  wire _62835 = uncoded_block[155] ^ uncoded_block[170];
  wire _62836 = _5469 ^ _62835;
  wire _62837 = _59682 ^ _3283;
  wire _62838 = _62836 ^ _62837;
  wire _62839 = uncoded_block[196] ^ uncoded_block[202];
  wire _62840 = _62839 ^ _30963;
  wire _62841 = _59688 ^ _34724;
  wire _62842 = _62840 ^ _62841;
  wire _62843 = _62838 ^ _62842;
  wire _62844 = _59691 ^ _4084;
  wire _62845 = _14116 ^ _31834;
  wire _62846 = _62844 ^ _62845;
  wire _62847 = uncoded_block[261] ^ uncoded_block[271];
  wire _62848 = _62847 ^ _10303;
  wire _62849 = uncoded_block[287] ^ uncoded_block[293];
  wire _62850 = _5515 ^ _62849;
  wire _62851 = _62848 ^ _62850;
  wire _62852 = _62846 ^ _62851;
  wire _62853 = _62843 ^ _62852;
  wire _62854 = _62834 ^ _62853;
  wire _62855 = _28065 ^ _3337;
  wire _62856 = _59706 ^ _33112;
  wire _62857 = _62855 ^ _62856;
  wire _62858 = uncoded_block[336] ^ uncoded_block[344];
  wire _62859 = _62858 ^ _8652;
  wire _62860 = _19092 ^ _10898;
  wire _62861 = _62859 ^ _62860;
  wire _62862 = _62857 ^ _62861;
  wire _62863 = uncoded_block[410] ^ uncoded_block[421];
  wire _62864 = _62863 ^ _37209;
  wire _62865 = _59713 ^ _62864;
  wire _62866 = _27350 ^ _12559;
  wire _62867 = uncoded_block[452] ^ uncoded_block[460];
  wire _62868 = _58123 ^ _62867;
  wire _62869 = _62866 ^ _62868;
  wire _62870 = _62865 ^ _62869;
  wire _62871 = _62862 ^ _62870;
  wire _62872 = _13665 ^ _59726;
  wire _62873 = _8694 ^ _4195;
  wire _62874 = _62872 ^ _62873;
  wire _62875 = uncoded_block[519] ^ uncoded_block[526];
  wire _62876 = _8705 ^ _62875;
  wire _62877 = _59731 ^ _62876;
  wire _62878 = _62874 ^ _62877;
  wire _62879 = uncoded_block[535] ^ uncoded_block[545];
  wire _62880 = _26081 ^ _62879;
  wire _62881 = _62880 ^ _58141;
  wire _62882 = uncoded_block[575] ^ uncoded_block[584];
  wire _62883 = _62882 ^ _58147;
  wire _62884 = _12608 ^ _23400;
  wire _62885 = _62883 ^ _62884;
  wire _62886 = _62881 ^ _62885;
  wire _62887 = _62878 ^ _62886;
  wire _62888 = _62871 ^ _62887;
  wire _62889 = _62854 ^ _62888;
  wire _62890 = _44924 ^ _34028;
  wire _62891 = _59750 ^ _62890;
  wire _62892 = _16752 ^ _33194;
  wire _62893 = _58158 ^ _62892;
  wire _62894 = _62891 ^ _62893;
  wire _62895 = _19191 ^ _18249;
  wire _62896 = _1186 ^ _14766;
  wire _62897 = _62895 ^ _62896;
  wire _62898 = _48929 ^ _59764;
  wire _62899 = _62898 ^ _59766;
  wire _62900 = _62897 ^ _62899;
  wire _62901 = _62894 ^ _62900;
  wire _62902 = _32372 ^ _31542;
  wire _62903 = _59769 ^ _62902;
  wire _62904 = _5723 ^ _22071;
  wire _62905 = _32377 ^ _62904;
  wire _62906 = _62903 ^ _62905;
  wire _62907 = _16791 ^ _16793;
  wire _62908 = _7632 ^ _7634;
  wire _62909 = _62907 ^ _62908;
  wire _62910 = _59782 ^ _33239;
  wire _62911 = uncoded_block[851] ^ uncoded_block[860];
  wire _62912 = _62911 ^ _2827;
  wire _62913 = _62910 ^ _62912;
  wire _62914 = _62909 ^ _62913;
  wire _62915 = _62906 ^ _62914;
  wire _62916 = _62901 ^ _62915;
  wire _62917 = uncoded_block[868] ^ uncoded_block[890];
  wire _62918 = _62917 ^ _31988;
  wire _62919 = _62918 ^ _1286;
  wire _62920 = _12712 ^ _2073;
  wire _62921 = _29379 ^ _9971;
  wire _62922 = _62920 ^ _62921;
  wire _62923 = _62919 ^ _62922;
  wire _62924 = uncoded_block[947] ^ uncoded_block[956];
  wire _62925 = uncoded_block[964] ^ uncoded_block[971];
  wire _62926 = _62924 ^ _62925;
  wire _62927 = _5112 ^ _5114;
  wire _62928 = _62926 ^ _62927;
  wire _62929 = _7093 ^ _2105;
  wire _62930 = uncoded_block[994] ^ uncoded_block[1001];
  wire _62931 = _62930 ^ _22122;
  wire _62932 = _62929 ^ _62931;
  wire _62933 = _62928 ^ _62932;
  wire _62934 = _62923 ^ _62933;
  wire _62935 = _2890 ^ _2894;
  wire _62936 = uncoded_block[1037] ^ uncoded_block[1042];
  wire _62937 = _2127 ^ _62936;
  wire _62938 = _62935 ^ _62937;
  wire _62939 = _1356 ^ _8311;
  wire _62940 = _62939 ^ _59818;
  wire _62941 = _62938 ^ _62940;
  wire _62942 = _5163 ^ _13857;
  wire _62943 = uncoded_block[1096] ^ uncoded_block[1101];
  wire _62944 = _62943 ^ _8914;
  wire _62945 = _62942 ^ _62944;
  wire _62946 = uncoded_block[1111] ^ uncoded_block[1125];
  wire _62947 = _62946 ^ _13866;
  wire _62948 = uncoded_block[1135] ^ uncoded_block[1151];
  wire _62949 = _62948 ^ _577;
  wire _62950 = _62947 ^ _62949;
  wire _62951 = _62945 ^ _62950;
  wire _62952 = _62941 ^ _62951;
  wire _62953 = _62934 ^ _62952;
  wire _62954 = _62916 ^ _62953;
  wire _62955 = _62889 ^ _62954;
  wire _62956 = _59827 ^ _59830;
  wire _62957 = _46078 ^ _60701;
  wire _62958 = _35360 ^ _50262;
  wire _62959 = _62957 ^ _62958;
  wire _62960 = _62956 ^ _62959;
  wire _62961 = _15927 ^ _59838;
  wire _62962 = _2232 ^ _59840;
  wire _62963 = _62961 ^ _62962;
  wire _62964 = uncoded_block[1261] ^ uncoded_block[1268];
  wire _62965 = _62964 ^ _16419;
  wire _62966 = _7792 ^ _59848;
  wire _62967 = _62965 ^ _62966;
  wire _62968 = _62963 ^ _62967;
  wire _62969 = _62960 ^ _62968;
  wire _62970 = uncoded_block[1308] ^ uncoded_block[1313];
  wire _62971 = _20812 ^ _62970;
  wire _62972 = _6574 ^ _29481;
  wire _62973 = _62971 ^ _62972;
  wire _62974 = _9564 ^ _5269;
  wire _62975 = _3035 ^ _62974;
  wire _62976 = _62973 ^ _62975;
  wire _62977 = _33363 ^ _5273;
  wire _62978 = uncoded_block[1361] ^ uncoded_block[1381];
  wire _62979 = _62978 ^ _59860;
  wire _62980 = _62977 ^ _62979;
  wire _62981 = _3846 ^ _1523;
  wire _62982 = _59865 ^ _62981;
  wire _62983 = _62980 ^ _62982;
  wire _62984 = _62976 ^ _62983;
  wire _62985 = _62969 ^ _62984;
  wire _62986 = _59867 ^ _7844;
  wire _62987 = _47970 ^ _59872;
  wire _62988 = _62986 ^ _62987;
  wire _62989 = _59873 ^ _14985;
  wire _62990 = uncoded_block[1473] ^ uncoded_block[1488];
  wire _62991 = _20855 ^ _62990;
  wire _62992 = _62989 ^ _62991;
  wire _62993 = _62988 ^ _62992;
  wire _62994 = _7259 ^ _5334;
  wire _62995 = _58295 ^ _62994;
  wire _62996 = _19429 ^ _4620;
  wire _62997 = _62996 ^ _59888;
  wire _62998 = _62995 ^ _62997;
  wire _62999 = _62993 ^ _62998;
  wire _63000 = _15009 ^ _7274;
  wire _63001 = uncoded_block[1568] ^ uncoded_block[1580];
  wire _63002 = _13472 ^ _63001;
  wire _63003 = _63000 ^ _63002;
  wire _63004 = uncoded_block[1581] ^ uncoded_block[1589];
  wire _63005 = _63004 ^ _791;
  wire _63006 = uncoded_block[1611] ^ uncoded_block[1624];
  wire _63007 = _800 ^ _63006;
  wire _63008 = _63005 ^ _63007;
  wire _63009 = _63003 ^ _63008;
  wire _63010 = _12947 ^ _7306;
  wire _63011 = uncoded_block[1648] ^ uncoded_block[1652];
  wire _63012 = _12955 ^ _63011;
  wire _63013 = _63010 ^ _63012;
  wire _63014 = uncoded_block[1669] ^ uncoded_block[1675];
  wire _63015 = _4687 ^ _63014;
  wire _63016 = uncoded_block[1698] ^ uncoded_block[1706];
  wire _63017 = _63016 ^ _39871;
  wire _63018 = _63015 ^ _63017;
  wire _63019 = _63013 ^ _63018;
  wire _63020 = _63009 ^ _63019;
  wire _63021 = _62999 ^ _63020;
  wire _63022 = _62985 ^ _63021;
  wire _63023 = _63022 ^ _4704;
  wire _63024 = _62955 ^ _63023;
  wire _63025 = uncoded_block[6] ^ uncoded_block[16];
  wire _63026 = uncoded_block[57] ^ uncoded_block[73];
  wire _63027 = _63025 ^ _63026;
  wire _63028 = uncoded_block[78] ^ uncoded_block[91];
  wire _63029 = uncoded_block[95] ^ uncoded_block[109];
  wire _63030 = _63028 ^ _63029;
  wire _63031 = _63027 ^ _63030;
  wire _63032 = _29611 ^ _15114;
  wire _63033 = uncoded_block[147] ^ uncoded_block[164];
  wire _63034 = uncoded_block[172] ^ uncoded_block[196];
  wire _63035 = _63033 ^ _63034;
  wire _63036 = _63032 ^ _63035;
  wire _63037 = _63031 ^ _63036;
  wire _63038 = uncoded_block[204] ^ uncoded_block[218];
  wire _63039 = _63038 ^ _29642;
  wire _63040 = uncoded_block[258] ^ uncoded_block[271];
  wire _63041 = _44837 ^ _63040;
  wire _63042 = _63039 ^ _63041;
  wire _63043 = uncoded_block[284] ^ uncoded_block[299];
  wire _63044 = _63043 ^ _17639;
  wire _63045 = uncoded_block[309] ^ uncoded_block[318];
  wire _63046 = uncoded_block[341] ^ uncoded_block[357];
  wire _63047 = _63045 ^ _63046;
  wire _63048 = _63044 ^ _63047;
  wire _63049 = _63042 ^ _63048;
  wire _63050 = _63037 ^ _63049;
  wire _63051 = uncoded_block[359] ^ uncoded_block[367];
  wire _63052 = uncoded_block[368] ^ uncoded_block[373];
  wire _63053 = _63051 ^ _63052;
  wire _63054 = uncoded_block[400] ^ uncoded_block[410];
  wire _63055 = _1849 ^ _63054;
  wire _63056 = _63053 ^ _63055;
  wire _63057 = uncoded_block[423] ^ uncoded_block[443];
  wire _63058 = _63057 ^ _3411;
  wire _63059 = uncoded_block[465] ^ uncoded_block[477];
  wire _63060 = _63059 ^ _9837;
  wire _63061 = _63058 ^ _63060;
  wire _63062 = _63056 ^ _63061;
  wire _63063 = uncoded_block[537] ^ uncoded_block[558];
  wire _63064 = _63063 ^ _1931;
  wire _63065 = _50113 ^ _63064;
  wire _63066 = uncoded_block[602] ^ uncoded_block[609];
  wire _63067 = uncoded_block[613] ^ uncoded_block[620];
  wire _63068 = _63066 ^ _63067;
  wire _63069 = uncoded_block[632] ^ uncoded_block[649];
  wire _63070 = uncoded_block[659] ^ uncoded_block[673];
  wire _63071 = _63069 ^ _63070;
  wire _63072 = _63068 ^ _63071;
  wire _63073 = _63065 ^ _63072;
  wire _63074 = _63062 ^ _63073;
  wire _63075 = _63050 ^ _63074;
  wire _63076 = uncoded_block[678] ^ uncoded_block[691];
  wire _63077 = uncoded_block[701] ^ uncoded_block[713];
  wire _63078 = _63076 ^ _63077;
  wire _63079 = uncoded_block[721] ^ uncoded_block[743];
  wire _63080 = _63079 ^ _58821;
  wire _63081 = _63078 ^ _63080;
  wire _63082 = uncoded_block[772] ^ uncoded_block[787];
  wire _63083 = _1217 ^ _63082;
  wire _63084 = uncoded_block[791] ^ uncoded_block[802];
  wire _63085 = uncoded_block[805] ^ uncoded_block[831];
  wire _63086 = _63084 ^ _63085;
  wire _63087 = _63083 ^ _63086;
  wire _63088 = _63081 ^ _63087;
  wire _63089 = uncoded_block[856] ^ uncoded_block[876];
  wire _63090 = _26164 ^ _63089;
  wire _63091 = uncoded_block[881] ^ uncoded_block[895];
  wire _63092 = _63091 ^ _4368;
  wire _63093 = _63090 ^ _63092;
  wire _63094 = uncoded_block[938] ^ uncoded_block[951];
  wire _63095 = _2858 ^ _63094;
  wire _63096 = uncoded_block[965] ^ uncoded_block[971];
  wire _63097 = uncoded_block[977] ^ uncoded_block[992];
  wire _63098 = _63096 ^ _63097;
  wire _63099 = _63095 ^ _63098;
  wire _63100 = _63093 ^ _63099;
  wire _63101 = _63088 ^ _63100;
  wire _63102 = uncoded_block[998] ^ uncoded_block[1024];
  wire _63103 = _63102 ^ _9455;
  wire _63104 = uncoded_block[1037] ^ uncoded_block[1053];
  wire _63105 = _63104 ^ _38137;
  wire _63106 = _63103 ^ _63105;
  wire _63107 = uncoded_block[1079] ^ uncoded_block[1093];
  wire _63108 = uncoded_block[1100] ^ uncoded_block[1108];
  wire _63109 = _63107 ^ _63108;
  wire _63110 = uncoded_block[1121] ^ uncoded_block[1129];
  wire _63111 = _7132 ^ _63110;
  wire _63112 = _63109 ^ _63111;
  wire _63113 = _63106 ^ _63112;
  wire _63114 = uncoded_block[1156] ^ uncoded_block[1172];
  wire _63115 = _4462 ^ _63114;
  wire _63116 = uncoded_block[1191] ^ uncoded_block[1203];
  wire _63117 = uncoded_block[1207] ^ uncoded_block[1217];
  wire _63118 = _63116 ^ _63117;
  wire _63119 = _63115 ^ _63118;
  wire _63120 = uncoded_block[1238] ^ uncoded_block[1249];
  wire _63121 = _59835 ^ _63120;
  wire _63122 = uncoded_block[1272] ^ uncoded_block[1287];
  wire _63123 = _63122 ^ _10646;
  wire _63124 = _63121 ^ _63123;
  wire _63125 = _63119 ^ _63124;
  wire _63126 = _63113 ^ _63125;
  wire _63127 = _63101 ^ _63126;
  wire _63128 = _63075 ^ _63127;
  wire _63129 = uncoded_block[1309] ^ uncoded_block[1317];
  wire _63130 = uncoded_block[1320] ^ uncoded_block[1335];
  wire _63131 = _63129 ^ _63130;
  wire _63132 = uncoded_block[1339] ^ uncoded_block[1351];
  wire _63133 = _63132 ^ _11220;
  wire _63134 = _63131 ^ _63133;
  wire _63135 = uncoded_block[1359] ^ uncoded_block[1392];
  wire _63136 = _63135 ^ _15970;
  wire _63137 = uncoded_block[1404] ^ uncoded_block[1447];
  wire _63138 = uncoded_block[1451] ^ uncoded_block[1457];
  wire _63139 = _63137 ^ _63138;
  wire _63140 = _63136 ^ _63139;
  wire _63141 = _63134 ^ _63140;
  wire _63142 = uncoded_block[1459] ^ uncoded_block[1468];
  wire _63143 = _63142 ^ _1551;
  wire _63144 = _13966 ^ _36653;
  wire _63145 = _63143 ^ _63144;
  wire _63146 = uncoded_block[1523] ^ uncoded_block[1538];
  wire _63147 = uncoded_block[1546] ^ uncoded_block[1555];
  wire _63148 = _63146 ^ _63147;
  wire _63149 = uncoded_block[1597] ^ uncoded_block[1618];
  wire _63150 = _774 ^ _63149;
  wire _63151 = _63148 ^ _63150;
  wire _63152 = _63145 ^ _63151;
  wire _63153 = _63141 ^ _63152;
  wire _63154 = uncoded_block[1639] ^ uncoded_block[1683];
  wire _63155 = _11853 ^ _63154;
  wire _63156 = uncoded_block[1697] ^ uncoded_block[1713];
  wire _63157 = _20429 ^ _63156;
  wire _63158 = _63155 ^ _63157;
  wire _63159 = _33025 ^ uncoded_block[1722];
  wire _63160 = _63158 ^ _63159;
  wire _63161 = _63153 ^ _63160;
  wire _63162 = _63128 ^ _63161;
  wire _63163 = uncoded_block[13] ^ uncoded_block[22];
  wire _63164 = _1683 ^ _63163;
  wire _63165 = uncoded_block[30] ^ uncoded_block[41];
  wire _63166 = _9694 ^ _63165;
  wire _63167 = _63164 ^ _63166;
  wire _63168 = _22 ^ _7968;
  wire _63169 = uncoded_block[56] ^ uncoded_block[61];
  wire _63170 = _63169 ^ _2474;
  wire _63171 = _63168 ^ _63170;
  wire _63172 = _63167 ^ _63171;
  wire _63173 = _7367 ^ _11904;
  wire _63174 = _6755 ^ _5449;
  wire _63175 = _63173 ^ _63174;
  wire _63176 = _1721 ^ _46546;
  wire _63177 = _3256 ^ _21898;
  wire _63178 = _63176 ^ _63177;
  wire _63179 = _63175 ^ _63178;
  wire _63180 = _63172 ^ _63179;
  wire _63181 = uncoded_block[140] ^ uncoded_block[144];
  wire _63182 = _20969 ^ _63181;
  wire _63183 = _9182 ^ _21906;
  wire _63184 = _63182 ^ _63183;
  wire _63185 = _2517 ^ _5476;
  wire _63186 = uncoded_block[181] ^ uncoded_block[189];
  wire _63187 = _63186 ^ _13038;
  wire _63188 = _63185 ^ _63187;
  wire _63189 = _63184 ^ _63188;
  wire _63190 = _1766 ^ _6161;
  wire _63191 = _39928 ^ _6814;
  wire _63192 = _63190 ^ _63191;
  wire _63193 = _33088 ^ _9761;
  wire _63194 = uncoded_block[258] ^ uncoded_block[265];
  wire _63195 = _63194 ^ _4099;
  wire _63196 = _63193 ^ _63195;
  wire _63197 = _63192 ^ _63196;
  wire _63198 = _63189 ^ _63197;
  wire _63199 = _63180 ^ _63198;
  wire _63200 = _49519 ^ _12516;
  wire _63201 = _10875 ^ _63200;
  wire _63202 = uncoded_block[316] ^ uncoded_block[323];
  wire _63203 = uncoded_block[324] ^ uncoded_block[330];
  wire _63204 = _63202 ^ _63203;
  wire _63205 = uncoded_block[340] ^ uncoded_block[351];
  wire _63206 = uncoded_block[352] ^ uncoded_block[358];
  wire _63207 = _63205 ^ _63206;
  wire _63208 = _63204 ^ _63207;
  wire _63209 = _63201 ^ _63208;
  wire _63210 = _8075 ^ _4854;
  wire _63211 = _6235 ^ _3380;
  wire _63212 = _63210 ^ _63211;
  wire _63213 = uncoded_block[388] ^ uncoded_block[395];
  wire _63214 = _63213 ^ _2626;
  wire _63215 = _19613 ^ _2638;
  wire _63216 = _63214 ^ _63215;
  wire _63217 = _63212 ^ _63216;
  wire _63218 = _63209 ^ _63217;
  wire _63219 = uncoded_block[433] ^ uncoded_block[442];
  wire _63220 = _63219 ^ _20574;
  wire _63221 = _8681 ^ _6906;
  wire _63222 = _63220 ^ _63221;
  wire _63223 = _59473 ^ _7516;
  wire _63224 = _6277 ^ _19135;
  wire _63225 = _63223 ^ _63224;
  wire _63226 = _63222 ^ _63225;
  wire _63227 = _6922 ^ _7531;
  wire _63228 = uncoded_block[518] ^ uncoded_block[525];
  wire _63229 = _8122 ^ _63228;
  wire _63230 = _63227 ^ _63229;
  wire _63231 = _60972 ^ _55228;
  wire _63232 = uncoded_block[563] ^ uncoded_block[570];
  wire _63233 = _52786 ^ _63232;
  wire _63234 = _63231 ^ _63233;
  wire _63235 = _63230 ^ _63234;
  wire _63236 = _63226 ^ _63235;
  wire _63237 = _63218 ^ _63236;
  wire _63238 = _63199 ^ _63237;
  wire _63239 = _6945 ^ _8143;
  wire _63240 = uncoded_block[588] ^ uncoded_block[593];
  wire _63241 = _63240 ^ _6952;
  wire _63242 = _63239 ^ _63241;
  wire _63243 = _63242 ^ _6962;
  wire _63244 = uncoded_block[634] ^ uncoded_block[640];
  wire _63245 = _8159 ^ _63244;
  wire _63246 = _296 ^ _19181;
  wire _63247 = _63245 ^ _63246;
  wire _63248 = uncoded_block[671] ^ uncoded_block[677];
  wire _63249 = _4264 ^ _63248;
  wire _63250 = uncoded_block[678] ^ uncoded_block[682];
  wire _63251 = uncoded_block[684] ^ uncoded_block[691];
  wire _63252 = _63250 ^ _63251;
  wire _63253 = _63249 ^ _63252;
  wire _63254 = _63247 ^ _63253;
  wire _63255 = _63243 ^ _63254;
  wire _63256 = uncoded_block[692] ^ uncoded_block[704];
  wire _63257 = _63256 ^ _46294;
  wire _63258 = _1983 ^ _51258;
  wire _63259 = _63257 ^ _63258;
  wire _63260 = uncoded_block[726] ^ uncoded_block[739];
  wire _63261 = _63260 ^ _21600;
  wire _63262 = _61467 ^ _9914;
  wire _63263 = _63261 ^ _63262;
  wire _63264 = _63259 ^ _63263;
  wire _63265 = _1221 ^ _19217;
  wire _63266 = _3570 ^ _7622;
  wire _63267 = _63265 ^ _63266;
  wire _63268 = uncoded_block[798] ^ uncoded_block[807];
  wire _63269 = _11024 ^ _63268;
  wire _63270 = uncoded_block[815] ^ uncoded_block[822];
  wire _63271 = _11029 ^ _63270;
  wire _63272 = _63269 ^ _63271;
  wire _63273 = _63267 ^ _63272;
  wire _63274 = _63264 ^ _63273;
  wire _63275 = _63255 ^ _63274;
  wire _63276 = uncoded_block[835] ^ uncoded_block[841];
  wire _63277 = uncoded_block[849] ^ uncoded_block[859];
  wire _63278 = _63276 ^ _63277;
  wire _63279 = _41994 ^ _63278;
  wire _63280 = _2824 ^ _16815;
  wire _63281 = _11059 ^ _45738;
  wire _63282 = _63280 ^ _63281;
  wire _63283 = _63279 ^ _63282;
  wire _63284 = _428 ^ _18311;
  wire _63285 = uncoded_block[912] ^ uncoded_block[923];
  wire _63286 = _3623 ^ _63285;
  wire _63287 = _63284 ^ _63286;
  wire _63288 = _3637 ^ _2863;
  wire _63289 = uncoded_block[947] ^ uncoded_block[955];
  wire _63290 = uncoded_block[958] ^ uncoded_block[962];
  wire _63291 = _63289 ^ _63290;
  wire _63292 = _63288 ^ _63291;
  wire _63293 = _63287 ^ _63292;
  wire _63294 = _63283 ^ _63293;
  wire _63295 = uncoded_block[972] ^ uncoded_block[977];
  wire _63296 = _63295 ^ _57438;
  wire _63297 = _63296 ^ _38920;
  wire _63298 = uncoded_block[994] ^ uncoded_block[1012];
  wire _63299 = _63298 ^ _2893;
  wire _63300 = uncoded_block[1019] ^ uncoded_block[1027];
  wire _63301 = uncoded_block[1029] ^ uncoded_block[1035];
  wire _63302 = _63300 ^ _63301;
  wire _63303 = _63299 ^ _63302;
  wire _63304 = _63297 ^ _63303;
  wire _63305 = _23498 ^ _23964;
  wire _63306 = _7117 ^ _1366;
  wire _63307 = _63305 ^ _63306;
  wire _63308 = _12770 ^ _26664;
  wire _63309 = uncoded_block[1102] ^ uncoded_block[1109];
  wire _63310 = _5843 ^ _63309;
  wire _63311 = _63308 ^ _63310;
  wire _63312 = _63307 ^ _63311;
  wire _63313 = _63304 ^ _63312;
  wire _63314 = _63294 ^ _63313;
  wire _63315 = _63275 ^ _63314;
  wire _63316 = _63238 ^ _63315;
  wire _63317 = uncoded_block[1114] ^ uncoded_block[1122];
  wire _63318 = uncoded_block[1123] ^ uncoded_block[1133];
  wire _63319 = _63317 ^ _63318;
  wire _63320 = uncoded_block[1137] ^ uncoded_block[1143];
  wire _63321 = _63320 ^ _574;
  wire _63322 = _63319 ^ _63321;
  wire _63323 = uncoded_block[1148] ^ uncoded_block[1158];
  wire _63324 = uncoded_block[1159] ^ uncoded_block[1165];
  wire _63325 = _63323 ^ _63324;
  wire _63326 = _2192 ^ _58887;
  wire _63327 = _63325 ^ _63326;
  wire _63328 = _63322 ^ _63327;
  wire _63329 = _14398 ^ _30344;
  wire _63330 = _30766 ^ _63329;
  wire _63331 = uncoded_block[1222] ^ uncoded_block[1239];
  wire _63332 = _63331 ^ _5229;
  wire _63333 = _7780 ^ _3008;
  wire _63334 = _63332 ^ _63333;
  wire _63335 = _63330 ^ _63334;
  wire _63336 = _63328 ^ _63335;
  wire _63337 = _6554 ^ _57499;
  wire _63338 = _28317 ^ _18866;
  wire _63339 = _63337 ^ _63338;
  wire _63340 = _3017 ^ _5917;
  wire _63341 = uncoded_block[1322] ^ uncoded_block[1328];
  wire _63342 = _20314 ^ _63341;
  wire _63343 = _63340 ^ _63342;
  wire _63344 = _63339 ^ _63343;
  wire _63345 = uncoded_block[1330] ^ uncoded_block[1340];
  wire _63346 = uncoded_block[1345] ^ uncoded_block[1348];
  wire _63347 = _63345 ^ _63346;
  wire _63348 = _25393 ^ _10665;
  wire _63349 = _63347 ^ _63348;
  wire _63350 = _12302 ^ _1509;
  wire _63351 = _58634 ^ _2293;
  wire _63352 = _63350 ^ _63351;
  wire _63353 = _63349 ^ _63352;
  wire _63354 = _63344 ^ _63353;
  wire _63355 = _63336 ^ _63354;
  wire _63356 = uncoded_block[1398] ^ uncoded_block[1404];
  wire _63357 = uncoded_block[1413] ^ uncoded_block[1422];
  wire _63358 = _63356 ^ _63357;
  wire _63359 = _14466 ^ _29508;
  wire _63360 = _63358 ^ _63359;
  wire _63361 = uncoded_block[1445] ^ uncoded_block[1458];
  wire _63362 = _10130 ^ _63361;
  wire _63363 = _3093 ^ _1555;
  wire _63364 = _63362 ^ _63363;
  wire _63365 = _63360 ^ _63364;
  wire _63366 = _43199 ^ _27184;
  wire _63367 = _63366 ^ _7257;
  wire _63368 = _1571 ^ _18478;
  wire _63369 = _63368 ^ _34222;
  wire _63370 = _63367 ^ _63369;
  wire _63371 = _63365 ^ _63370;
  wire _63372 = uncoded_block[1525] ^ uncoded_block[1530];
  wire _63373 = _5999 ^ _63372;
  wire _63374 = _3905 ^ _15009;
  wire _63375 = _63373 ^ _63374;
  wire _63376 = uncoded_block[1554] ^ uncoded_block[1560];
  wire _63377 = uncoded_block[1565] ^ uncoded_block[1576];
  wire _63378 = _63376 ^ _63377;
  wire _63379 = _47615 ^ _63378;
  wire _63380 = _63375 ^ _63379;
  wire _63381 = uncoded_block[1581] ^ uncoded_block[1595];
  wire _63382 = _63381 ^ _14517;
  wire _63383 = _63382 ^ _22290;
  wire _63384 = uncoded_block[1617] ^ uncoded_block[1622];
  wire _63385 = _63384 ^ _22292;
  wire _63386 = _4667 ^ _62118;
  wire _63387 = _63385 ^ _63386;
  wire _63388 = _63383 ^ _63387;
  wire _63389 = _63380 ^ _63388;
  wire _63390 = _63371 ^ _63389;
  wire _63391 = _63355 ^ _63390;
  wire _63392 = _39465 ^ _6055;
  wire _63393 = uncoded_block[1674] ^ uncoded_block[1683];
  wire _63394 = _6058 ^ _63393;
  wire _63395 = _63392 ^ _63394;
  wire _63396 = uncoded_block[1687] ^ uncoded_block[1694];
  wire _63397 = _63396 ^ _9677;
  wire _63398 = _10778 ^ uncoded_block[1717];
  wire _63399 = _63397 ^ _63398;
  wire _63400 = _63395 ^ _63399;
  wire _63401 = _63391 ^ _63400;
  wire _63402 = _63316 ^ _63401;
  wire _63403 = uncoded_block[0] ^ uncoded_block[21];
  wire _63404 = _63403 ^ _18;
  wire _63405 = uncoded_block[51] ^ uncoded_block[65];
  wire _63406 = _56408 ^ _63405;
  wire _63407 = _63404 ^ _63406;
  wire _63408 = _42 ^ _44806;
  wire _63409 = _22806 ^ _63408;
  wire _63410 = _63407 ^ _63409;
  wire _63411 = _59257 ^ _59259;
  wire _63412 = uncoded_block[151] ^ uncoded_block[158];
  wire _63413 = uncoded_block[169] ^ uncoded_block[179];
  wire _63414 = _63412 ^ _63413;
  wire _63415 = _63411 ^ _63414;
  wire _63416 = _42607 ^ _2531;
  wire _63417 = _59265 ^ _50418;
  wire _63418 = _63416 ^ _63417;
  wire _63419 = _63415 ^ _63418;
  wire _63420 = _63410 ^ _63419;
  wire _63421 = uncoded_block[249] ^ uncoded_block[260];
  wire _63422 = _63421 ^ _56436;
  wire _63423 = _63422 ^ _56440;
  wire _63424 = uncoded_block[324] ^ uncoded_block[333];
  wire _63425 = _59270 ^ _63424;
  wire _63426 = _6859 ^ _10329;
  wire _63427 = _63425 ^ _63426;
  wire _63428 = _63423 ^ _63427;
  wire _63429 = uncoded_block[373] ^ uncoded_block[388];
  wire _63430 = _56450 ^ _63429;
  wire _63431 = uncoded_block[396] ^ uncoded_block[404];
  wire _63432 = uncoded_block[407] ^ uncoded_block[419];
  wire _63433 = _63431 ^ _63432;
  wire _63434 = _63430 ^ _63433;
  wire _63435 = uncoded_block[440] ^ uncoded_block[456];
  wire _63436 = _6894 ^ _63435;
  wire _63437 = uncoded_block[477] ^ uncoded_block[488];
  wire _63438 = _4185 ^ _63437;
  wire _63439 = _63436 ^ _63438;
  wire _63440 = _63434 ^ _63439;
  wire _63441 = _63428 ^ _63440;
  wire _63442 = _63420 ^ _63441;
  wire _63443 = _6919 ^ _18669;
  wire _63444 = _63443 ^ _59289;
  wire _63445 = uncoded_block[559] ^ uncoded_block[575];
  wire _63446 = _63445 ^ _26096;
  wire _63447 = _1938 ^ _56478;
  wire _63448 = _63446 ^ _63447;
  wire _63449 = _63444 ^ _63448;
  wire _63450 = _14218 ^ _15261;
  wire _63451 = _3502 ^ _22954;
  wire _63452 = _63450 ^ _63451;
  wire _63453 = _19674 ^ _15774;
  wire _63454 = uncoded_block[675] ^ uncoded_block[689];
  wire _63455 = uncoded_block[693] ^ uncoded_block[717];
  wire _63456 = _63454 ^ _63455;
  wire _63457 = _63453 ^ _63456;
  wire _63458 = _63452 ^ _63457;
  wire _63459 = _63449 ^ _63458;
  wire _63460 = uncoded_block[720] ^ uncoded_block[729];
  wire _63461 = _63460 ^ _9908;
  wire _63462 = uncoded_block[750] ^ uncoded_block[767];
  wire _63463 = _5013 ^ _63462;
  wire _63464 = _63461 ^ _63463;
  wire _63465 = uncoded_block[779] ^ uncoded_block[784];
  wire _63466 = _7617 ^ _63465;
  wire _63467 = _7026 ^ _59316;
  wire _63468 = _63466 ^ _63467;
  wire _63469 = _63464 ^ _63468;
  wire _63470 = uncoded_block[811] ^ uncoded_block[831];
  wire _63471 = uncoded_block[832] ^ uncoded_block[835];
  wire _63472 = _63470 ^ _63471;
  wire _63473 = uncoded_block[862] ^ uncoded_block[881];
  wire _63474 = _2814 ^ _63473;
  wire _63475 = _63472 ^ _63474;
  wire _63476 = uncoded_block[901] ^ uncoded_block[912];
  wire _63477 = _58838 ^ _63476;
  wire _63478 = _52872 ^ _25736;
  wire _63479 = _63477 ^ _63478;
  wire _63480 = _63475 ^ _63479;
  wire _63481 = _63469 ^ _63480;
  wire _63482 = _63459 ^ _63481;
  wire _63483 = _63442 ^ _63482;
  wire _63484 = _43454 ^ _12179;
  wire _63485 = uncoded_block[980] ^ uncoded_block[988];
  wire _63486 = _5786 ^ _63485;
  wire _63487 = _63484 ^ _63486;
  wire _63488 = _35704 ^ _5129;
  wire _63489 = _63488 ^ _59336;
  wire _63490 = _63487 ^ _63489;
  wire _63491 = _59337 ^ _56543;
  wire _63492 = _22145 ^ _6486;
  wire _63493 = _63491 ^ _63492;
  wire _63494 = uncoded_block[1080] ^ uncoded_block[1096];
  wire _63495 = _63494 ^ _19794;
  wire _63496 = _63495 ^ _56554;
  wire _63497 = _63493 ^ _63496;
  wire _63498 = _63490 ^ _63497;
  wire _63499 = _46389 ^ _14894;
  wire _63500 = uncoded_block[1187] ^ uncoded_block[1196];
  wire _63501 = _43127 ^ _63500;
  wire _63502 = _63499 ^ _63501;
  wire _63503 = _32484 ^ _21263;
  wire _63504 = _5218 ^ _15441;
  wire _63505 = _63503 ^ _63504;
  wire _63506 = _63502 ^ _63505;
  wire _63507 = uncoded_block[1279] ^ uncoded_block[1298];
  wire _63508 = _63507 ^ _18870;
  wire _63509 = _59359 ^ _63508;
  wire _63510 = _62421 ^ _34581;
  wire _63511 = _24951 ^ _11776;
  wire _63512 = _63510 ^ _63511;
  wire _63513 = _63509 ^ _63512;
  wire _63514 = _63506 ^ _63513;
  wire _63515 = _63498 ^ _63514;
  wire _63516 = uncoded_block[1372] ^ uncoded_block[1377];
  wire _63517 = uncoded_block[1391] ^ uncoded_block[1400];
  wire _63518 = _63516 ^ _63517;
  wire _63519 = uncoded_block[1414] ^ uncoded_block[1429];
  wire _63520 = _25406 ^ _63519;
  wire _63521 = _63518 ^ _63520;
  wire _63522 = uncoded_block[1438] ^ uncoded_block[1447];
  wire _63523 = _59615 ^ _63522;
  wire _63524 = _3865 ^ _6622;
  wire _63525 = _63523 ^ _63524;
  wire _63526 = _63521 ^ _63525;
  wire _63527 = _4601 ^ _3884;
  wire _63528 = _9042 ^ _1563;
  wire _63529 = _63527 ^ _63528;
  wire _63530 = uncoded_block[1498] ^ uncoded_block[1511];
  wire _63531 = _63530 ^ _15004;
  wire _63532 = _1582 ^ _24994;
  wire _63533 = _63531 ^ _63532;
  wire _63534 = _63529 ^ _63533;
  wire _63535 = _63526 ^ _63534;
  wire _63536 = uncoded_block[1566] ^ uncoded_block[1575];
  wire _63537 = _5347 ^ _63536;
  wire _63538 = _63537 ^ _59388;
  wire _63539 = uncoded_block[1599] ^ uncoded_block[1615];
  wire _63540 = uncoded_block[1625] ^ uncoded_block[1633];
  wire _63541 = _63539 ^ _63540;
  wire _63542 = uncoded_block[1643] ^ uncoded_block[1652];
  wire _63543 = _63542 ^ _53026;
  wire _63544 = _63541 ^ _63543;
  wire _63545 = _63538 ^ _63544;
  wire _63546 = _56628 ^ _2429;
  wire _63547 = _11327 ^ uncoded_block[1714];
  wire _63548 = _63546 ^ _63547;
  wire _63549 = _63545 ^ _63548;
  wire _63550 = _63535 ^ _63549;
  wire _63551 = _63515 ^ _63550;
  wire _63552 = _63483 ^ _63551;
  wire _63553 = uncoded_block[12] ^ uncoded_block[22];
  wire _63554 = _27241 ^ _63553;
  wire _63555 = _63554 ^ _58051;
  wire _63556 = _2475 ^ _6745;
  wire _63557 = uncoded_block[75] ^ uncoded_block[83];
  wire _63558 = uncoded_block[86] ^ uncoded_block[100];
  wire _63559 = _63557 ^ _63558;
  wire _63560 = _63556 ^ _63559;
  wire _63561 = _63555 ^ _63560;
  wire _63562 = uncoded_block[102] ^ uncoded_block[108];
  wire _63563 = uncoded_block[114] ^ uncoded_block[126];
  wire _63564 = _63562 ^ _63563;
  wire _63565 = _32634 ^ _22819;
  wire _63566 = _63564 ^ _63565;
  wire _63567 = uncoded_block[154] ^ uncoded_block[160];
  wire _63568 = _15620 ^ _63567;
  wire _63569 = uncoded_block[161] ^ uncoded_block[169];
  wire _63570 = uncoded_block[181] ^ uncoded_block[187];
  wire _63571 = _63569 ^ _63570;
  wire _63572 = _63568 ^ _63571;
  wire _63573 = _63566 ^ _63572;
  wire _63574 = _63561 ^ _63573;
  wire _63575 = uncoded_block[189] ^ uncoded_block[195];
  wire _63576 = _63575 ^ _25983;
  wire _63577 = _4070 ^ _35134;
  wire _63578 = _63576 ^ _63577;
  wire _63579 = _48830 ^ _8028;
  wire _63580 = uncoded_block[234] ^ uncoded_block[243];
  wire _63581 = _63580 ^ _16129;
  wire _63582 = _63579 ^ _63581;
  wire _63583 = _63578 ^ _63582;
  wire _63584 = uncoded_block[259] ^ uncoded_block[271];
  wire _63585 = _19061 ^ _63584;
  wire _63586 = _17142 ^ _3334;
  wire _63587 = _63585 ^ _63586;
  wire _63588 = _21942 ^ _11444;
  wire _63589 = _3352 ^ _10323;
  wire _63590 = _63588 ^ _63589;
  wire _63591 = _63587 ^ _63590;
  wire _63592 = _63583 ^ _63591;
  wire _63593 = _63574 ^ _63592;
  wire _63594 = uncoded_block[378] ^ uncoded_block[384];
  wire _63595 = _56700 ^ _63594;
  wire _63596 = _1045 ^ _1849;
  wire _63597 = _63595 ^ _63596;
  wire _63598 = _13646 ^ _184;
  wire _63599 = uncoded_block[410] ^ uncoded_block[425];
  wire _63600 = _63599 ^ _6894;
  wire _63601 = _63598 ^ _63600;
  wire _63602 = _63597 ^ _63601;
  wire _63603 = _39976 ^ _1866;
  wire _63604 = uncoded_block[454] ^ uncoded_block[466];
  wire _63605 = uncoded_block[479] ^ uncoded_block[488];
  wire _63606 = _63604 ^ _63605;
  wire _63607 = _63603 ^ _63606;
  wire _63608 = _10937 ^ _9294;
  wire _63609 = _1895 ^ _20603;
  wire _63610 = _63608 ^ _63609;
  wire _63611 = _63607 ^ _63610;
  wire _63612 = _63602 ^ _63611;
  wire _63613 = uncoded_block[534] ^ uncoded_block[542];
  wire _63614 = _63613 ^ _2687;
  wire _63615 = uncoded_block[564] ^ uncoded_block[572];
  wire _63616 = _15236 ^ _63615;
  wire _63617 = _63614 ^ _63616;
  wire _63618 = _263 ^ _24289;
  wire _63619 = uncoded_block[608] ^ uncoded_block[615];
  wire _63620 = _9330 ^ _63619;
  wire _63621 = _63618 ^ _63620;
  wire _63622 = _63617 ^ _63621;
  wire _63623 = uncoded_block[633] ^ uncoded_block[644];
  wire _63624 = _27797 ^ _63623;
  wire _63625 = _3514 ^ _7582;
  wire _63626 = _63624 ^ _63625;
  wire _63627 = _28158 ^ _1968;
  wire _63628 = uncoded_block[681] ^ uncoded_block[695];
  wire _63629 = _63628 ^ _333;
  wire _63630 = _63627 ^ _63629;
  wire _63631 = _63626 ^ _63630;
  wire _63632 = _63622 ^ _63631;
  wire _63633 = _63612 ^ _63632;
  wire _63634 = _63593 ^ _63633;
  wire _63635 = _24320 ^ _4998;
  wire _63636 = uncoded_block[719] ^ uncoded_block[725];
  wire _63637 = uncoded_block[729] ^ uncoded_block[737];
  wire _63638 = _63636 ^ _63637;
  wire _63639 = _63635 ^ _63638;
  wire _63640 = uncoded_block[763] ^ uncoded_block[772];
  wire _63641 = _12109 ^ _63640;
  wire _63642 = _41197 ^ _63641;
  wire _63643 = _63639 ^ _63642;
  wire _63644 = uncoded_block[773] ^ uncoded_block[785];
  wire _63645 = _63644 ^ _5032;
  wire _63646 = _26589 ^ _10486;
  wire _63647 = _63645 ^ _63646;
  wire _63648 = _48953 ^ _23003;
  wire _63649 = uncoded_block[846] ^ uncoded_block[856];
  wire _63650 = _38481 ^ _63649;
  wire _63651 = _63648 ^ _63650;
  wire _63652 = _63647 ^ _63651;
  wire _63653 = _63643 ^ _63652;
  wire _63654 = _6415 ^ _29803;
  wire _63655 = uncoded_block[890] ^ uncoded_block[904];
  wire _63656 = _1272 ^ _63655;
  wire _63657 = _63654 ^ _63656;
  wire _63658 = _23917 ^ _17820;
  wire _63659 = uncoded_block[932] ^ uncoded_block[942];
  wire _63660 = _63659 ^ _27476;
  wire _63661 = _63658 ^ _63660;
  wire _63662 = _63657 ^ _63661;
  wire _63663 = uncoded_block[961] ^ uncoded_block[969];
  wire _63664 = uncoded_block[972] ^ uncoded_block[980];
  wire _63665 = _63663 ^ _63664;
  wire _63666 = uncoded_block[982] ^ uncoded_block[1009];
  wire _63667 = _63666 ^ _13283;
  wire _63668 = _63665 ^ _63667;
  wire _63669 = uncoded_block[1018] ^ uncoded_block[1024];
  wire _63670 = _9996 ^ _63669;
  wire _63671 = uncoded_block[1056] ^ uncoded_block[1064];
  wire _63672 = _11677 ^ _63671;
  wire _63673 = _63670 ^ _63672;
  wire _63674 = _63668 ^ _63673;
  wire _63675 = _63662 ^ _63674;
  wire _63676 = _63653 ^ _63675;
  wire _63677 = uncoded_block[1069] ^ uncoded_block[1088];
  wire _63678 = _8889 ^ _63677;
  wire _63679 = uncoded_block[1092] ^ uncoded_block[1098];
  wire _63680 = uncoded_block[1104] ^ uncoded_block[1114];
  wire _63681 = _63679 ^ _63680;
  wire _63682 = _63678 ^ _63681;
  wire _63683 = _62076 ^ _20269;
  wire _63684 = _9502 ^ _15907;
  wire _63685 = _63683 ^ _63684;
  wire _63686 = _63682 ^ _63685;
  wire _63687 = _41296 ^ _44670;
  wire _63688 = _63687 ^ _27547;
  wire _63689 = uncoded_block[1211] ^ uncoded_block[1229];
  wire _63690 = _30346 ^ _63689;
  wire _63691 = uncoded_block[1243] ^ uncoded_block[1252];
  wire _63692 = uncoded_block[1254] ^ uncoded_block[1263];
  wire _63693 = _63691 ^ _63692;
  wire _63694 = _63690 ^ _63693;
  wire _63695 = _63688 ^ _63694;
  wire _63696 = _63686 ^ _63695;
  wire _63697 = uncoded_block[1272] ^ uncoded_block[1284];
  wire _63698 = _30363 ^ _63697;
  wire _63699 = uncoded_block[1285] ^ uncoded_block[1305];
  wire _63700 = uncoded_block[1308] ^ uncoded_block[1314];
  wire _63701 = _63699 ^ _63700;
  wire _63702 = _63698 ^ _63701;
  wire _63703 = uncoded_block[1329] ^ uncoded_block[1334];
  wire _63704 = _9555 ^ _63703;
  wire _63705 = uncoded_block[1344] ^ uncoded_block[1351];
  wire _63706 = _63705 ^ _673;
  wire _63707 = _63704 ^ _63706;
  wire _63708 = _63702 ^ _63707;
  wire _63709 = uncoded_block[1379] ^ uncoded_block[1384];
  wire _63710 = _46826 ^ _63709;
  wire _63711 = uncoded_block[1400] ^ uncoded_block[1405];
  wire _63712 = _20834 ^ _63711;
  wire _63713 = _63710 ^ _63712;
  wire _63714 = uncoded_block[1407] ^ uncoded_block[1418];
  wire _63715 = uncoded_block[1419] ^ uncoded_block[1432];
  wire _63716 = _63714 ^ _63715;
  wire _63717 = _10124 ^ _13432;
  wire _63718 = _63716 ^ _63717;
  wire _63719 = _63713 ^ _63718;
  wire _63720 = _63708 ^ _63719;
  wire _63721 = _63696 ^ _63720;
  wire _63722 = _63676 ^ _63721;
  wire _63723 = _63634 ^ _63722;
  wire _63724 = _8450 ^ _20852;
  wire _63725 = uncoded_block[1473] ^ uncoded_block[1486];
  wire _63726 = _8455 ^ _63725;
  wire _63727 = _63724 ^ _63726;
  wire _63728 = uncoded_block[1496] ^ uncoded_block[1503];
  wire _63729 = uncoded_block[1516] ^ uncoded_block[1532];
  wire _63730 = _63728 ^ _63729;
  wire _63731 = uncoded_block[1533] ^ uncoded_block[1540];
  wire _63732 = _63731 ^ _15020;
  wire _63733 = _63730 ^ _63732;
  wire _63734 = _63727 ^ _63733;
  wire _63735 = _22731 ^ _3141;
  wire _63736 = _15535 ^ _21821;
  wire _63737 = _63735 ^ _63736;
  wire _63738 = _11849 ^ _60726;
  wire _63739 = uncoded_block[1616] ^ uncoded_block[1628];
  wire _63740 = _63739 ^ _3948;
  wire _63741 = _63738 ^ _63740;
  wire _63742 = _63737 ^ _63741;
  wire _63743 = _63734 ^ _63742;
  wire _63744 = uncoded_block[1647] ^ uncoded_block[1653];
  wire _63745 = _815 ^ _63744;
  wire _63746 = uncoded_block[1658] ^ uncoded_block[1664];
  wire _63747 = _10760 ^ _63746;
  wire _63748 = _63745 ^ _63747;
  wire _63749 = _41412 ^ _830;
  wire _63750 = uncoded_block[1677] ^ uncoded_block[1684];
  wire _63751 = _63750 ^ _11324;
  wire _63752 = _63749 ^ _63751;
  wire _63753 = _63748 ^ _63752;
  wire _63754 = uncoded_block[1693] ^ uncoded_block[1700];
  wire _63755 = uncoded_block[1703] ^ uncoded_block[1707];
  wire _63756 = _63754 ^ _63755;
  wire _63757 = _30027 ^ uncoded_block[1718];
  wire _63758 = _63756 ^ _63757;
  wire _63759 = _63753 ^ _63758;
  wire _63760 = _63743 ^ _63759;
  wire _63761 = _63723 ^ _63760;
  wire _63762 = _3212 ^ _2454;
  wire _63763 = _46150 ^ _22790;
  wire _63764 = _63762 ^ _63763;
  wire _63765 = uncoded_block[37] ^ uncoded_block[51];
  wire _63766 = _22333 ^ _63765;
  wire _63767 = _63766 ^ _51115;
  wire _63768 = _63764 ^ _63767;
  wire _63769 = _1714 ^ _28438;
  wire _63770 = _42591 ^ _7981;
  wire _63771 = _63769 ^ _63770;
  wire _63772 = _20952 ^ _15101;
  wire _63773 = _63772 ^ _17089;
  wire _63774 = _63771 ^ _63773;
  wire _63775 = _63768 ^ _63774;
  wire _63776 = _25967 ^ _31392;
  wire _63777 = _33069 ^ _19539;
  wire _63778 = _63776 ^ _63777;
  wire _63779 = uncoded_block[179] ^ uncoded_block[189];
  wire _63780 = _63779 ^ _33077;
  wire _63781 = uncoded_block[198] ^ uncoded_block[208];
  wire _63782 = _63781 ^ _4071;
  wire _63783 = _63780 ^ _63782;
  wire _63784 = _63778 ^ _63783;
  wire _63785 = _10854 ^ _11945;
  wire _63786 = _63785 ^ _45193;
  wire _63787 = uncoded_block[240] ^ uncoded_block[247];
  wire _63788 = _63787 ^ _2556;
  wire _63789 = _33510 ^ _37959;
  wire _63790 = _63788 ^ _63789;
  wire _63791 = _63786 ^ _63790;
  wire _63792 = _63784 ^ _63791;
  wire _63793 = _63775 ^ _63792;
  wire _63794 = uncoded_block[272] ^ uncoded_block[279];
  wire _63795 = _63794 ^ _29238;
  wire _63796 = uncoded_block[295] ^ uncoded_block[305];
  wire _63797 = _4819 ^ _63796;
  wire _63798 = _63795 ^ _63797;
  wire _63799 = _21017 ^ _1813;
  wire _63800 = _11441 ^ _12521;
  wire _63801 = _63799 ^ _63800;
  wire _63802 = _63798 ^ _63801;
  wire _63803 = _38366 ^ _54294;
  wire _63804 = _17650 ^ _63803;
  wire _63805 = uncoded_block[371] ^ uncoded_block[378];
  wire _63806 = _63805 ^ _6876;
  wire _63807 = uncoded_block[394] ^ uncoded_block[412];
  wire _63808 = _10907 ^ _63807;
  wire _63809 = _63806 ^ _63808;
  wire _63810 = _63804 ^ _63809;
  wire _63811 = _63802 ^ _63810;
  wire _63812 = uncoded_block[418] ^ uncoded_block[426];
  wire _63813 = _5565 ^ _63812;
  wire _63814 = _14687 ^ _16187;
  wire _63815 = _63813 ^ _63814;
  wire _63816 = _17181 ^ _7498;
  wire _63817 = uncoded_block[451] ^ uncoded_block[457];
  wire _63818 = _63817 ^ _10926;
  wire _63819 = _63816 ^ _63818;
  wire _63820 = _63815 ^ _63819;
  wire _63821 = uncoded_block[471] ^ uncoded_block[482];
  wire _63822 = _63821 ^ _9291;
  wire _63823 = _20081 ^ _63822;
  wire _63824 = _30167 ^ _1892;
  wire _63825 = uncoded_block[511] ^ uncoded_block[515];
  wire _63826 = uncoded_block[516] ^ uncoded_block[525];
  wire _63827 = _63825 ^ _63826;
  wire _63828 = _63824 ^ _63827;
  wire _63829 = _63823 ^ _63828;
  wire _63830 = _63820 ^ _63829;
  wire _63831 = _63811 ^ _63830;
  wire _63832 = _63793 ^ _63831;
  wire _63833 = _6292 ^ _28882;
  wire _63834 = _1118 ^ _48152;
  wire _63835 = _63833 ^ _63834;
  wire _63836 = _20110 ^ _4941;
  wire _63837 = _10400 ^ _4946;
  wire _63838 = _63836 ^ _63837;
  wire _63839 = _63835 ^ _63838;
  wire _63840 = uncoded_block[586] ^ uncoded_block[593];
  wire _63841 = _63840 ^ _7558;
  wire _63842 = uncoded_block[603] ^ uncoded_block[615];
  wire _63843 = _63842 ^ _15261;
  wire _63844 = _63841 ^ _63843;
  wire _63845 = _3502 ^ _50498;
  wire _63846 = _8755 ^ _2739;
  wire _63847 = _63845 ^ _63846;
  wire _63848 = _63844 ^ _63847;
  wire _63849 = _63839 ^ _63848;
  wire _63850 = _309 ^ _40427;
  wire _63851 = _6983 ^ _17753;
  wire _63852 = _63850 ^ _63851;
  wire _63853 = uncoded_block[697] ^ uncoded_block[709];
  wire _63854 = _63853 ^ _2762;
  wire _63855 = _2763 ^ _5691;
  wire _63856 = _63854 ^ _63855;
  wire _63857 = _63852 ^ _63856;
  wire _63858 = _59509 ^ _11576;
  wire _63859 = uncoded_block[754] ^ uncoded_block[764];
  wire _63860 = _8209 ^ _63859;
  wire _63861 = _63858 ^ _63860;
  wire _63862 = _13215 ^ _39661;
  wire _63863 = uncoded_block[791] ^ uncoded_block[798];
  wire _63864 = _49309 ^ _63863;
  wire _63865 = _63862 ^ _63864;
  wire _63866 = _63861 ^ _63865;
  wire _63867 = _63857 ^ _63866;
  wire _63868 = _63849 ^ _63867;
  wire _63869 = _35268 ^ _6398;
  wire _63870 = _397 ^ _53188;
  wire _63871 = _63869 ^ _63870;
  wire _63872 = _3599 ^ _6406;
  wire _63873 = _46322 ^ _63872;
  wire _63874 = _63871 ^ _63873;
  wire _63875 = uncoded_block[855] ^ uncoded_block[871];
  wire _63876 = _63875 ^ _6416;
  wire _63877 = uncoded_block[877] ^ uncoded_block[891];
  wire _63878 = _63877 ^ _12704;
  wire _63879 = _63876 ^ _63878;
  wire _63880 = uncoded_block[894] ^ uncoded_block[898];
  wire _63881 = uncoded_block[902] ^ uncoded_block[913];
  wire _63882 = _63880 ^ _63881;
  wire _63883 = _8256 ^ _25736;
  wire _63884 = _63882 ^ _63883;
  wire _63885 = _63879 ^ _63884;
  wire _63886 = _63874 ^ _63885;
  wire _63887 = _32828 ^ _51310;
  wire _63888 = uncoded_block[958] ^ uncoded_block[966];
  wire _63889 = _4382 ^ _63888;
  wire _63890 = _4390 ^ _29832;
  wire _63891 = _63889 ^ _63890;
  wire _63892 = _63887 ^ _63891;
  wire _63893 = _5798 ^ _4404;
  wire _63894 = _8866 ^ _9993;
  wire _63895 = _63893 ^ _63894;
  wire _63896 = _492 ^ _498;
  wire _63897 = _4418 ^ _16864;
  wire _63898 = _63896 ^ _63897;
  wire _63899 = _63895 ^ _63898;
  wire _63900 = _63892 ^ _63899;
  wire _63901 = _63886 ^ _63900;
  wire _63902 = _63868 ^ _63901;
  wire _63903 = _63832 ^ _63902;
  wire _63904 = _2913 ^ _14355;
  wire _63905 = _522 ^ _13851;
  wire _63906 = _63904 ^ _63905;
  wire _63907 = _2147 ^ _19301;
  wire _63908 = uncoded_block[1093] ^ uncoded_block[1099];
  wire _63909 = _10021 ^ _63908;
  wire _63910 = _63907 ^ _63909;
  wire _63911 = _63906 ^ _63910;
  wire _63912 = uncoded_block[1100] ^ uncoded_block[1123];
  wire _63913 = _63912 ^ _5178;
  wire _63914 = _63913 ^ _48274;
  wire _63915 = uncoded_block[1161] ^ uncoded_block[1168];
  wire _63916 = _578 ^ _63915;
  wire _63917 = _63916 ^ _43886;
  wire _63918 = _63914 ^ _63917;
  wire _63919 = _63911 ^ _63918;
  wire _63920 = uncoded_block[1182] ^ uncoded_block[1187];
  wire _63921 = _63920 ^ _40904;
  wire _63922 = uncoded_block[1213] ^ uncoded_block[1217];
  wire _63923 = _14912 ^ _63922;
  wire _63924 = _63921 ^ _63923;
  wire _63925 = _4499 ^ _55360;
  wire _63926 = uncoded_block[1256] ^ uncoded_block[1260];
  wire _63927 = _31231 ^ _63926;
  wire _63928 = _63925 ^ _63927;
  wire _63929 = _63924 ^ _63928;
  wire _63930 = uncoded_block[1271] ^ uncoded_block[1280];
  wire _63931 = _4516 ^ _63930;
  wire _63932 = _4525 ^ _29913;
  wire _63933 = _63931 ^ _63932;
  wire _63934 = uncoded_block[1310] ^ uncoded_block[1324];
  wire _63935 = _23131 ^ _63934;
  wire _63936 = _42101 ^ _63935;
  wire _63937 = _63933 ^ _63936;
  wire _63938 = _63929 ^ _63937;
  wire _63939 = _63919 ^ _63938;
  wire _63940 = _15467 ^ _661;
  wire _63941 = _55382 ^ _672;
  wire _63942 = _63940 ^ _63941;
  wire _63943 = _54880 ^ _3054;
  wire _63944 = uncoded_block[1381] ^ uncoded_block[1396];
  wire _63945 = _63944 ^ _695;
  wire _63946 = _63943 ^ _63945;
  wire _63947 = _63942 ^ _63946;
  wire _63948 = uncoded_block[1410] ^ uncoded_block[1417];
  wire _63949 = _63948 ^ _1526;
  wire _63950 = uncoded_block[1441] ^ uncoded_block[1449];
  wire _63951 = _13951 ^ _63950;
  wire _63952 = _63949 ^ _63951;
  wire _63953 = uncoded_block[1453] ^ uncoded_block[1461];
  wire _63954 = _63953 ^ _20362;
  wire _63955 = uncoded_block[1472] ^ uncoded_block[1481];
  wire _63956 = _18919 ^ _63955;
  wire _63957 = _63954 ^ _63956;
  wire _63958 = _63952 ^ _63957;
  wire _63959 = _63947 ^ _63958;
  wire _63960 = uncoded_block[1507] ^ uncoded_block[1516];
  wire _63961 = _7861 ^ _63960;
  wire _63962 = _9624 ^ _46860;
  wire _63963 = _63961 ^ _63962;
  wire _63964 = uncoded_block[1542] ^ uncoded_block[1546];
  wire _63965 = _36656 ^ _63964;
  wire _63966 = uncoded_block[1555] ^ uncoded_block[1562];
  wire _63967 = _29977 ^ _63966;
  wire _63968 = _63965 ^ _63967;
  wire _63969 = _63963 ^ _63968;
  wire _63970 = _16019 ^ _7891;
  wire _63971 = uncoded_block[1580] ^ uncoded_block[1588];
  wire _63972 = _63971 ^ _791;
  wire _63973 = _63970 ^ _63972;
  wire _63974 = uncoded_block[1594] ^ uncoded_block[1599];
  wire _63975 = uncoded_block[1611] ^ uncoded_block[1616];
  wire _63976 = _63974 ^ _63975;
  wire _63977 = _63976 ^ _42174;
  wire _63978 = _63973 ^ _63977;
  wire _63979 = _63969 ^ _63978;
  wire _63980 = _63959 ^ _63979;
  wire _63981 = _63939 ^ _63980;
  wire _63982 = uncoded_block[1629] ^ uncoded_block[1640];
  wire _63983 = _14525 ^ _63982;
  wire _63984 = _63983 ^ _52332;
  wire _63985 = uncoded_block[1660] ^ uncoded_block[1671];
  wire _63986 = _63985 ^ _37094;
  wire _63987 = _20418 ^ _63986;
  wire _63988 = _63984 ^ _63987;
  wire _63989 = uncoded_block[1681] ^ uncoded_block[1690];
  wire _63990 = _63989 ^ _11327;
  wire _63991 = uncoded_block[1708] ^ uncoded_block[1720];
  wire _63992 = _63991 ^ uncoded_block[1721];
  wire _63993 = _63990 ^ _63992;
  wire _63994 = _63988 ^ _63993;
  wire _63995 = _63981 ^ _63994;
  wire _63996 = _63903 ^ _63995;
  wire _63997 = uncoded_block[7] ^ uncoded_block[14];
  wire _63998 = uncoded_block[16] ^ uncoded_block[27];
  wire _63999 = _63997 ^ _63998;
  wire _64000 = _15594 ^ _48418;
  wire _64001 = _63999 ^ _64000;
  wire _64002 = _58054 ^ _12438;
  wire _64003 = uncoded_block[98] ^ uncoded_block[116];
  wire _64004 = _7374 ^ _64003;
  wire _64005 = _64002 ^ _64004;
  wire _64006 = _64001 ^ _64005;
  wire _64007 = uncoded_block[124] ^ uncoded_block[132];
  wire _64008 = _13571 ^ _64007;
  wire _64009 = uncoded_block[137] ^ uncoded_block[148];
  wire _64010 = uncoded_block[149] ^ uncoded_block[174];
  wire _64011 = _64009 ^ _64010;
  wire _64012 = _64008 ^ _64011;
  wire _64013 = uncoded_block[199] ^ uncoded_block[205];
  wire _64014 = _49664 ^ _64013;
  wire _64015 = uncoded_block[213] ^ uncoded_block[225];
  wire _64016 = _98 ^ _64015;
  wire _64017 = _64014 ^ _64016;
  wire _64018 = _64012 ^ _64017;
  wire _64019 = _64006 ^ _64018;
  wire _64020 = uncoded_block[233] ^ uncoded_block[242];
  wire _64021 = uncoded_block[248] ^ uncoded_block[256];
  wire _64022 = _64020 ^ _64021;
  wire _64023 = uncoded_block[270] ^ uncoded_block[281];
  wire _64024 = _64023 ^ _49687;
  wire _64025 = _64022 ^ _64024;
  wire _64026 = uncoded_block[292] ^ uncoded_block[305];
  wire _64027 = _64026 ^ _149;
  wire _64028 = _59955 ^ _38366;
  wire _64029 = _64027 ^ _64028;
  wire _64030 = _64025 ^ _64029;
  wire _64031 = uncoded_block[382] ^ uncoded_block[392];
  wire _64032 = _39567 ^ _64031;
  wire _64033 = uncoded_block[395] ^ uncoded_block[412];
  wire _64034 = _64033 ^ _3397;
  wire _64035 = _64032 ^ _64034;
  wire _64036 = uncoded_block[440] ^ uncoded_block[476];
  wire _64037 = uncoded_block[483] ^ uncoded_block[488];
  wire _64038 = _64036 ^ _64037;
  wire _64039 = _64038 ^ _17202;
  wire _64040 = _64035 ^ _64039;
  wire _64041 = _64030 ^ _64040;
  wire _64042 = _64019 ^ _64041;
  wire _64043 = uncoded_block[503] ^ uncoded_block[512];
  wire _64044 = _64043 ^ _17702;
  wire _64045 = uncoded_block[537] ^ uncoded_block[572];
  wire _64046 = _1108 ^ _64045;
  wire _64047 = _64044 ^ _64046;
  wire _64048 = uncoded_block[577] ^ uncoded_block[583];
  wire _64049 = _4941 ^ _64048;
  wire _64050 = uncoded_block[600] ^ uncoded_block[613];
  wire _64051 = _64050 ^ _2720;
  wire _64052 = _64049 ^ _64051;
  wire _64053 = _64047 ^ _64052;
  wire _64054 = uncoded_block[635] ^ uncoded_block[650];
  wire _64055 = _64054 ^ _302;
  wire _64056 = _309 ^ _4265;
  wire _64057 = _64055 ^ _64056;
  wire _64058 = _8761 ^ _4984;
  wire _64059 = _18721 ^ _21596;
  wire _64060 = _64058 ^ _64059;
  wire _64061 = _64057 ^ _64060;
  wire _64062 = _64053 ^ _64061;
  wire _64063 = _14264 ^ _12663;
  wire _64064 = _51267 ^ _3567;
  wire _64065 = _64063 ^ _64064;
  wire _64066 = uncoded_block[788] ^ uncoded_block[796];
  wire _64067 = _4309 ^ _64066;
  wire _64068 = uncoded_block[801] ^ uncoded_block[822];
  wire _64069 = _64068 ^ _10490;
  wire _64070 = _64067 ^ _64069;
  wire _64071 = _64065 ^ _64070;
  wire _64072 = uncoded_block[852] ^ uncoded_block[858];
  wire _64073 = _4336 ^ _64072;
  wire _64074 = uncoded_block[871] ^ uncoded_block[878];
  wire _64075 = _64074 ^ _21172;
  wire _64076 = _64073 ^ _64075;
  wire _64077 = uncoded_block[896] ^ uncoded_block[908];
  wire _64078 = _64077 ^ _63285;
  wire _64079 = uncoded_block[940] ^ uncoded_block[948];
  wire _64080 = _2083 ^ _64079;
  wire _64081 = _64078 ^ _64080;
  wire _64082 = _64076 ^ _64081;
  wire _64083 = _64071 ^ _64082;
  wire _64084 = _64062 ^ _64083;
  wire _64085 = _64042 ^ _64084;
  wire _64086 = uncoded_block[959] ^ uncoded_block[976];
  wire _64087 = _7083 ^ _64086;
  wire _64088 = uncoded_block[999] ^ uncoded_block[1007];
  wire _64089 = _2100 ^ _64088;
  wire _64090 = _64087 ^ _64089;
  wire _64091 = uncoded_block[1012] ^ uncoded_block[1028];
  wire _64092 = _64091 ^ _21218;
  wire _64093 = uncoded_block[1048] ^ uncoded_block[1060];
  wire _64094 = _12208 ^ _64093;
  wire _64095 = _64092 ^ _64094;
  wire _64096 = _64090 ^ _64095;
  wire _64097 = _8889 ^ _23505;
  wire _64098 = uncoded_block[1111] ^ uncoded_block[1121];
  wire _64099 = _5166 ^ _64098;
  wire _64100 = _64097 ^ _64099;
  wire _64101 = _8933 ^ _11711;
  wire _64102 = uncoded_block[1171] ^ uncoded_block[1183];
  wire _64103 = _5869 ^ _64102;
  wire _64104 = _64101 ^ _64103;
  wire _64105 = _64100 ^ _64104;
  wire _64106 = _64096 ^ _64105;
  wire _64107 = uncoded_block[1186] ^ uncoded_block[1202];
  wire _64108 = uncoded_block[1227] ^ uncoded_block[1239];
  wire _64109 = _64107 ^ _64108;
  wire _64110 = _17911 ^ _60875;
  wire _64111 = _64109 ^ _64110;
  wire _64112 = uncoded_block[1279] ^ uncoded_block[1289];
  wire _64113 = _64112 ^ _3017;
  wire _64114 = _17435 ^ _60071;
  wire _64115 = _64113 ^ _64114;
  wire _64116 = _64111 ^ _64115;
  wire _64117 = uncoded_block[1350] ^ uncoded_block[1356];
  wire _64118 = _63345 ^ _64117;
  wire _64119 = _64118 ^ _24043;
  wire _64120 = _61219 ^ _2299;
  wire _64121 = _13422 ^ _29508;
  wire _64122 = _64120 ^ _64121;
  wire _64123 = _64119 ^ _64122;
  wire _64124 = _64116 ^ _64123;
  wire _64125 = _64106 ^ _64124;
  wire _64126 = uncoded_block[1446] ^ uncoded_block[1462];
  wire _64127 = _64126 ^ _11255;
  wire _64128 = uncoded_block[1480] ^ uncoded_block[1500];
  wire _64129 = _64128 ^ _23624;
  wire _64130 = _64127 ^ _64129;
  wire _64131 = _7264 ^ _6643;
  wire _64132 = uncoded_block[1525] ^ uncoded_block[1531];
  wire _64133 = _5999 ^ _64132;
  wire _64134 = _64131 ^ _64133;
  wire _64135 = _64130 ^ _64134;
  wire _64136 = _38240 ^ _58311;
  wire _64137 = uncoded_block[1579] ^ uncoded_block[1587];
  wire _64138 = _64137 ^ _11295;
  wire _64139 = _64136 ^ _64138;
  wire _64140 = uncoded_block[1617] ^ uncoded_block[1625];
  wire _64141 = _4660 ^ _64140;
  wire _64142 = uncoded_block[1633] ^ uncoded_block[1640];
  wire _64143 = _64142 ^ _5399;
  wire _64144 = _64141 ^ _64143;
  wire _64145 = _64139 ^ _64144;
  wire _64146 = _64135 ^ _64145;
  wire _64147 = _7323 ^ _63754;
  wire _64148 = uncoded_block[1713] ^ uncoded_block[1718];
  wire _64149 = _851 ^ _64148;
  wire _64150 = _64147 ^ _64149;
  wire _64151 = _64150 ^ uncoded_block[1721];
  wire _64152 = _64146 ^ _64151;
  wire _64153 = _64125 ^ _64152;
  wire _64154 = _64085 ^ _64153;
  wire _64155 = _57589 ^ _9139;
  wire _64156 = _13543 ^ _3230;
  wire _64157 = _64155 ^ _64156;
  wire _64158 = uncoded_block[42] ^ uncoded_block[60];
  wire _64159 = _64158 ^ _11363;
  wire _64160 = _13558 ^ _56649;
  wire _64161 = _64159 ^ _64160;
  wire _64162 = _64157 ^ _64161;
  wire _64163 = uncoded_block[117] ^ uncoded_block[121];
  wire _64164 = _57601 ^ _64163;
  wire _64165 = uncoded_block[126] ^ uncoded_block[130];
  wire _64166 = uncoded_block[139] ^ uncoded_block[149];
  wire _64167 = _64165 ^ _64166;
  wire _64168 = _64164 ^ _64167;
  wire _64169 = uncoded_block[164] ^ uncoded_block[171];
  wire _64170 = _19040 ^ _64169;
  wire _64171 = _64170 ^ _57613;
  wire _64172 = _64168 ^ _64171;
  wire _64173 = _64162 ^ _64172;
  wire _64174 = uncoded_block[205] ^ uncoded_block[216];
  wire _64175 = _57614 ^ _64174;
  wire _64176 = _105 ^ _30087;
  wire _64177 = _64175 ^ _64176;
  wire _64178 = uncoded_block[240] ^ uncoded_block[250];
  wire _64179 = _64178 ^ _63584;
  wire _64180 = _2568 ^ _12506;
  wire _64181 = _64179 ^ _64180;
  wire _64182 = _64177 ^ _64181;
  wire _64183 = uncoded_block[302] ^ uncoded_block[325];
  wire _64184 = _138 ^ _64183;
  wire _64185 = _57625 ^ _64184;
  wire _64186 = _57630 ^ _11987;
  wire _64187 = _4844 ^ _20056;
  wire _64188 = _64186 ^ _64187;
  wire _64189 = _64185 ^ _64188;
  wire _64190 = _64182 ^ _64189;
  wire _64191 = _64173 ^ _64190;
  wire _64192 = uncoded_block[380] ^ uncoded_block[388];
  wire _64193 = _64192 ^ _10908;
  wire _64194 = uncoded_block[395] ^ uncoded_block[407];
  wire _64195 = uncoded_block[413] ^ uncoded_block[426];
  wire _64196 = _64194 ^ _64195;
  wire _64197 = _64193 ^ _64196;
  wire _64198 = _14690 ^ _14169;
  wire _64199 = uncoded_block[446] ^ uncoded_block[467];
  wire _64200 = _64199 ^ _6266;
  wire _64201 = _64198 ^ _64200;
  wire _64202 = _64197 ^ _64201;
  wire _64203 = uncoded_block[496] ^ uncoded_block[503];
  wire _64204 = _64203 ^ _14707;
  wire _64205 = _27767 ^ _64204;
  wire _64206 = uncoded_block[520] ^ uncoded_block[535];
  wire _64207 = _57045 ^ _64206;
  wire _64208 = _64207 ^ _57658;
  wire _64209 = _64205 ^ _64208;
  wire _64210 = _64202 ^ _64209;
  wire _64211 = uncoded_block[559] ^ uncoded_block[567];
  wire _64212 = _8724 ^ _64211;
  wire _64213 = _57661 ^ _277;
  wire _64214 = _64212 ^ _64213;
  wire _64215 = uncoded_block[621] ^ uncoded_block[629];
  wire _64216 = _14223 ^ _64215;
  wire _64217 = uncoded_block[638] ^ uncoded_block[647];
  wire _64218 = _57666 ^ _64217;
  wire _64219 = _64216 ^ _64218;
  wire _64220 = _64214 ^ _64219;
  wire _64221 = _297 ^ _3514;
  wire _64222 = _38439 ^ _8760;
  wire _64223 = _64221 ^ _64222;
  wire _64224 = _23863 ^ _2765;
  wire _64225 = _57678 ^ _64224;
  wire _64226 = _64223 ^ _64225;
  wire _64227 = _64220 ^ _64226;
  wire _64228 = _64210 ^ _64227;
  wire _64229 = _64191 ^ _64228;
  wire _64230 = _8204 ^ _13208;
  wire _64231 = uncoded_block[748] ^ uncoded_block[758];
  wire _64232 = _64231 ^ _49305;
  wire _64233 = _64230 ^ _64232;
  wire _64234 = _30234 ^ _57090;
  wire _64235 = _57684 ^ _31551;
  wire _64236 = _64234 ^ _64235;
  wire _64237 = _64233 ^ _64236;
  wire _64238 = uncoded_block[814] ^ uncoded_block[825];
  wire _64239 = _16791 ^ _64238;
  wire _64240 = uncoded_block[827] ^ uncoded_block[841];
  wire _64241 = _64240 ^ _14812;
  wire _64242 = _64239 ^ _64241;
  wire _64243 = _57695 ^ _57698;
  wire _64244 = _64242 ^ _64243;
  wire _64245 = _64237 ^ _64244;
  wire _64246 = _7665 ^ _8259;
  wire _64247 = _57699 ^ _64246;
  wire _64248 = uncoded_block[929] ^ uncoded_block[944];
  wire _64249 = uncoded_block[961] ^ uncoded_block[965];
  wire _64250 = _64248 ^ _64249;
  wire _64251 = _5785 ^ _468;
  wire _64252 = _64250 ^ _64251;
  wire _64253 = _64247 ^ _64252;
  wire _64254 = _3657 ^ _23939;
  wire _64255 = _59127 ^ _27077;
  wire _64256 = _64254 ^ _64255;
  wire _64257 = uncoded_block[1013] ^ uncoded_block[1050];
  wire _64258 = _64257 ^ _7717;
  wire _64259 = uncoded_block[1065] ^ uncoded_block[1076];
  wire _64260 = uncoded_block[1079] ^ uncoded_block[1085];
  wire _64261 = _64259 ^ _64260;
  wire _64262 = _64258 ^ _64261;
  wire _64263 = _64256 ^ _64262;
  wire _64264 = _64253 ^ _64263;
  wire _64265 = _64245 ^ _64264;
  wire _64266 = uncoded_block[1146] ^ uncoded_block[1154];
  wire _64267 = _10593 ^ _64266;
  wire _64268 = _64267 ^ _57727;
  wire _64269 = _57724 ^ _64268;
  wire _64270 = _11171 ^ _27911;
  wire _64271 = _12815 ^ _17907;
  wire _64272 = _64270 ^ _64271;
  wire _64273 = _57735 ^ _64272;
  wire _64274 = _64269 ^ _64273;
  wire _64275 = uncoded_block[1237] ^ uncoded_block[1250];
  wire _64276 = _64275 ^ _3780;
  wire _64277 = _64276 ^ _38581;
  wire _64278 = _1458 ^ _2247;
  wire _64279 = uncoded_block[1279] ^ uncoded_block[1287];
  wire _64280 = uncoded_block[1288] ^ uncoded_block[1293];
  wire _64281 = _64279 ^ _64280;
  wire _64282 = _64278 ^ _64281;
  wire _64283 = _64277 ^ _64282;
  wire _64284 = _35380 ^ _4539;
  wire _64285 = uncoded_block[1334] ^ uncoded_block[1340];
  wire _64286 = _59852 ^ _64285;
  wire _64287 = _64284 ^ _64286;
  wire _64288 = _29486 ^ _4564;
  wire _64289 = _25399 ^ _38613;
  wire _64290 = _64288 ^ _64289;
  wire _64291 = _64287 ^ _64290;
  wire _64292 = _64283 ^ _64291;
  wire _64293 = _64274 ^ _64292;
  wire _64294 = _64265 ^ _64293;
  wire _64295 = _64229 ^ _64294;
  wire _64296 = uncoded_block[1399] ^ uncoded_block[1408];
  wire _64297 = uncoded_block[1411] ^ uncoded_block[1425];
  wire _64298 = _64296 ^ _64297;
  wire _64299 = uncoded_block[1452] ^ uncoded_block[1467];
  wire _64300 = _17470 ^ _64299;
  wire _64301 = _64298 ^ _64300;
  wire _64302 = uncoded_block[1468] ^ uncoded_block[1495];
  wire _64303 = uncoded_block[1496] ^ uncoded_block[1504];
  wire _64304 = _64302 ^ _64303;
  wire _64305 = uncoded_block[1505] ^ uncoded_block[1515];
  wire _64306 = _64305 ^ _56921;
  wire _64307 = _64304 ^ _64306;
  wire _64308 = _64301 ^ _64307;
  wire _64309 = _38240 ^ _32975;
  wire _64310 = _4634 ^ _10724;
  wire _64311 = _64309 ^ _64310;
  wire _64312 = _10161 ^ _57779;
  wire _64313 = _64312 ^ _47246;
  wire _64314 = _64311 ^ _64313;
  wire _64315 = _64308 ^ _64314;
  wire _64316 = _25454 ^ _5373;
  wire _64317 = _6677 ^ _63975;
  wire _64318 = _64316 ^ _64317;
  wire _64319 = _38668 ^ _4667;
  wire _64320 = _57790 ^ _32178;
  wire _64321 = _64319 ^ _64320;
  wire _64322 = _64318 ^ _64321;
  wire _64323 = uncoded_block[1672] ^ uncoded_block[1680];
  wire _64324 = _64323 ^ _7933;
  wire _64325 = uncoded_block[1688] ^ uncoded_block[1708];
  wire _64326 = uncoded_block[1709] ^ uncoded_block[1715];
  wire _64327 = _64325 ^ _64326;
  wire _64328 = _64324 ^ _64327;
  wire _64329 = _64328 ^ _5416;
  wire _64330 = _64322 ^ _64329;
  wire _64331 = _64315 ^ _64330;
  wire _64332 = _64295 ^ _64331;
  wire _64333 = _14565 ^ _14048;
  wire _64334 = _14055 ^ _2480;
  wire _64335 = _64333 ^ _64334;
  wire _64336 = uncoded_block[76] ^ uncoded_block[105];
  wire _64337 = _64336 ^ _4034;
  wire _64338 = uncoded_block[134] ^ uncoded_block[162];
  wire _64339 = _64338 ^ _58738;
  wire _64340 = _64337 ^ _64339;
  wire _64341 = _64335 ^ _64340;
  wire _64342 = uncoded_block[199] ^ uncoded_block[208];
  wire _64343 = _64342 ^ _10854;
  wire _64344 = uncoded_block[234] ^ uncoded_block[252];
  wire _64345 = _33504 ^ _64344;
  wire _64346 = _64343 ^ _64345;
  wire _64347 = uncoded_block[254] ^ uncoded_block[269];
  wire _64348 = uncoded_block[284] ^ uncoded_block[289];
  wire _64349 = _64347 ^ _64348;
  wire _64350 = uncoded_block[316] ^ uncoded_block[328];
  wire _64351 = _15163 ^ _64350;
  wire _64352 = _64349 ^ _64351;
  wire _64353 = _64346 ^ _64352;
  wire _64354 = _64341 ^ _64353;
  wire _64355 = uncoded_block[352] ^ uncoded_block[379];
  wire _64356 = _7463 ^ _64355;
  wire _64357 = uncoded_block[383] ^ uncoded_block[390];
  wire _64358 = _64357 ^ _3394;
  wire _64359 = _64356 ^ _64358;
  wire _64360 = uncoded_block[415] ^ uncoded_block[426];
  wire _64361 = _64360 ^ _23349;
  wire _64362 = uncoded_block[449] ^ uncoded_block[460];
  wire _64363 = uncoded_block[469] ^ uncoded_block[484];
  wire _64364 = _64362 ^ _64363;
  wire _64365 = _64361 ^ _64364;
  wire _64366 = _64359 ^ _64365;
  wire _64367 = _228 ^ _10948;
  wire _64368 = uncoded_block[531] ^ uncoded_block[543];
  wire _64369 = _64368 ^ _5628;
  wire _64370 = _64367 ^ _64369;
  wire _64371 = uncoded_block[579] ^ uncoded_block[599];
  wire _64372 = _1130 ^ _64371;
  wire _64373 = uncoded_block[618] ^ uncoded_block[657];
  wire _64374 = _30624 ^ _64373;
  wire _64375 = _64372 ^ _64374;
  wire _64376 = _64370 ^ _64375;
  wire _64377 = _64366 ^ _64376;
  wire _64378 = _64354 ^ _64377;
  wire _64379 = _10440 ^ _9895;
  wire _64380 = uncoded_block[696] ^ uncoded_block[718];
  wire _64381 = _64380 ^ _32779;
  wire _64382 = _64379 ^ _64381;
  wire _64383 = uncoded_block[739] ^ uncoded_block[745];
  wire _64384 = _64383 ^ _4311;
  wire _64385 = uncoded_block[796] ^ uncoded_block[814];
  wire _64386 = _64385 ^ _60834;
  wire _64387 = _64384 ^ _64386;
  wire _64388 = _64382 ^ _64387;
  wire _64389 = uncoded_block[859] ^ uncoded_block[875];
  wire _64390 = _64389 ^ _8820;
  wire _64391 = uncoded_block[917] ^ uncoded_block[932];
  wire _64392 = _60999 ^ _64391;
  wire _64393 = _64390 ^ _64392;
  wire _64394 = _2083 ^ _11643;
  wire _64395 = uncoded_block[965] ^ uncoded_block[977];
  wire _64396 = _64395 ^ _47871;
  wire _64397 = _64394 ^ _64396;
  wire _64398 = _64393 ^ _64397;
  wire _64399 = _64388 ^ _64398;
  wire _64400 = uncoded_block[1011] ^ uncoded_block[1022];
  wire _64401 = uncoded_block[1031] ^ uncoded_block[1042];
  wire _64402 = _64400 ^ _64401;
  wire _64403 = uncoded_block[1062] ^ uncoded_block[1072];
  wire _64404 = _23966 ^ _64403;
  wire _64405 = _64402 ^ _64404;
  wire _64406 = uncoded_block[1077] ^ uncoded_block[1102];
  wire _64407 = uncoded_block[1121] ^ uncoded_block[1126];
  wire _64408 = _64406 ^ _64407;
  wire _64409 = uncoded_block[1146] ^ uncoded_block[1169];
  wire _64410 = _56555 ^ _64409;
  wire _64411 = _64408 ^ _64410;
  wire _64412 = _64405 ^ _64411;
  wire _64413 = _60866 ^ _11722;
  wire _64414 = uncoded_block[1253] ^ uncoded_block[1258];
  wire _64415 = _5901 ^ _64414;
  wire _64416 = _64413 ^ _64415;
  wire _64417 = uncoded_block[1297] ^ uncoded_block[1317];
  wire _64418 = _64417 ^ _48319;
  wire _64419 = _11207 ^ _2276;
  wire _64420 = _64418 ^ _64419;
  wire _64421 = _64416 ^ _64420;
  wire _64422 = _64412 ^ _64421;
  wire _64423 = _64399 ^ _64422;
  wire _64424 = _64378 ^ _64423;
  wire _64425 = uncoded_block[1348] ^ uncoded_block[1360];
  wire _64426 = uncoded_block[1361] ^ uncoded_block[1386];
  wire _64427 = _64425 ^ _64426;
  wire _64428 = uncoded_block[1387] ^ uncoded_block[1396];
  wire _64429 = uncoded_block[1406] ^ uncoded_block[1417];
  wire _64430 = _64428 ^ _64429;
  wire _64431 = _64427 ^ _64430;
  wire _64432 = uncoded_block[1422] ^ uncoded_block[1440];
  wire _64433 = _64432 ^ _5305;
  wire _64434 = uncoded_block[1461] ^ uncoded_block[1474];
  wire _64435 = uncoded_block[1484] ^ uncoded_block[1507];
  wire _64436 = _64434 ^ _64435;
  wire _64437 = _64433 ^ _64436;
  wire _64438 = _64431 ^ _64437;
  wire _64439 = _11266 ^ _5343;
  wire _64440 = _49954 ^ _62592;
  wire _64441 = _64439 ^ _64440;
  wire _64442 = uncoded_block[1577] ^ uncoded_block[1582];
  wire _64443 = uncoded_block[1604] ^ uncoded_block[1620];
  wire _64444 = _64442 ^ _64443;
  wire _64445 = uncoded_block[1623] ^ uncoded_block[1633];
  wire _64446 = _64445 ^ _26354;
  wire _64447 = _64444 ^ _64446;
  wire _64448 = _64441 ^ _64447;
  wire _64449 = _64438 ^ _64448;
  wire _64450 = uncoded_block[1666] ^ uncoded_block[1674];
  wire _64451 = _64450 ^ _41416;
  wire _64452 = uncoded_block[1692] ^ uncoded_block[1710];
  wire _64453 = _64452 ^ uncoded_block[1714];
  wire _64454 = _64451 ^ _64453;
  wire _64455 = _64449 ^ _64454;
  wire _64456 = _64424 ^ _64455;
  wire _64457 = uncoded_block[14] ^ uncoded_block[17];
  wire _64458 = _46913 ^ _64457;
  wire _64459 = uncoded_block[29] ^ uncoded_block[35];
  wire _64460 = _64459 ^ _31365;
  wire _64461 = _64458 ^ _64460;
  wire _64462 = uncoded_block[77] ^ uncoded_block[90];
  wire _64463 = _28008 ^ _64462;
  wire _64464 = uncoded_block[91] ^ uncoded_block[105];
  wire _64465 = _64464 ^ _16589;
  wire _64466 = _64463 ^ _64465;
  wire _64467 = _64461 ^ _64466;
  wire _64468 = uncoded_block[118] ^ uncoded_block[125];
  wire _64469 = uncoded_block[153] ^ uncoded_block[158];
  wire _64470 = _64468 ^ _64469;
  wire _64471 = uncoded_block[174] ^ uncoded_block[182];
  wire _64472 = _1749 ^ _64471;
  wire _64473 = _64470 ^ _64472;
  wire _64474 = uncoded_block[184] ^ uncoded_block[187];
  wire _64475 = uncoded_block[192] ^ uncoded_block[197];
  wire _64476 = _64474 ^ _64475;
  wire _64477 = uncoded_block[212] ^ uncoded_block[221];
  wire _64478 = uncoded_block[225] ^ uncoded_block[236];
  wire _64479 = _64477 ^ _64478;
  wire _64480 = _64476 ^ _64479;
  wire _64481 = _64473 ^ _64480;
  wire _64482 = _64467 ^ _64481;
  wire _64483 = uncoded_block[253] ^ uncoded_block[273];
  wire _64484 = _20021 ^ _64483;
  wire _64485 = _15159 ^ _35929;
  wire _64486 = _64484 ^ _64485;
  wire _64487 = uncoded_block[298] ^ uncoded_block[306];
  wire _64488 = _64487 ^ _48476;
  wire _64489 = uncoded_block[335] ^ uncoded_block[340];
  wire _64490 = uncoded_block[354] ^ uncoded_block[371];
  wire _64491 = _64489 ^ _64490;
  wire _64492 = _64488 ^ _64491;
  wire _64493 = _64486 ^ _64492;
  wire _64494 = uncoded_block[373] ^ uncoded_block[384];
  wire _64495 = _64494 ^ _12006;
  wire _64496 = uncoded_block[406] ^ uncoded_block[427];
  wire _64497 = _64496 ^ _42300;
  wire _64498 = _64495 ^ _64497;
  wire _64499 = uncoded_block[449] ^ uncoded_block[479];
  wire _64500 = _64499 ^ _2660;
  wire _64501 = _45982 ^ _8120;
  wire _64502 = _64500 ^ _64501;
  wire _64503 = _64498 ^ _64502;
  wire _64504 = _64493 ^ _64503;
  wire _64505 = _64482 ^ _64504;
  wire _64506 = uncoded_block[516] ^ uncoded_block[527];
  wire _64507 = _64506 ^ _35602;
  wire _64508 = uncoded_block[537] ^ uncoded_block[542];
  wire _64509 = uncoded_block[543] ^ uncoded_block[557];
  wire _64510 = _64508 ^ _64509;
  wire _64511 = _64507 ^ _64510;
  wire _64512 = _52447 ^ _6312;
  wire _64513 = uncoded_block[612] ^ uncoded_block[625];
  wire _64514 = _13705 ^ _64513;
  wire _64515 = _64512 ^ _64514;
  wire _64516 = _64511 ^ _64515;
  wire _64517 = _6966 ^ _42674;
  wire _64518 = uncoded_block[658] ^ uncoded_block[661];
  wire _64519 = _64518 ^ _7586;
  wire _64520 = _64517 ^ _64519;
  wire _64521 = uncoded_block[684] ^ uncoded_block[689];
  wire _64522 = _64521 ^ _9896;
  wire _64523 = uncoded_block[703] ^ uncoded_block[710];
  wire _64524 = uncoded_block[712] ^ uncoded_block[722];
  wire _64525 = _64523 ^ _64524;
  wire _64526 = _64522 ^ _64525;
  wire _64527 = _64520 ^ _64526;
  wire _64528 = _64516 ^ _64527;
  wire _64529 = uncoded_block[737] ^ uncoded_block[764];
  wire _64530 = _32779 ^ _64529;
  wire _64531 = uncoded_block[779] ^ uncoded_block[799];
  wire _64532 = _61850 ^ _64531;
  wire _64533 = _64530 ^ _64532;
  wire _64534 = uncoded_block[818] ^ uncoded_block[828];
  wire _64535 = _61859 ^ _64534;
  wire _64536 = uncoded_block[836] ^ uncoded_block[847];
  wire _64537 = _64536 ^ _16808;
  wire _64538 = _64535 ^ _64537;
  wire _64539 = _64533 ^ _64538;
  wire _64540 = uncoded_block[875] ^ uncoded_block[885];
  wire _64541 = _7650 ^ _64540;
  wire _64542 = uncoded_block[915] ^ uncoded_block[930];
  wire _64543 = _16312 ^ _64542;
  wire _64544 = _64541 ^ _64543;
  wire _64545 = _13809 ^ _7673;
  wire _64546 = uncoded_block[944] ^ uncoded_block[950];
  wire _64547 = uncoded_block[964] ^ uncoded_block[977];
  wire _64548 = _64546 ^ _64547;
  wire _64549 = _64545 ^ _64548;
  wire _64550 = _64544 ^ _64549;
  wire _64551 = _64539 ^ _64550;
  wire _64552 = _64528 ^ _64551;
  wire _64553 = _64505 ^ _64552;
  wire _64554 = uncoded_block[980] ^ uncoded_block[993];
  wire _64555 = uncoded_block[1008] ^ uncoded_block[1023];
  wire _64556 = _64554 ^ _64555;
  wire _64557 = uncoded_block[1026] ^ uncoded_block[1035];
  wire _64558 = _64557 ^ _2133;
  wire _64559 = _64556 ^ _64558;
  wire _64560 = _30731 ^ _2922;
  wire _64561 = _62070 ^ _534;
  wire _64562 = _64560 ^ _64561;
  wire _64563 = _64559 ^ _64562;
  wire _64564 = uncoded_block[1099] ^ uncoded_block[1107];
  wire _64565 = _64564 ^ _8920;
  wire _64566 = _56845 ^ _56555;
  wire _64567 = _64565 ^ _64566;
  wire _64568 = uncoded_block[1152] ^ uncoded_block[1159];
  wire _64569 = _64568 ^ _7151;
  wire _64570 = uncoded_block[1173] ^ uncoded_block[1187];
  wire _64571 = uncoded_block[1190] ^ uncoded_block[1199];
  wire _64572 = _64570 ^ _64571;
  wire _64573 = _64569 ^ _64572;
  wire _64574 = _64567 ^ _64573;
  wire _64575 = _64563 ^ _64574;
  wire _64576 = _49397 ^ _2989;
  wire _64577 = uncoded_block[1239] ^ uncoded_block[1252];
  wire _64578 = uncoded_block[1254] ^ uncoded_block[1261];
  wire _64579 = _64577 ^ _64578;
  wire _64580 = _64576 ^ _64579;
  wire _64581 = uncoded_block[1285] ^ uncoded_block[1294];
  wire _64582 = _59846 ^ _64581;
  wire _64583 = _4532 ^ _2254;
  wire _64584 = _64582 ^ _64583;
  wire _64585 = _64580 ^ _64584;
  wire _64586 = uncoded_block[1308] ^ uncoded_block[1318];
  wire _64587 = _64586 ^ _2277;
  wire _64588 = uncoded_block[1344] ^ uncoded_block[1356];
  wire _64589 = uncoded_block[1360] ^ uncoded_block[1373];
  wire _64590 = _64588 ^ _64589;
  wire _64591 = _64587 ^ _64590;
  wire _64592 = uncoded_block[1379] ^ uncoded_block[1387];
  wire _64593 = uncoded_block[1391] ^ uncoded_block[1397];
  wire _64594 = _64592 ^ _64593;
  wire _64595 = uncoded_block[1400] ^ uncoded_block[1414];
  wire _64596 = _64595 ^ _29508;
  wire _64597 = _64594 ^ _64596;
  wire _64598 = _64591 ^ _64597;
  wire _64599 = _64585 ^ _64598;
  wire _64600 = _64575 ^ _64599;
  wire _64601 = uncoded_block[1439] ^ uncoded_block[1446];
  wire _64602 = _64601 ^ _61370;
  wire _64603 = uncoded_block[1458] ^ uncoded_block[1489];
  wire _64604 = uncoded_block[1494] ^ uncoded_block[1505];
  wire _64605 = _64603 ^ _64604;
  wire _64606 = _64602 ^ _64605;
  wire _64607 = uncoded_block[1519] ^ uncoded_block[1534];
  wire _64608 = _64607 ^ _16995;
  wire _64609 = _4640 ^ _1612;
  wire _64610 = _64608 ^ _64609;
  wire _64611 = _64606 ^ _64610;
  wire _64612 = _3146 ^ _63974;
  wire _64613 = uncoded_block[1600] ^ uncoded_block[1611];
  wire _64614 = _64613 ^ _10745;
  wire _64615 = _64612 ^ _64614;
  wire _64616 = _14006 ^ _2405;
  wire _64617 = uncoded_block[1651] ^ uncoded_block[1658];
  wire _64618 = _64617 ^ _48771;
  wire _64619 = _64616 ^ _64618;
  wire _64620 = _64615 ^ _64619;
  wire _64621 = _64611 ^ _64620;
  wire _64622 = uncoded_block[1679] ^ uncoded_block[1688];
  wire _64623 = _64622 ^ _1669;
  wire _64624 = _64623 ^ uncoded_block[1704];
  wire _64625 = _64621 ^ _64624;
  wire _64626 = _64600 ^ _64625;
  wire _64627 = _64553 ^ _64626;
  wire _64628 = uncoded_block[9] ^ uncoded_block[18];
  wire _64629 = _64628 ^ _6728;
  wire _64630 = uncoded_block[36] ^ uncoded_block[50];
  wire _64631 = uncoded_block[60] ^ uncoded_block[73];
  wire _64632 = _64630 ^ _64631;
  wire _64633 = _64629 ^ _64632;
  wire _64634 = uncoded_block[94] ^ uncoded_block[106];
  wire _64635 = _58993 ^ _64634;
  wire _64636 = uncoded_block[121] ^ uncoded_block[129];
  wire _64637 = _35117 ^ _64636;
  wire _64638 = _64635 ^ _64637;
  wire _64639 = _64633 ^ _64638;
  wire _64640 = uncoded_block[140] ^ uncoded_block[156];
  wire _64641 = _64640 ^ _19536;
  wire _64642 = _4766 ^ _941;
  wire _64643 = _64641 ^ _64642;
  wire _64644 = uncoded_block[200] ^ uncoded_block[211];
  wire _64645 = _16114 ^ _64644;
  wire _64646 = uncoded_block[236] ^ uncoded_block[240];
  wire _64647 = _64646 ^ _8616;
  wire _64648 = _64645 ^ _64647;
  wire _64649 = _64643 ^ _64648;
  wire _64650 = _64639 ^ _64649;
  wire _64651 = uncoded_block[256] ^ uncoded_block[279];
  wire _64652 = _6182 ^ _64651;
  wire _64653 = _19072 ^ _13615;
  wire _64654 = _64652 ^ _64653;
  wire _64655 = _9779 ^ _1819;
  wire _64656 = _64489 ^ _38366;
  wire _64657 = _64655 ^ _64656;
  wire _64658 = _64654 ^ _64657;
  wire _64659 = _39961 ^ _10340;
  wire _64660 = uncoded_block[426] ^ uncoded_block[439];
  wire _64661 = _4874 ^ _64660;
  wire _64662 = _64659 ^ _64661;
  wire _64663 = uncoded_block[449] ^ uncoded_block[457];
  wire _64664 = _5580 ^ _64663;
  wire _64665 = uncoded_block[462] ^ uncoded_block[468];
  wire _64666 = _64665 ^ _14176;
  wire _64667 = _64664 ^ _64666;
  wire _64668 = _64662 ^ _64667;
  wire _64669 = _64658 ^ _64668;
  wire _64670 = _64650 ^ _64669;
  wire _64671 = uncoded_block[510] ^ uncoded_block[520];
  wire _64672 = _3424 ^ _64671;
  wire _64673 = uncoded_block[525] ^ uncoded_block[530];
  wire _64674 = _64673 ^ _18670;
  wire _64675 = _64672 ^ _64674;
  wire _64676 = _61290 ^ _7550;
  wire _64677 = uncoded_block[586] ^ uncoded_block[598];
  wire _64678 = _62676 ^ _64677;
  wire _64679 = _64676 ^ _64678;
  wire _64680 = _64675 ^ _64679;
  wire _64681 = uncoded_block[606] ^ uncoded_block[615];
  wire _64682 = _64681 ^ _12071;
  wire _64683 = uncoded_block[636] ^ uncoded_block[648];
  wire _64684 = _64683 ^ _34829;
  wire _64685 = _64682 ^ _64684;
  wire _64686 = uncoded_block[685] ^ uncoded_block[692];
  wire _64687 = _43772 ^ _64686;
  wire _64688 = uncoded_block[706] ^ uncoded_block[714];
  wire _64689 = _55600 ^ _64688;
  wire _64690 = _64687 ^ _64689;
  wire _64691 = _64685 ^ _64690;
  wire _64692 = _64680 ^ _64691;
  wire _64693 = uncoded_block[731] ^ uncoded_block[743];
  wire _64694 = _64693 ^ _11012;
  wire _64695 = _13215 ^ _58824;
  wire _64696 = _64694 ^ _64695;
  wire _64697 = _19705 ^ _33218;
  wire _64698 = uncoded_block[799] ^ uncoded_block[812];
  wire _64699 = _64698 ^ _31971;
  wire _64700 = _64697 ^ _64699;
  wire _64701 = _64696 ^ _64700;
  wire _64702 = uncoded_block[847] ^ uncoded_block[854];
  wire _64703 = _11607 ^ _64702;
  wire _64704 = uncoded_block[855] ^ uncoded_block[875];
  wire _64705 = uncoded_block[897] ^ uncoded_block[902];
  wire _64706 = _64704 ^ _64705;
  wire _64707 = _64703 ^ _64706;
  wire _64708 = uncoded_block[931] ^ uncoded_block[941];
  wire _64709 = _61669 ^ _64708;
  wire _64710 = _9433 ^ _2871;
  wire _64711 = _64709 ^ _64710;
  wire _64712 = _64707 ^ _64711;
  wire _64713 = _64701 ^ _64712;
  wire _64714 = _64692 ^ _64713;
  wire _64715 = _64670 ^ _64714;
  wire _64716 = _10537 ^ _24400;
  wire _64717 = _61684 ^ _50575;
  wire _64718 = _64716 ^ _64717;
  wire _64719 = _58865 ^ _8892;
  wire _64720 = uncoded_block[1082] ^ uncoded_block[1094];
  wire _64721 = _64720 ^ _2938;
  wire _64722 = _64719 ^ _64721;
  wire _64723 = _64718 ^ _64722;
  wire _64724 = uncoded_block[1140] ^ uncoded_block[1154];
  wire _64725 = _56845 ^ _64724;
  wire _64726 = _2964 ^ _10608;
  wire _64727 = _64725 ^ _64726;
  wire _64728 = uncoded_block[1189] ^ uncoded_block[1211];
  wire _64729 = _64728 ^ _49397;
  wire _64730 = _64729 ^ _58894;
  wire _64731 = _64727 ^ _64730;
  wire _64732 = _64723 ^ _64731;
  wire _64733 = _19827 ^ _60702;
  wire _64734 = uncoded_block[1263] ^ uncoded_block[1282];
  wire _64735 = _64734 ^ _18866;
  wire _64736 = _64733 ^ _64735;
  wire _64737 = _21741 ^ _10081;
  wire _64738 = uncoded_block[1308] ^ uncoded_block[1327];
  wire _64739 = uncoded_block[1335] ^ uncoded_block[1341];
  wire _64740 = _64738 ^ _64739;
  wire _64741 = _64737 ^ _64740;
  wire _64742 = _64736 ^ _64741;
  wire _64743 = _46096 ^ _15477;
  wire _64744 = _4564 ^ _1517;
  wire _64745 = _64743 ^ _64744;
  wire _64746 = _10678 ^ _3850;
  wire _64747 = uncoded_block[1439] ^ uncoded_block[1459];
  wire _64748 = uncoded_block[1465] ^ uncoded_block[1475];
  wire _64749 = _64747 ^ _64748;
  wire _64750 = _64746 ^ _64749;
  wire _64751 = _64745 ^ _64750;
  wire _64752 = _64742 ^ _64751;
  wire _64753 = _64732 ^ _64752;
  wire _64754 = uncoded_block[1491] ^ uncoded_block[1513];
  wire _64755 = uncoded_block[1519] ^ uncoded_block[1541];
  wire _64756 = _64754 ^ _64755;
  wire _64757 = uncoded_block[1545] ^ uncoded_block[1554];
  wire _64758 = _64757 ^ _48748;
  wire _64759 = _64756 ^ _64758;
  wire _64760 = uncoded_block[1567] ^ uncoded_block[1590];
  wire _64761 = _5361 ^ _64760;
  wire _64762 = _12935 ^ _6674;
  wire _64763 = _64761 ^ _64762;
  wire _64764 = _64759 ^ _64763;
  wire _64765 = uncoded_block[1602] ^ uncoded_block[1613];
  wire _64766 = _64765 ^ _24115;
  wire _64767 = uncoded_block[1656] ^ uncoded_block[1666];
  wire _64768 = _59903 ^ _64767;
  wire _64769 = _64766 ^ _64768;
  wire _64770 = uncoded_block[1681] ^ uncoded_block[1694];
  wire _64771 = _8521 ^ _64770;
  wire _64772 = _64771 ^ _3989;
  wire _64773 = _64769 ^ _64772;
  wire _64774 = _64764 ^ _64773;
  wire _64775 = _64753 ^ _64774;
  wire _64776 = _64715 ^ _64775;
  wire _64777 = uncoded_block[20] ^ uncoded_block[47];
  wire _64778 = uncoded_block[51] ^ uncoded_block[62];
  wire _64779 = _64777 ^ _64778;
  wire _64780 = uncoded_block[85] ^ uncoded_block[104];
  wire _64781 = uncoded_block[136] ^ uncoded_block[166];
  wire _64782 = _64780 ^ _64781;
  wire _64783 = _64779 ^ _64782;
  wire _64784 = uncoded_block[168] ^ uncoded_block[194];
  wire _64785 = uncoded_block[195] ^ uncoded_block[206];
  wire _64786 = _64784 ^ _64785;
  wire _64787 = uncoded_block[232] ^ uncoded_block[246];
  wire _64788 = uncoded_block[266] ^ uncoded_block[281];
  wire _64789 = _64787 ^ _64788;
  wire _64790 = _64786 ^ _64789;
  wire _64791 = _64783 ^ _64790;
  wire _64792 = uncoded_block[301] ^ uncoded_block[317];
  wire _64793 = uncoded_block[363] ^ uncoded_block[386];
  wire _64794 = _64792 ^ _64793;
  wire _64795 = uncoded_block[389] ^ uncoded_block[407];
  wire _64796 = uncoded_block[428] ^ uncoded_block[436];
  wire _64797 = _64795 ^ _64796;
  wire _64798 = _64794 ^ _64797;
  wire _64799 = uncoded_block[450] ^ uncoded_block[463];
  wire _64800 = uncoded_block[502] ^ uncoded_block[536];
  wire _64801 = _64799 ^ _64800;
  wire _64802 = uncoded_block[542] ^ uncoded_block[556];
  wire _64803 = _64802 ^ _17221;
  wire _64804 = _64801 ^ _64803;
  wire _64805 = _64798 ^ _64804;
  wire _64806 = _64791 ^ _64805;
  wire _64807 = uncoded_block[593] ^ uncoded_block[624];
  wire _64808 = uncoded_block[629] ^ uncoded_block[641];
  wire _64809 = _64807 ^ _64808;
  wire _64810 = uncoded_block[671] ^ uncoded_block[713];
  wire _64811 = uncoded_block[715] ^ uncoded_block[732];
  wire _64812 = _64810 ^ _64811;
  wire _64813 = _64809 ^ _64812;
  wire _64814 = uncoded_block[798] ^ uncoded_block[822];
  wire _64815 = _60534 ^ _64814;
  wire _64816 = uncoded_block[857] ^ uncoded_block[878];
  wire _64817 = _54070 ^ _64816;
  wire _64818 = _64815 ^ _64817;
  wire _64819 = _64813 ^ _64818;
  wire _64820 = uncoded_block[898] ^ uncoded_block[921];
  wire _64821 = uncoded_block[933] ^ uncoded_block[948];
  wire _64822 = _64820 ^ _64821;
  wire _64823 = uncoded_block[959] ^ uncoded_block[999];
  wire _64824 = _64823 ^ _49571;
  wire _64825 = _64822 ^ _64824;
  wire _64826 = uncoded_block[1050] ^ uncoded_block[1063];
  wire _64827 = uncoded_block[1076] ^ uncoded_block[1099];
  wire _64828 = _64826 ^ _64827;
  wire _64829 = uncoded_block[1108] ^ uncoded_block[1141];
  wire _64830 = uncoded_block[1162] ^ uncoded_block[1173];
  wire _64831 = _64829 ^ _64830;
  wire _64832 = _64828 ^ _64831;
  wire _64833 = _64825 ^ _64832;
  wire _64834 = _64819 ^ _64833;
  wire _64835 = _64806 ^ _64834;
  wire _64836 = _1428 ^ _17910;
  wire _64837 = uncoded_block[1248] ^ uncoded_block[1303];
  wire _64838 = uncoded_block[1314] ^ uncoded_block[1331];
  wire _64839 = _64837 ^ _64838;
  wire _64840 = _64836 ^ _64839;
  wire _64841 = uncoded_block[1354] ^ uncoded_block[1388];
  wire _64842 = uncoded_block[1414] ^ uncoded_block[1431];
  wire _64843 = _64841 ^ _64842;
  wire _64844 = uncoded_block[1448] ^ uncoded_block[1464];
  wire _64845 = uncoded_block[1484] ^ uncoded_block[1495];
  wire _64846 = _64844 ^ _64845;
  wire _64847 = _64843 ^ _64846;
  wire _64848 = _64840 ^ _64847;
  wire _64849 = uncoded_block[1511] ^ uncoded_block[1532];
  wire _64850 = _64849 ^ _14506;
  wire _64851 = uncoded_block[1606] ^ uncoded_block[1614];
  wire _64852 = uncoded_block[1624] ^ uncoded_block[1652];
  wire _64853 = _64851 ^ _64852;
  wire _64854 = _64850 ^ _64853;
  wire _64855 = uncoded_block[1661] ^ uncoded_block[1690];
  wire _64856 = _64855 ^ uncoded_block[1708];
  wire _64857 = _64854 ^ _64856;
  wire _64858 = _64848 ^ _64857;
  wire _64859 = _64835 ^ _64858;
  wire _64860 = _32201 ^ _42204;
  wire _64861 = uncoded_block[29] ^ uncoded_block[37];
  wire _64862 = uncoded_block[52] ^ uncoded_block[61];
  wire _64863 = _64861 ^ _64862;
  wire _64864 = _64860 ^ _64863;
  wire _64865 = uncoded_block[66] ^ uncoded_block[71];
  wire _64866 = _64865 ^ _6113;
  wire _64867 = uncoded_block[98] ^ uncoded_block[105];
  wire _64868 = _7374 ^ _64867;
  wire _64869 = _64866 ^ _64868;
  wire _64870 = _64864 ^ _64869;
  wire _64871 = uncoded_block[117] ^ uncoded_block[130];
  wire _64872 = _64871 ^ _4761;
  wire _64873 = _39508 ^ _64872;
  wire _64874 = uncoded_block[151] ^ uncoded_block[174];
  wire _64875 = _14082 ^ _64874;
  wire _64876 = uncoded_block[181] ^ uncoded_block[194];
  wire _64877 = _64876 ^ _95;
  wire _64878 = _64875 ^ _64877;
  wire _64879 = _64873 ^ _64878;
  wire _64880 = _64870 ^ _64879;
  wire _64881 = _9747 ^ _6161;
  wire _64882 = uncoded_block[221] ^ uncoded_block[232];
  wire _64883 = _64882 ^ _35141;
  wire _64884 = _64881 ^ _64883;
  wire _64885 = uncoded_block[248] ^ uncoded_block[254];
  wire _64886 = _63787 ^ _64885;
  wire _64887 = uncoded_block[267] ^ uncoded_block[287];
  wire _64888 = _64887 ^ _38762;
  wire _64889 = _64886 ^ _64888;
  wire _64890 = _64884 ^ _64889;
  wire _64891 = uncoded_block[308] ^ uncoded_block[316];
  wire _64892 = _21016 ^ _64891;
  wire _64893 = uncoded_block[319] ^ uncoded_block[326];
  wire _64894 = uncoded_block[331] ^ uncoded_block[336];
  wire _64895 = _64893 ^ _64894;
  wire _64896 = _64892 ^ _64895;
  wire _64897 = uncoded_block[345] ^ uncoded_block[361];
  wire _64898 = uncoded_block[362] ^ uncoded_block[368];
  wire _64899 = _64897 ^ _64898;
  wire _64900 = uncoded_block[374] ^ uncoded_block[379];
  wire _64901 = uncoded_block[386] ^ uncoded_block[392];
  wire _64902 = _64900 ^ _64901;
  wire _64903 = _64899 ^ _64902;
  wire _64904 = _64896 ^ _64903;
  wire _64905 = _64890 ^ _64904;
  wire _64906 = _64880 ^ _64905;
  wire _64907 = uncoded_block[411] ^ uncoded_block[415];
  wire _64908 = _10910 ^ _64907;
  wire _64909 = uncoded_block[418] ^ uncoded_block[438];
  wire _64910 = _64909 ^ _3405;
  wire _64911 = _64908 ^ _64910;
  wire _64912 = uncoded_block[443] ^ uncoded_block[454];
  wire _64913 = _64912 ^ _1871;
  wire _64914 = uncoded_block[463] ^ uncoded_block[473];
  wire _64915 = uncoded_block[474] ^ uncoded_block[484];
  wire _64916 = _64914 ^ _64915;
  wire _64917 = _64913 ^ _64916;
  wire _64918 = _64911 ^ _64917;
  wire _64919 = uncoded_block[488] ^ uncoded_block[496];
  wire _64920 = _64919 ^ _64043;
  wire _64921 = _26080 ^ _24279;
  wire _64922 = _64920 ^ _64921;
  wire _64923 = _6945 ^ _19652;
  wire _64924 = _2689 ^ _64923;
  wire _64925 = _64922 ^ _64924;
  wire _64926 = _64918 ^ _64925;
  wire _64927 = uncoded_block[606] ^ uncoded_block[613];
  wire _64928 = _56740 ^ _64927;
  wire _64929 = uncoded_block[617] ^ uncoded_block[625];
  wire _64930 = _64929 ^ _45999;
  wire _64931 = _64928 ^ _64930;
  wire _64932 = uncoded_block[636] ^ uncoded_block[650];
  wire _64933 = uncoded_block[651] ^ uncoded_block[666];
  wire _64934 = _64932 ^ _64933;
  wire _64935 = _4265 ^ _3527;
  wire _64936 = _64934 ^ _64935;
  wire _64937 = _64931 ^ _64936;
  wire _64938 = uncoded_block[692] ^ uncoded_block[721];
  wire _64939 = _64938 ^ _1991;
  wire _64940 = uncoded_block[742] ^ uncoded_block[754];
  wire _64941 = _23870 ^ _64940;
  wire _64942 = _64939 ^ _64941;
  wire _64943 = _13219 ^ _8790;
  wire _64944 = uncoded_block[797] ^ uncoded_block[803];
  wire _64945 = uncoded_block[814] ^ uncoded_block[819];
  wire _64946 = _64944 ^ _64945;
  wire _64947 = _64943 ^ _64946;
  wire _64948 = _64942 ^ _64947;
  wire _64949 = _64937 ^ _64948;
  wire _64950 = _64926 ^ _64949;
  wire _64951 = _64906 ^ _64950;
  wire _64952 = _3590 ^ _35668;
  wire _64953 = uncoded_block[841] ^ uncoded_block[854];
  wire _64954 = uncoded_block[859] ^ uncoded_block[868];
  wire _64955 = _64953 ^ _64954;
  wire _64956 = _64952 ^ _64955;
  wire _64957 = uncoded_block[871] ^ uncoded_block[881];
  wire _64958 = uncoded_block[883] ^ uncoded_block[891];
  wire _64959 = _64957 ^ _64958;
  wire _64960 = uncoded_block[897] ^ uncoded_block[904];
  wire _64961 = uncoded_block[907] ^ uncoded_block[912];
  wire _64962 = _64960 ^ _64961;
  wire _64963 = _64959 ^ _64962;
  wire _64964 = _64956 ^ _64963;
  wire _64965 = uncoded_block[937] ^ uncoded_block[957];
  wire _64966 = _49563 ^ _64965;
  wire _64967 = _4385 ^ _24388;
  wire _64968 = _64966 ^ _64967;
  wire _64969 = _5789 ^ _61177;
  wire _64970 = uncoded_block[998] ^ uncoded_block[1017];
  wire _64971 = _64970 ^ _2121;
  wire _64972 = _64969 ^ _64971;
  wire _64973 = _64968 ^ _64972;
  wire _64974 = _64964 ^ _64973;
  wire _64975 = uncoded_block[1040] ^ uncoded_block[1057];
  wire _64976 = _9461 ^ _64975;
  wire _64977 = uncoded_block[1059] ^ uncoded_block[1067];
  wire _64978 = _64977 ^ _13851;
  wire _64979 = _64976 ^ _64978;
  wire _64980 = _61689 ^ _23071;
  wire _64981 = _64980 ^ _11144;
  wire _64982 = _64979 ^ _64981;
  wire _64983 = uncoded_block[1117] ^ uncoded_block[1127];
  wire _64984 = uncoded_block[1130] ^ uncoded_block[1146];
  wire _64985 = _64983 ^ _64984;
  wire _64986 = _7143 ^ _12243;
  wire _64987 = _64985 ^ _64986;
  wire _64988 = _7151 ^ _3742;
  wire _64989 = _1417 ^ _10612;
  wire _64990 = _64988 ^ _64989;
  wire _64991 = _64987 ^ _64990;
  wire _64992 = _64982 ^ _64991;
  wire _64993 = _64974 ^ _64992;
  wire _64994 = uncoded_block[1239] ^ uncoded_block[1245];
  wire _64995 = _21723 ^ _64994;
  wire _64996 = _3783 ^ _57498;
  wire _64997 = _64995 ^ _64996;
  wire _64998 = uncoded_block[1288] ^ uncoded_block[1298];
  wire _64999 = _64998 ^ _648;
  wire _65000 = uncoded_block[1311] ^ uncoded_block[1320];
  wire _65001 = _65000 ^ _19375;
  wire _65002 = _64999 ^ _65001;
  wire _65003 = _64997 ^ _65002;
  wire _65004 = uncoded_block[1327] ^ uncoded_block[1339];
  wire _65005 = _65004 ^ _46096;
  wire _65006 = _11218 ^ _21762;
  wire _65007 = _65005 ^ _65006;
  wire _65008 = _57192 ^ _9578;
  wire _65009 = _16458 ^ _57527;
  wire _65010 = _65008 ^ _65009;
  wire _65011 = _65007 ^ _65010;
  wire _65012 = _65003 ^ _65011;
  wire _65013 = uncoded_block[1422] ^ uncoded_block[1428];
  wire _65014 = _8438 ^ _65013;
  wire _65015 = uncoded_block[1442] ^ uncoded_block[1460];
  wire _65016 = _13432 ^ _65015;
  wire _65017 = _65014 ^ _65016;
  wire _65018 = uncoded_block[1466] ^ uncoded_block[1472];
  wire _65019 = uncoded_block[1475] ^ uncoded_block[1480];
  wire _65020 = _65018 ^ _65019;
  wire _65021 = _5320 ^ _1562;
  wire _65022 = _65020 ^ _65021;
  wire _65023 = _65017 ^ _65022;
  wire _65024 = uncoded_block[1492] ^ uncoded_block[1497];
  wire _65025 = _65024 ^ _9618;
  wire _65026 = _8467 ^ _12352;
  wire _65027 = _65025 ^ _65026;
  wire _65028 = _19899 ^ _31309;
  wire _65029 = _3131 ^ _55416;
  wire _65030 = _65028 ^ _65029;
  wire _65031 = _65027 ^ _65030;
  wire _65032 = _65023 ^ _65031;
  wire _65033 = _65012 ^ _65032;
  wire _65034 = _64993 ^ _65033;
  wire _65035 = _64951 ^ _65034;
  wire _65036 = _16515 ^ _11294;
  wire _65037 = uncoded_block[1599] ^ uncoded_block[1610];
  wire _65038 = _65037 ^ _6046;
  wire _65039 = _65036 ^ _65038;
  wire _65040 = uncoded_block[1633] ^ uncoded_block[1639];
  wire _65041 = _65040 ^ _43612;
  wire _65042 = _19471 ^ _31339;
  wire _65043 = _65041 ^ _65042;
  wire _65044 = _65039 ^ _65043;
  wire _65045 = _14545 ^ _5409;
  wire _65046 = uncoded_block[1700] ^ uncoded_block[1717];
  wire _65047 = _65046 ^ uncoded_block[1722];
  wire _65048 = _65045 ^ _65047;
  wire _65049 = _65044 ^ _65048;
  wire _65050 = _65035 ^ _65049;
  wire _65051 = uncoded_block[3] ^ uncoded_block[10];
  wire _65052 = _65051 ^ _34676;
  wire _65053 = uncoded_block[23] ^ uncoded_block[34];
  wire _65054 = _65053 ^ _879;
  wire _65055 = _65052 ^ _65054;
  wire _65056 = _18 ^ _62130;
  wire _65057 = _65056 ^ _42859;
  wire _65058 = _65055 ^ _65057;
  wire _65059 = uncoded_block[61] ^ uncoded_block[66];
  wire _65060 = uncoded_block[68] ^ uncoded_block[94];
  wire _65061 = _65059 ^ _65060;
  wire _65062 = _15097 ^ _58998;
  wire _65063 = _65061 ^ _65062;
  wire _65064 = _2497 ^ _1730;
  wire _65065 = uncoded_block[136] ^ uncoded_block[142];
  wire _65066 = _923 ^ _65065;
  wire _65067 = _65064 ^ _65066;
  wire _65068 = _65063 ^ _65067;
  wire _65069 = _65058 ^ _65068;
  wire _65070 = uncoded_block[152] ^ uncoded_block[163];
  wire _65071 = _15622 ^ _65070;
  wire _65072 = uncoded_block[168] ^ uncoded_block[173];
  wire _65073 = _65072 ^ _7403;
  wire _65074 = _65071 ^ _65073;
  wire _65075 = _28037 ^ _89;
  wire _65076 = uncoded_block[198] ^ uncoded_block[207];
  wire _65077 = _65076 ^ _21459;
  wire _65078 = _65075 ^ _65077;
  wire _65079 = _65074 ^ _65078;
  wire _65080 = _24657 ^ _10292;
  wire _65081 = _6180 ^ _64885;
  wire _65082 = _65080 ^ _65081;
  wire _65083 = uncoded_block[266] ^ uncoded_block[272];
  wire _65084 = _6185 ^ _65083;
  wire _65085 = uncoded_block[273] ^ uncoded_block[285];
  wire _65086 = _65085 ^ _56439;
  wire _65087 = _65084 ^ _65086;
  wire _65088 = _65082 ^ _65087;
  wire _65089 = _65079 ^ _65088;
  wire _65090 = _65069 ^ _65089;
  wire _65091 = _40724 ^ _40726;
  wire _65092 = _41502 ^ _9782;
  wire _65093 = _65091 ^ _65092;
  wire _65094 = _25577 ^ _6857;
  wire _65095 = uncoded_block[349] ^ uncoded_block[360];
  wire _65096 = _37186 ^ _65095;
  wire _65097 = _65094 ^ _65096;
  wire _65098 = _65093 ^ _65097;
  wire _65099 = _30569 ^ _4853;
  wire _65100 = uncoded_block[389] ^ uncoded_block[395];
  wire _65101 = _35563 ^ _65100;
  wire _65102 = _65099 ^ _65101;
  wire _65103 = _180 ^ _2625;
  wire _65104 = _1054 ^ _193;
  wire _65105 = _65103 ^ _65104;
  wire _65106 = _65102 ^ _65105;
  wire _65107 = _65098 ^ _65106;
  wire _65108 = _24707 ^ _17177;
  wire _65109 = uncoded_block[431] ^ uncoded_block[453];
  wire _65110 = _65109 ^ _13662;
  wire _65111 = _65108 ^ _65110;
  wire _65112 = uncoded_block[464] ^ uncoded_block[471];
  wire _65113 = _65112 ^ _2657;
  wire _65114 = uncoded_block[486] ^ uncoded_block[494];
  wire _65115 = _1086 ^ _65114;
  wire _65116 = _65113 ^ _65115;
  wire _65117 = _65111 ^ _65116;
  wire _65118 = uncoded_block[504] ^ uncoded_block[514];
  wire _65119 = _65118 ^ _6286;
  wire _65120 = uncoded_block[523] ^ uncoded_block[531];
  wire _65121 = _65120 ^ _44903;
  wire _65122 = _65119 ^ _65121;
  wire _65123 = _18670 ^ _43741;
  wire _65124 = uncoded_block[565] ^ uncoded_block[570];
  wire _65125 = _31907 ^ _65124;
  wire _65126 = _65123 ^ _65125;
  wire _65127 = _65122 ^ _65126;
  wire _65128 = _65117 ^ _65127;
  wire _65129 = _65107 ^ _65128;
  wire _65130 = _65090 ^ _65129;
  wire _65131 = _3475 ^ _37247;
  wire _65132 = _65131 ^ _25193;
  wire _65133 = uncoded_block[602] ^ uncoded_block[607];
  wire _65134 = _65133 ^ _6957;
  wire _65135 = uncoded_block[624] ^ uncoded_block[630];
  wire _65136 = _43759 ^ _65135;
  wire _65137 = _65134 ^ _65136;
  wire _65138 = _65132 ^ _65137;
  wire _65139 = _4972 ^ _41955;
  wire _65140 = _24303 ^ _65139;
  wire _65141 = _6342 ^ _20643;
  wire _65142 = _1178 ^ _8761;
  wire _65143 = _65141 ^ _65142;
  wire _65144 = _65140 ^ _65143;
  wire _65145 = _65138 ^ _65144;
  wire _65146 = _9891 ^ _5685;
  wire _65147 = uncoded_block[718] ^ uncoded_block[724];
  wire _65148 = _6366 ^ _65147;
  wire _65149 = _65146 ^ _65148;
  wire _65150 = uncoded_block[738] ^ uncoded_block[750];
  wire _65151 = _65150 ^ _15310;
  wire _65152 = _46301 ^ _65151;
  wire _65153 = _65149 ^ _65152;
  wire _65154 = uncoded_block[776] ^ uncoded_block[781];
  wire _65155 = _65154 ^ _25694;
  wire _65156 = _374 ^ _11024;
  wire _65157 = _65155 ^ _65156;
  wire _65158 = uncoded_block[804] ^ uncoded_block[818];
  wire _65159 = _7029 ^ _65158;
  wire _65160 = _45332 ^ _17793;
  wire _65161 = _65159 ^ _65160;
  wire _65162 = _65157 ^ _65161;
  wire _65163 = _65153 ^ _65162;
  wire _65164 = _65145 ^ _65163;
  wire _65165 = _33659 ^ _23010;
  wire _65166 = _413 ^ _1266;
  wire _65167 = _65165 ^ _65166;
  wire _65168 = uncoded_block[887] ^ uncoded_block[893];
  wire _65169 = _423 ^ _65168;
  wire _65170 = _39682 ^ _65169;
  wire _65171 = _65167 ^ _65170;
  wire _65172 = _45355 ^ _1281;
  wire _65173 = _435 ^ _18775;
  wire _65174 = _65172 ^ _65173;
  wire _65175 = uncoded_block[934] ^ uncoded_block[940];
  wire _65176 = _26623 ^ _65175;
  wire _65177 = _48621 ^ _14329;
  wire _65178 = _65176 ^ _65177;
  wire _65179 = _65174 ^ _65178;
  wire _65180 = _65171 ^ _65179;
  wire _65181 = uncoded_block[960] ^ uncoded_block[968];
  wire _65182 = _7680 ^ _65181;
  wire _65183 = _61678 ^ _6451;
  wire _65184 = _65182 ^ _65183;
  wire _65185 = uncoded_block[991] ^ uncoded_block[998];
  wire _65186 = _65185 ^ _1326;
  wire _65187 = _13835 ^ _61684;
  wire _65188 = _65186 ^ _65187;
  wire _65189 = _65184 ^ _65188;
  wire _65190 = _12752 ^ _8875;
  wire _65191 = _5806 ^ _12758;
  wire _65192 = _65190 ^ _65191;
  wire _65193 = uncoded_block[1054] ^ uncoded_block[1070];
  wire _65194 = _22135 ^ _65193;
  wire _65195 = _527 ^ _17363;
  wire _65196 = _65194 ^ _65195;
  wire _65197 = _65192 ^ _65196;
  wire _65198 = _65189 ^ _65197;
  wire _65199 = _65180 ^ _65198;
  wire _65200 = _65164 ^ _65199;
  wire _65201 = _65130 ^ _65200;
  wire _65202 = _52906 ^ _46770;
  wire _65203 = uncoded_block[1109] ^ uncoded_block[1114];
  wire _65204 = _65203 ^ _3713;
  wire _65205 = _65202 ^ _65204;
  wire _65206 = uncoded_block[1127] ^ uncoded_block[1132];
  wire _65207 = _46066 ^ _65206;
  wire _65208 = uncoded_block[1133] ^ uncoded_block[1140];
  wire _65209 = _65208 ^ _43874;
  wire _65210 = _65207 ^ _65209;
  wire _65211 = _65205 ^ _65210;
  wire _65212 = uncoded_block[1153] ^ uncoded_block[1162];
  wire _65213 = _65212 ^ _2964;
  wire _65214 = _17390 ^ _585;
  wire _65215 = _65213 ^ _65214;
  wire _65216 = _5200 ^ _1418;
  wire _65217 = uncoded_block[1200] ^ uncoded_block[1209];
  wire _65218 = _2971 ^ _65217;
  wire _65219 = _65216 ^ _65218;
  wire _65220 = _65215 ^ _65219;
  wire _65221 = _65211 ^ _65220;
  wire _65222 = _40908 ^ _5215;
  wire _65223 = _612 ^ _17908;
  wire _65224 = _65222 ^ _65223;
  wire _65225 = uncoded_block[1246] ^ uncoded_block[1254];
  wire _65226 = _17910 ^ _65225;
  wire _65227 = uncoded_block[1274] ^ uncoded_block[1281];
  wire _65228 = _46419 ^ _65227;
  wire _65229 = _65226 ^ _65228;
  wire _65230 = _65224 ^ _65229;
  wire _65231 = _1471 ^ _3807;
  wire _65232 = _56878 ^ _65231;
  wire _65233 = uncoded_block[1313] ^ uncoded_block[1323];
  wire _65234 = _13917 ^ _65233;
  wire _65235 = uncoded_block[1328] ^ uncoded_block[1333];
  wire _65236 = _65235 ^ _4551;
  wire _65237 = _65234 ^ _65236;
  wire _65238 = _65232 ^ _65237;
  wire _65239 = _65230 ^ _65238;
  wire _65240 = _65221 ^ _65239;
  wire _65241 = _20327 ^ _3047;
  wire _65242 = _7816 ^ _65241;
  wire _65243 = uncoded_block[1382] ^ uncoded_block[1391];
  wire _65244 = _57192 ^ _65243;
  wire _65245 = _30821 ^ _701;
  wire _65246 = _65244 ^ _65245;
  wire _65247 = _65242 ^ _65246;
  wire _65248 = uncoded_block[1427] ^ uncoded_block[1433];
  wire _65249 = _6606 ^ _65248;
  wire _65250 = _65249 ^ _21789;
  wire _65251 = uncoded_block[1449] ^ uncoded_block[1455];
  wire _65252 = _65251 ^ _12335;
  wire _65253 = _24071 ^ _5316;
  wire _65254 = _65252 ^ _65253;
  wire _65255 = _65250 ^ _65254;
  wire _65256 = _65247 ^ _65255;
  wire _65257 = uncoded_block[1483] ^ uncoded_block[1491];
  wire _65258 = _13963 ^ _65257;
  wire _65259 = _9614 ^ _747;
  wire _65260 = _65258 ^ _65259;
  wire _65261 = _4616 ^ _17499;
  wire _65262 = uncoded_block[1551] ^ uncoded_block[1558];
  wire _65263 = _65262 ^ _28386;
  wire _65264 = _65261 ^ _65263;
  wire _65265 = _65260 ^ _65264;
  wire _65266 = _60599 ^ _13479;
  wire _65267 = _65266 ^ _21828;
  wire _65268 = uncoded_block[1603] ^ uncoded_block[1611];
  wire _65269 = _65268 ^ _20409;
  wire _65270 = uncoded_block[1626] ^ uncoded_block[1633];
  wire _65271 = _27215 ^ _65270;
  wire _65272 = _65269 ^ _65271;
  wire _65273 = _65267 ^ _65272;
  wire _65274 = _65265 ^ _65273;
  wire _65275 = _65256 ^ _65274;
  wire _65276 = _65240 ^ _65275;
  wire _65277 = _4668 ^ _44393;
  wire _65278 = _4674 ^ _30008;
  wire _65279 = _65277 ^ _65278;
  wire _65280 = uncoded_block[1662] ^ uncoded_block[1669];
  wire _65281 = _65280 ^ _19471;
  wire _65282 = _61978 ^ _16060;
  wire _65283 = _65281 ^ _65282;
  wire _65284 = _65279 ^ _65283;
  wire _65285 = _3972 ^ _8533;
  wire _65286 = _2438 ^ uncoded_block[1719];
  wire _65287 = _65285 ^ _65286;
  wire _65288 = _65284 ^ _65287;
  wire _65289 = _65276 ^ _65288;
  wire _65290 = _65201 ^ _65289;
  wire _65291 = uncoded_block[10] ^ uncoded_block[90];
  wire _65292 = uncoded_block[98] ^ uncoded_block[113];
  wire _65293 = _65291 ^ _65292;
  wire _65294 = uncoded_block[142] ^ uncoded_block[194];
  wire _65295 = uncoded_block[200] ^ uncoded_block[234];
  wire _65296 = _65294 ^ _65295;
  wire _65297 = _65293 ^ _65296;
  wire _65298 = uncoded_block[240] ^ uncoded_block[298];
  wire _65299 = uncoded_block[326] ^ uncoded_block[374];
  wire _65300 = _65298 ^ _65299;
  wire _65301 = uncoded_block[418] ^ uncoded_block[439];
  wire _65302 = uncoded_block[458] ^ uncoded_block[474];
  wire _65303 = _65301 ^ _65302;
  wire _65304 = _65300 ^ _65303;
  wire _65305 = _65297 ^ _65304;
  wire _65306 = uncoded_block[550] ^ uncoded_block[590];
  wire _65307 = uncoded_block[606] ^ uncoded_block[617];
  wire _65308 = _65306 ^ _65307;
  wire _65309 = uncoded_block[636] ^ uncoded_block[685];
  wire _65310 = uncoded_block[702] ^ uncoded_block[734];
  wire _65311 = _65309 ^ _65310;
  wire _65312 = _65308 ^ _65311;
  wire _65313 = uncoded_block[767] ^ uncoded_block[803];
  wire _65314 = uncoded_block[814] ^ uncoded_block[840];
  wire _65315 = _65313 ^ _65314;
  wire _65316 = uncoded_block[854] ^ uncoded_block[897];
  wire _65317 = uncoded_block[919] ^ uncoded_block[961];
  wire _65318 = _65316 ^ _65317;
  wire _65319 = _65315 ^ _65318;
  wire _65320 = _65312 ^ _65319;
  wire _65321 = _65305 ^ _65320;
  wire _65322 = uncoded_block[963] ^ uncoded_block[1035];
  wire _65323 = uncoded_block[1040] ^ uncoded_block[1086];
  wire _65324 = _65322 ^ _65323;
  wire _65325 = uncoded_block[1094] ^ uncoded_block[1127];
  wire _65326 = uncoded_block[1150] ^ uncoded_block[1181];
  wire _65327 = _65325 ^ _65326;
  wire _65328 = _65324 ^ _65327;
  wire _65329 = uncoded_block[1263] ^ uncoded_block[1325];
  wire _65330 = _65329 ^ _49595;
  wire _65331 = uncoded_block[1378] ^ uncoded_block[1390];
  wire _65332 = _65331 ^ _60896;
  wire _65333 = _65330 ^ _65332;
  wire _65334 = _65328 ^ _65333;
  wire _65335 = uncoded_block[1497] ^ uncoded_block[1517];
  wire _65336 = uncoded_block[1521] ^ uncoded_block[1554];
  wire _65337 = _65335 ^ _65336;
  wire _65338 = uncoded_block[1556] ^ uncoded_block[1564];
  wire _65339 = _65338 ^ _16515;
  wire _65340 = _65337 ^ _65339;
  wire _65341 = _6685 ^ _62342;
  wire _65342 = _65341 ^ uncoded_block[1722];
  wire _65343 = _65340 ^ _65342;
  wire _65344 = _65334 ^ _65343;
  wire _65345 = _65321 ^ _65344;
  wire _65346 = uncoded_block[38] ^ uncoded_block[63];
  wire _65347 = _2459 ^ _65346;
  wire _65348 = _41044 ^ _62463;
  wire _65349 = _65347 ^ _65348;
  wire _65350 = uncoded_block[162] ^ uncoded_block[181];
  wire _65351 = uncoded_block[184] ^ uncoded_block[190];
  wire _65352 = _65350 ^ _65351;
  wire _65353 = uncoded_block[254] ^ uncoded_block[291];
  wire _65354 = _968 ^ _65353;
  wire _65355 = _65352 ^ _65354;
  wire _65356 = _65349 ^ _65355;
  wire _65357 = uncoded_block[339] ^ uncoded_block[352];
  wire _65358 = _5525 ^ _65357;
  wire _65359 = uncoded_block[380] ^ uncoded_block[420];
  wire _65360 = uncoded_block[421] ^ uncoded_block[443];
  wire _65361 = _65359 ^ _65360;
  wire _65362 = _65358 ^ _65361;
  wire _65363 = uncoded_block[476] ^ uncoded_block[520];
  wire _65364 = _62492 ^ _65363;
  wire _65365 = _65364 ^ _62501;
  wire _65366 = _65362 ^ _65365;
  wire _65367 = _65356 ^ _65366;
  wire _65368 = uncoded_block[611] ^ uncoded_block[618];
  wire _65369 = uncoded_block[621] ^ uncoded_block[647];
  wire _65370 = _65368 ^ _65369;
  wire _65371 = uncoded_block[678] ^ uncoded_block[699];
  wire _65372 = uncoded_block[715] ^ uncoded_block[729];
  wire _65373 = _65371 ^ _65372;
  wire _65374 = _65370 ^ _65373;
  wire _65375 = uncoded_block[732] ^ uncoded_block[770];
  wire _65376 = _65375 ^ _5035;
  wire _65377 = uncoded_block[814] ^ uncoded_block[863];
  wire _65378 = _65377 ^ _417;
  wire _65379 = _65376 ^ _65378;
  wire _65380 = _65374 ^ _65379;
  wire _65381 = uncoded_block[905] ^ uncoded_block[932];
  wire _65382 = uncoded_block[949] ^ uncoded_block[984];
  wire _65383 = _65381 ^ _65382;
  wire _65384 = uncoded_block[995] ^ uncoded_block[1031];
  wire _65385 = _65384 ^ _11116;
  wire _65386 = _65383 ^ _65385;
  wire _65387 = uncoded_block[1059] ^ uncoded_block[1086];
  wire _65388 = uncoded_block[1098] ^ uncoded_block[1119];
  wire _65389 = _65387 ^ _65388;
  wire _65390 = uncoded_block[1127] ^ uncoded_block[1145];
  wire _65391 = _65390 ^ _585;
  wire _65392 = _65389 ^ _65391;
  wire _65393 = _65386 ^ _65392;
  wire _65394 = _65380 ^ _65393;
  wire _65395 = _65367 ^ _65394;
  wire _65396 = uncoded_block[1189] ^ uncoded_block[1236];
  wire _65397 = _65396 ^ _62562;
  wire _65398 = uncoded_block[1307] ^ uncoded_block[1313];
  wire _65399 = uncoded_block[1346] ^ uncoded_block[1355];
  wire _65400 = _65398 ^ _65399;
  wire _65401 = _65397 ^ _65400;
  wire _65402 = uncoded_block[1406] ^ uncoded_block[1433];
  wire _65403 = uncoded_block[1444] ^ uncoded_block[1455];
  wire _65404 = _65402 ^ _65403;
  wire _65405 = uncoded_block[1457] ^ uncoded_block[1487];
  wire _65406 = uncoded_block[1507] ^ uncoded_block[1528];
  wire _65407 = _65405 ^ _65406;
  wire _65408 = _65404 ^ _65407;
  wire _65409 = _65401 ^ _65408;
  wire _65410 = _60436 ^ _62592;
  wire _65411 = uncoded_block[1623] ^ uncoded_block[1657];
  wire _65412 = _62595 ^ _65411;
  wire _65413 = _65410 ^ _65412;
  wire _65414 = uncoded_block[1665] ^ uncoded_block[1684];
  wire _65415 = _65414 ^ uncoded_block[1706];
  wire _65416 = _65413 ^ _65415;
  wire _65417 = _65409 ^ _65416;
  wire _65418 = _65395 ^ _65417;
  wire _65419 = uncoded_block[36] ^ uncoded_block[46];
  wire _65420 = uncoded_block[78] ^ uncoded_block[94];
  wire _65421 = _65419 ^ _65420;
  wire _65422 = uncoded_block[123] ^ uncoded_block[148];
  wire _65423 = _65422 ^ _30963;
  wire _65424 = _65421 ^ _65423;
  wire _65425 = uncoded_block[225] ^ uncoded_block[272];
  wire _65426 = uncoded_block[293] ^ uncoded_block[318];
  wire _65427 = _65425 ^ _65426;
  wire _65428 = uncoded_block[341] ^ uncoded_block[361];
  wire _65429 = uncoded_block[393] ^ uncoded_block[446];
  wire _65430 = _65428 ^ _65429;
  wire _65431 = _65427 ^ _65430;
  wire _65432 = _65424 ^ _65431;
  wire _65433 = uncoded_block[461] ^ uncoded_block[502];
  wire _65434 = uncoded_block[521] ^ uncoded_block[557];
  wire _65435 = _65433 ^ _65434;
  wire _65436 = uncoded_block[585] ^ uncoded_block[612];
  wire _65437 = uncoded_block[634] ^ uncoded_block[654];
  wire _65438 = _65436 ^ _65437;
  wire _65439 = _65435 ^ _65438;
  wire _65440 = uncoded_block[674] ^ uncoded_block[701];
  wire _65441 = uncoded_block[746] ^ uncoded_block[777];
  wire _65442 = _65440 ^ _65441;
  wire _65443 = uncoded_block[783] ^ uncoded_block[837];
  wire _65444 = uncoded_block[870] ^ uncoded_block[911];
  wire _65445 = _65443 ^ _65444;
  wire _65446 = _65442 ^ _65445;
  wire _65447 = _65439 ^ _65446;
  wire _65448 = _65432 ^ _65447;
  wire _65449 = uncoded_block[913] ^ uncoded_block[956];
  wire _65450 = uncoded_block[974] ^ uncoded_block[1008];
  wire _65451 = _65449 ^ _65450;
  wire _65452 = uncoded_block[1038] ^ uncoded_block[1061];
  wire _65453 = uncoded_block[1066] ^ uncoded_block[1122];
  wire _65454 = _65452 ^ _65453;
  wire _65455 = _65451 ^ _65454;
  wire _65456 = uncoded_block[1151] ^ uncoded_block[1182];
  wire _65457 = uncoded_block[1186] ^ uncoded_block[1244];
  wire _65458 = _65456 ^ _65457;
  wire _65459 = uncoded_block[1262] ^ uncoded_block[1310];
  wire _65460 = uncoded_block[1349] ^ uncoded_block[1371];
  wire _65461 = _65459 ^ _65460;
  wire _65462 = _65458 ^ _65461;
  wire _65463 = _65455 ^ _65462;
  wire _65464 = uncoded_block[1401] ^ uncoded_block[1428];
  wire _65465 = _65464 ^ _59201;
  wire _65466 = uncoded_block[1500] ^ uncoded_block[1527];
  wire _65467 = _3884 ^ _65466;
  wire _65468 = _65465 ^ _65467;
  wire _65469 = uncoded_block[1537] ^ uncoded_block[1632];
  wire _65470 = uncoded_block[1635] ^ uncoded_block[1698];
  wire _65471 = _65469 ^ _65470;
  wire _65472 = _65471 ^ uncoded_block[1699];
  wire _65473 = _65468 ^ _65472;
  wire _65474 = _65463 ^ _65473;
  wire _65475 = _65448 ^ _65474;
  wire _65476 = uncoded_block[3] ^ uncoded_block[36];
  wire _65477 = uncoded_block[41] ^ uncoded_block[78];
  wire _65478 = _65476 ^ _65477;
  wire _65479 = uncoded_block[86] ^ uncoded_block[106];
  wire _65480 = _65479 ^ _10821;
  wire _65481 = _65478 ^ _65480;
  wire _65482 = uncoded_block[146] ^ uncoded_block[174];
  wire _65483 = _65482 ^ _11943;
  wire _65484 = uncoded_block[225] ^ uncoded_block[265];
  wire _65485 = uncoded_block[270] ^ uncoded_block[293];
  wire _65486 = _65484 ^ _65485;
  wire _65487 = _65483 ^ _65486;
  wire _65488 = _65481 ^ _65487;
  wire _65489 = _61273 ^ _62010;
  wire _65490 = uncoded_block[384] ^ uncoded_block[393];
  wire _65491 = uncoded_block[408] ^ uncoded_block[437];
  wire _65492 = _65490 ^ _65491;
  wire _65493 = _65489 ^ _65492;
  wire _65494 = uncoded_block[481] ^ uncoded_block[509];
  wire _65495 = _13127 ^ _65494;
  wire _65496 = uncoded_block[571] ^ uncoded_block[585];
  wire _65497 = _61290 ^ _65496;
  wire _65498 = _65495 ^ _65497;
  wire _65499 = _65493 ^ _65498;
  wire _65500 = _65488 ^ _65499;
  wire _65501 = uncoded_block[588] ^ uncoded_block[619];
  wire _65502 = _65501 ^ _60523;
  wire _65503 = uncoded_block[674] ^ uncoded_block[699];
  wire _65504 = uncoded_block[710] ^ uncoded_block[740];
  wire _65505 = _65503 ^ _65504;
  wire _65506 = _65502 ^ _65505;
  wire _65507 = uncoded_block[746] ^ uncoded_block[761];
  wire _65508 = _65507 ^ _13768;
  wire _65509 = uncoded_block[810] ^ uncoded_block[835];
  wire _65510 = _65509 ^ _9938;
  wire _65511 = _65508 ^ _65510;
  wire _65512 = _65506 ^ _65511;
  wire _65513 = uncoded_block[889] ^ uncoded_block[912];
  wire _65514 = uncoded_block[913] ^ uncoded_block[974];
  wire _65515 = _65513 ^ _65514;
  wire _65516 = _4402 ^ _5801;
  wire _65517 = _65515 ^ _65516;
  wire _65518 = uncoded_block[1041] ^ uncoded_block[1061];
  wire _65519 = _65518 ^ _61337;
  wire _65520 = uncoded_block[1122] ^ uncoded_block[1143];
  wire _65521 = uncoded_block[1177] ^ uncoded_block[1186];
  wire _65522 = _65520 ^ _65521;
  wire _65523 = _65519 ^ _65522;
  wire _65524 = _65517 ^ _65523;
  wire _65525 = _65512 ^ _65524;
  wire _65526 = _65500 ^ _65525;
  wire _65527 = uncoded_block[1188] ^ uncoded_block[1257];
  wire _65528 = uncoded_block[1262] ^ uncoded_block[1268];
  wire _65529 = _65527 ^ _65528;
  wire _65530 = _61356 ^ _61360;
  wire _65531 = _65529 ^ _65530;
  wire _65532 = uncoded_block[1371] ^ uncoded_block[1420];
  wire _65533 = _65532 ^ _2311;
  wire _65534 = uncoded_block[1448] ^ uncoded_block[1460];
  wire _65535 = _65534 ^ _65019;
  wire _65536 = _65533 ^ _65535;
  wire _65537 = _65531 ^ _65536;
  wire _65538 = uncoded_block[1481] ^ uncoded_block[1513];
  wire _65539 = _65538 ^ _61378;
  wire _65540 = uncoded_block[1547] ^ uncoded_block[1609];
  wire _65541 = _65540 ^ _61384;
  wire _65542 = _65539 ^ _65541;
  wire _65543 = _2430 ^ uncoded_block[1715];
  wire _65544 = _65542 ^ _65543;
  wire _65545 = _65537 ^ _65544;
  wire _65546 = _65526 ^ _65545;
  wire _65547 = uncoded_block[7] ^ uncoded_block[87];
  wire _65548 = uncoded_block[97] ^ uncoded_block[111];
  wire _65549 = _65547 ^ _65548;
  wire _65550 = uncoded_block[157] ^ uncoded_block[198];
  wire _65551 = uncoded_block[222] ^ uncoded_block[237];
  wire _65552 = _65550 ^ _65551;
  wire _65553 = _65549 ^ _65552;
  wire _65554 = uncoded_block[263] ^ uncoded_block[283];
  wire _65555 = uncoded_block[323] ^ uncoded_block[359];
  wire _65556 = _65554 ^ _65555;
  wire _65557 = uncoded_block[371] ^ uncoded_block[437];
  wire _65558 = _65557 ^ _58123;
  wire _65559 = _65556 ^ _65558;
  wire _65560 = _65553 ^ _65559;
  wire _65561 = uncoded_block[471] ^ uncoded_block[512];
  wire _65562 = uncoded_block[547] ^ uncoded_block[595];
  wire _65563 = _65561 ^ _65562;
  wire _65564 = uncoded_block[603] ^ uncoded_block[619];
  wire _65565 = uncoded_block[633] ^ uncoded_block[682];
  wire _65566 = _65564 ^ _65565;
  wire _65567 = _65563 ^ _65566;
  wire _65568 = uncoded_block[709] ^ uncoded_block[751];
  wire _65569 = uncoded_block[764] ^ uncoded_block[811];
  wire _65570 = _65568 ^ _65569;
  wire _65571 = uncoded_block[828] ^ uncoded_block[851];
  wire _65572 = uncoded_block[865] ^ uncoded_block[894];
  wire _65573 = _65571 ^ _65572;
  wire _65574 = _65570 ^ _65573;
  wire _65575 = _65567 ^ _65574;
  wire _65576 = _65560 ^ _65575;
  wire _65577 = uncoded_block[925] ^ uncoded_block[958];
  wire _65578 = uncoded_block[982] ^ uncoded_block[1031];
  wire _65579 = _65577 ^ _65578;
  wire _65580 = uncoded_block[1033] ^ uncoded_block[1091];
  wire _65581 = uncoded_block[1098] ^ uncoded_block[1124];
  wire _65582 = _65580 ^ _65581;
  wire _65583 = _65579 ^ _65582;
  wire _65584 = uncoded_block[1126] ^ uncoded_block[1167];
  wire _65585 = uncoded_block[1178] ^ uncoded_block[1184];
  wire _65586 = _65584 ^ _65585;
  wire _65587 = uncoded_block[1301] ^ uncoded_block[1324];
  wire _65588 = _63926 ^ _65587;
  wire _65589 = _65586 ^ _65588;
  wire _65590 = _65583 ^ _65589;
  wire _65591 = uncoded_block[1331] ^ uncoded_block[1376];
  wire _65592 = uncoded_block[1396] ^ uncoded_block[1423];
  wire _65593 = _65591 ^ _65592;
  wire _65594 = uncoded_block[1562] ^ uncoded_block[1571];
  wire _65595 = _65594 ^ _15031;
  wire _65596 = _65593 ^ _65595;
  wire _65597 = uncoded_block[1613] ^ uncoded_block[1628];
  wire _65598 = uncoded_block[1708] ^ uncoded_block[1716];
  wire _65599 = _65597 ^ _65598;
  wire _65600 = _65599 ^ uncoded_block[1720];
  wire _65601 = _65596 ^ _65600;
  wire _65602 = _65590 ^ _65601;
  wire _65603 = _65576 ^ _65602;
  wire _65604 = uncoded_block[8] ^ uncoded_block[24];
  wire _65605 = uncoded_block[77] ^ uncoded_block[102];
  wire _65606 = _65604 ^ _65605;
  wire _65607 = uncoded_block[112] ^ uncoded_block[163];
  wire _65608 = uncoded_block[178] ^ uncoded_block[224];
  wire _65609 = _65607 ^ _65608;
  wire _65610 = _65606 ^ _65609;
  wire _65611 = uncoded_block[230] ^ uncoded_block[235];
  wire _65612 = uncoded_block[293] ^ uncoded_block[310];
  wire _65613 = _65611 ^ _65612;
  wire _65614 = uncoded_block[339] ^ uncoded_block[382];
  wire _65615 = _65614 ^ _13650;
  wire _65616 = _65613 ^ _65615;
  wire _65617 = _65610 ^ _65616;
  wire _65618 = uncoded_block[470] ^ uncoded_block[497];
  wire _65619 = uncoded_block[506] ^ uncoded_block[544];
  wire _65620 = _65618 ^ _65619;
  wire _65621 = uncoded_block[640] ^ uncoded_block[646];
  wire _65622 = _6947 ^ _65621;
  wire _65623 = _65620 ^ _65622;
  wire _65624 = uncoded_block[686] ^ uncoded_block[697];
  wire _65625 = uncoded_block[727] ^ uncoded_block[764];
  wire _65626 = _65624 ^ _65625;
  wire _65627 = uncoded_block[789] ^ uncoded_block[823];
  wire _65628 = _65627 ^ _64536;
  wire _65629 = _65626 ^ _65628;
  wire _65630 = _65623 ^ _65629;
  wire _65631 = _65617 ^ _65630;
  wire _65632 = uncoded_block[890] ^ uncoded_block[918];
  wire _65633 = uncoded_block[947] ^ uncoded_block[966];
  wire _65634 = _65632 ^ _65633;
  wire _65635 = uncoded_block[1003] ^ uncoded_block[1012];
  wire _65636 = uncoded_block[1027] ^ uncoded_block[1063];
  wire _65637 = _65635 ^ _65636;
  wire _65638 = _65634 ^ _65637;
  wire _65639 = uncoded_block[1078] ^ uncoded_block[1137];
  wire _65640 = uncoded_block[1144] ^ uncoded_block[1181];
  wire _65641 = _65639 ^ _65640;
  wire _65642 = uncoded_block[1208] ^ uncoded_block[1218];
  wire _65643 = uncoded_block[1265] ^ uncoded_block[1326];
  wire _65644 = _65642 ^ _65643;
  wire _65645 = _65641 ^ _65644;
  wire _65646 = _65638 ^ _65645;
  wire _65647 = uncoded_block[1337] ^ uncoded_block[1373];
  wire _65648 = uncoded_block[1407] ^ uncoded_block[1468];
  wire _65649 = _65647 ^ _65648;
  wire _65650 = uncoded_block[1475] ^ uncoded_block[1520];
  wire _65651 = uncoded_block[1546] ^ uncoded_block[1578];
  wire _65652 = _65650 ^ _65651;
  wire _65653 = _65649 ^ _65652;
  wire _65654 = uncoded_block[1592] ^ uncoded_block[1621];
  wire _65655 = uncoded_block[1642] ^ uncoded_block[1660];
  wire _65656 = _65654 ^ _65655;
  wire _65657 = _65656 ^ uncoded_block[1681];
  wire _65658 = _65653 ^ _65657;
  wire _65659 = _65646 ^ _65658;
  wire _65660 = _65631 ^ _65659;
  wire _65661 = uncoded_block[12] ^ uncoded_block[29];
  wire _65662 = uncoded_block[45] ^ uncoded_block[75];
  wire _65663 = _65661 ^ _65662;
  wire _65664 = uncoded_block[126] ^ uncoded_block[134];
  wire _65665 = _61771 ^ _65664;
  wire _65666 = _65663 ^ _65665;
  wire _65667 = uncoded_block[148] ^ uncoded_block[198];
  wire _65668 = _65667 ^ _14099;
  wire _65669 = uncoded_block[227] ^ uncoded_block[245];
  wire _65670 = uncoded_block[262] ^ uncoded_block[282];
  wire _65671 = _65669 ^ _65670;
  wire _65672 = _65668 ^ _65671;
  wire _65673 = _65666 ^ _65672;
  wire _65674 = uncoded_block[300] ^ uncoded_block[329];
  wire _65675 = uncoded_block[339] ^ uncoded_block[351];
  wire _65676 = _65674 ^ _65675;
  wire _65677 = uncoded_block[387] ^ uncoded_block[406];
  wire _65678 = uncoded_block[408] ^ uncoded_block[414];
  wire _65679 = _65677 ^ _65678;
  wire _65680 = _65676 ^ _65679;
  wire _65681 = uncoded_block[448] ^ uncoded_block[485];
  wire _65682 = uncoded_block[501] ^ uncoded_block[523];
  wire _65683 = _65681 ^ _65682;
  wire _65684 = uncoded_block[524] ^ uncoded_block[554];
  wire _65685 = uncoded_block[570] ^ uncoded_block[574];
  wire _65686 = _65684 ^ _65685;
  wire _65687 = _65683 ^ _65686;
  wire _65688 = _65680 ^ _65687;
  wire _65689 = _65673 ^ _65688;
  wire _65690 = uncoded_block[611] ^ uncoded_block[627];
  wire _65691 = uncoded_block[628] ^ uncoded_block[639];
  wire _65692 = _65690 ^ _65691;
  wire _65693 = uncoded_block[681] ^ uncoded_block[704];
  wire _65694 = uncoded_block[711] ^ uncoded_block[747];
  wire _65695 = _65693 ^ _65694;
  wire _65696 = _65692 ^ _65695;
  wire _65697 = uncoded_block[760] ^ uncoded_block[776];
  wire _65698 = _65697 ^ _3576;
  wire _65699 = uncoded_block[820] ^ uncoded_block[849];
  wire _65700 = _65699 ^ _47464;
  wire _65701 = _65698 ^ _65700;
  wire _65702 = _65696 ^ _65701;
  wire _65703 = uncoded_block[919] ^ uncoded_block[941];
  wire _65704 = _65703 ^ _21187;
  wire _65705 = uncoded_block[953] ^ uncoded_block[961];
  wire _65706 = _65705 ^ _47133;
  wire _65707 = _65704 ^ _65706;
  wire _65708 = uncoded_block[1044] ^ uncoded_block[1061];
  wire _65709 = uncoded_block[1078] ^ uncoded_block[1122];
  wire _65710 = _65708 ^ _65709;
  wire _65711 = uncoded_block[1129] ^ uncoded_block[1139];
  wire _65712 = uncoded_block[1194] ^ uncoded_block[1204];
  wire _65713 = _65711 ^ _65712;
  wire _65714 = _65710 ^ _65713;
  wire _65715 = _65707 ^ _65714;
  wire _65716 = _65702 ^ _65715;
  wire _65717 = _65689 ^ _65716;
  wire _65718 = uncoded_block[1210] ^ uncoded_block[1224];
  wire _65719 = _65718 ^ _14412;
  wire _65720 = uncoded_block[1266] ^ uncoded_block[1299];
  wire _65721 = uncoded_block[1323] ^ uncoded_block[1332];
  wire _65722 = _65720 ^ _65721;
  wire _65723 = _65719 ^ _65722;
  wire _65724 = _20329 ^ _11782;
  wire _65725 = uncoded_block[1446] ^ uncoded_block[1495];
  wire _65726 = uncoded_block[1508] ^ uncoded_block[1532];
  wire _65727 = _65725 ^ _65726;
  wire _65728 = _65724 ^ _65727;
  wire _65729 = _65723 ^ _65728;
  wire _65730 = uncoded_block[1542] ^ uncoded_block[1572];
  wire _65731 = uncoded_block[1576] ^ uncoded_block[1602];
  wire _65732 = _65730 ^ _65731;
  wire _65733 = uncoded_block[1606] ^ uncoded_block[1613];
  wire _65734 = uncoded_block[1628] ^ uncoded_block[1639];
  wire _65735 = _65733 ^ _65734;
  wire _65736 = _65732 ^ _65735;
  wire _65737 = uncoded_block[1667] ^ uncoded_block[1685];
  wire _65738 = _65737 ^ uncoded_block[1707];
  wire _65739 = _65736 ^ _65738;
  wire _65740 = _65729 ^ _65739;
  wire _65741 = _65717 ^ _65740;
  wire _65742 = uncoded_block[2] ^ uncoded_block[13];
  wire _65743 = _65742 ^ _1691;
  wire _65744 = _65743 ^ _63170;
  wire _65745 = uncoded_block[69] ^ uncoded_block[103];
  wire _65746 = uncoded_block[111] ^ uncoded_block[133];
  wire _65747 = _65745 ^ _65746;
  wire _65748 = uncoded_block[140] ^ uncoded_block[145];
  wire _65749 = _65748 ^ _57822;
  wire _65750 = _65747 ^ _65749;
  wire _65751 = _65744 ^ _65750;
  wire _65752 = uncoded_block[178] ^ uncoded_block[185];
  wire _65753 = _65752 ^ _53080;
  wire _65754 = uncoded_block[195] ^ uncoded_block[211];
  wire _65755 = uncoded_block[226] ^ uncoded_block[233];
  wire _65756 = _65754 ^ _65755;
  wire _65757 = _65753 ^ _65756;
  wire _65758 = uncoded_block[242] ^ uncoded_block[258];
  wire _65759 = uncoded_block[265] ^ uncoded_block[277];
  wire _65760 = _65758 ^ _65759;
  wire _65761 = uncoded_block[280] ^ uncoded_block[290];
  wire _65762 = uncoded_block[314] ^ uncoded_block[324];
  wire _65763 = _65761 ^ _65762;
  wire _65764 = _65760 ^ _65763;
  wire _65765 = _65757 ^ _65764;
  wire _65766 = _65751 ^ _65765;
  wire _65767 = uncoded_block[351] ^ uncoded_block[358];
  wire _65768 = uncoded_block[368] ^ uncoded_block[378];
  wire _65769 = _65767 ^ _65768;
  wire _65770 = uncoded_block[417] ^ uncoded_block[432];
  wire _65771 = _31005 ^ _65770;
  wire _65772 = _65769 ^ _65771;
  wire _65773 = _24711 ^ _32709;
  wire _65774 = uncoded_block[469] ^ uncoded_block[481];
  wire _65775 = uncoded_block[489] ^ uncoded_block[501];
  wire _65776 = _65774 ^ _65775;
  wire _65777 = _65773 ^ _65776;
  wire _65778 = _65772 ^ _65777;
  wire _65779 = uncoded_block[516] ^ uncoded_block[541];
  wire _65780 = _1893 ^ _65779;
  wire _65781 = uncoded_block[546] ^ uncoded_block[555];
  wire _65782 = uncoded_block[570] ^ uncoded_block[587];
  wire _65783 = _65781 ^ _65782;
  wire _65784 = _65780 ^ _65783;
  wire _65785 = _7556 ^ _18232;
  wire _65786 = uncoded_block[620] ^ uncoded_block[634];
  wire _65787 = _6959 ^ _65786;
  wire _65788 = _65785 ^ _65787;
  wire _65789 = _65784 ^ _65788;
  wire _65790 = _65778 ^ _65789;
  wire _65791 = _65766 ^ _65790;
  wire _65792 = uncoded_block[677] ^ uncoded_block[691];
  wire _65793 = _65621 ^ _65792;
  wire _65794 = uncoded_block[699] ^ uncoded_block[707];
  wire _65795 = uncoded_block[714] ^ uncoded_block[718];
  wire _65796 = _65794 ^ _65795;
  wire _65797 = _65793 ^ _65796;
  wire _65798 = uncoded_block[726] ^ uncoded_block[746];
  wire _65799 = uncoded_block[748] ^ uncoded_block[772];
  wire _65800 = _65798 ^ _65799;
  wire _65801 = uncoded_block[807] ^ uncoded_block[813];
  wire _65802 = _33218 ^ _65801;
  wire _65803 = _65800 ^ _65802;
  wire _65804 = _65797 ^ _65803;
  wire _65805 = uncoded_block[831] ^ uncoded_block[863];
  wire _65806 = _63270 ^ _65805;
  wire _65807 = uncoded_block[887] ^ uncoded_block[897];
  wire _65808 = _16815 ^ _65807;
  wire _65809 = _65806 ^ _65808;
  wire _65810 = uncoded_block[906] ^ uncoded_block[931];
  wire _65811 = _45355 ^ _65810;
  wire _65812 = uncoded_block[958] ^ uncoded_block[972];
  wire _65813 = _65812 ^ _8287;
  wire _65814 = _65811 ^ _65813;
  wire _65815 = _65809 ^ _65814;
  wire _65816 = _65804 ^ _65815;
  wire _65817 = uncoded_block[988] ^ uncoded_block[994];
  wire _65818 = uncoded_block[1018] ^ uncoded_block[1035];
  wire _65819 = _65817 ^ _65818;
  wire _65820 = _59138 ^ _6485;
  wire _65821 = _65819 ^ _65820;
  wire _65822 = uncoded_block[1075] ^ uncoded_block[1096];
  wire _65823 = uncoded_block[1098] ^ uncoded_block[1109];
  wire _65824 = _65822 ^ _65823;
  wire _65825 = uncoded_block[1137] ^ uncoded_block[1144];
  wire _65826 = uncoded_block[1158] ^ uncoded_block[1165];
  wire _65827 = _65825 ^ _65826;
  wire _65828 = _65824 ^ _65827;
  wire _65829 = _65821 ^ _65828;
  wire _65830 = _2192 ^ _7159;
  wire _65831 = uncoded_block[1198] ^ uncoded_block[1222];
  wire _65832 = _65831 ^ _64108;
  wire _65833 = _65830 ^ _65832;
  wire _65834 = uncoded_block[1270] ^ uncoded_block[1284];
  wire _65835 = _5229 ^ _65834;
  wire _65836 = uncoded_block[1298] ^ uncoded_block[1311];
  wire _65837 = uncoded_block[1313] ^ uncoded_block[1322];
  wire _65838 = _65836 ^ _65837;
  wire _65839 = _65835 ^ _65838;
  wire _65840 = _65833 ^ _65839;
  wire _65841 = _65829 ^ _65840;
  wire _65842 = _65816 ^ _65841;
  wire _65843 = _65791 ^ _65842;
  wire _65844 = uncoded_block[1330] ^ uncoded_block[1345];
  wire _65845 = uncoded_block[1357] ^ uncoded_block[1366];
  wire _65846 = _65844 ^ _65845;
  wire _65847 = _5281 ^ _3061;
  wire _65848 = _65846 ^ _65847;
  wire _65849 = uncoded_block[1404] ^ uncoded_block[1413];
  wire _65850 = _65849 ^ _716;
  wire _65851 = uncoded_block[1478] ^ uncoded_block[1502];
  wire _65852 = uncoded_block[1510] ^ uncoded_block[1524];
  wire _65853 = _65851 ^ _65852;
  wire _65854 = _65850 ^ _65853;
  wire _65855 = _65848 ^ _65854;
  wire _65856 = uncoded_block[1540] ^ uncoded_block[1552];
  wire _65857 = _60098 ^ _65856;
  wire _65858 = uncoded_block[1565] ^ uncoded_block[1575];
  wire _65859 = uncoded_block[1576] ^ uncoded_block[1595];
  wire _65860 = _65858 ^ _65859;
  wire _65861 = _65857 ^ _65860;
  wire _65862 = _54551 ^ _7300;
  wire _65863 = uncoded_block[1631] ^ uncoded_block[1660];
  wire _65864 = _4667 ^ _65863;
  wire _65865 = _65862 ^ _65864;
  wire _65866 = _65861 ^ _65865;
  wire _65867 = _65855 ^ _65866;
  wire _65868 = uncoded_block[1661] ^ uncoded_block[1683];
  wire _65869 = _65868 ^ _13519;
  wire _65870 = uncoded_block[1697] ^ uncoded_block[1706];
  wire _65871 = _65870 ^ uncoded_block[1709];
  wire _65872 = _65869 ^ _65871;
  wire _65873 = _65867 ^ _65872;
  wire _65874 = _65843 ^ _65873;
  wire _65875 = uncoded_block[0] ^ uncoded_block[19];
  wire _65876 = uncoded_block[96] ^ uncoded_block[106];
  wire _65877 = _65875 ^ _65876;
  wire _65878 = uncoded_block[193] ^ uncoded_block[223];
  wire _65879 = _61411 ^ _65878;
  wire _65880 = _65877 ^ _65879;
  wire _65881 = uncoded_block[226] ^ uncoded_block[249];
  wire _65882 = uncoded_block[318] ^ uncoded_block[354];
  wire _65883 = _65881 ^ _65882;
  wire _65884 = uncoded_block[377] ^ uncoded_block[439];
  wire _65885 = uncoded_block[444] ^ uncoded_block[484];
  wire _65886 = _65884 ^ _65885;
  wire _65887 = _65883 ^ _65886;
  wire _65888 = _65880 ^ _65887;
  wire _65889 = uncoded_block[487] ^ uncoded_block[545];
  wire _65890 = uncoded_block[558] ^ uncoded_block[590];
  wire _65891 = _65889 ^ _65890;
  wire _65892 = uncoded_block[603] ^ uncoded_block[629];
  wire _65893 = uncoded_block[658] ^ uncoded_block[673];
  wire _65894 = _65892 ^ _65893;
  wire _65895 = _65891 ^ _65894;
  wire _65896 = uncoded_block[689] ^ uncoded_block[726];
  wire _65897 = uncoded_block[757] ^ uncoded_block[783];
  wire _65898 = _65896 ^ _65897;
  wire _65899 = uncoded_block[796] ^ uncoded_block[850];
  wire _65900 = uncoded_block[867] ^ uncoded_block[896];
  wire _65901 = _65899 ^ _65900;
  wire _65902 = _65898 ^ _65901;
  wire _65903 = _65895 ^ _65902;
  wire _65904 = _65888 ^ _65903;
  wire _65905 = uncoded_block[909] ^ uncoded_block[973];
  wire _65906 = _65905 ^ _22585;
  wire _65907 = uncoded_block[1055] ^ uncoded_block[1080];
  wire _65908 = uncoded_block[1089] ^ uncoded_block[1125];
  wire _65909 = _65907 ^ _65908;
  wire _65910 = _65906 ^ _65909;
  wire _65911 = uncoded_block[1176] ^ uncoded_block[1205];
  wire _65912 = uncoded_block[1248] ^ uncoded_block[1305];
  wire _65913 = _65911 ^ _65912;
  wire _65914 = _61525 ^ _1523;
  wire _65915 = _65913 ^ _65914;
  wire _65916 = _65910 ^ _65915;
  wire _65917 = uncoded_block[1426] ^ uncoded_block[1450];
  wire _65918 = _65917 ^ _10699;
  wire _65919 = uncoded_block[1494] ^ uncoded_block[1512];
  wire _65920 = _65919 ^ _61543;
  wire _65921 = _65918 ^ _65920;
  wire _65922 = uncoded_block[1558] ^ uncoded_block[1568];
  wire _65923 = uncoded_block[1610] ^ uncoded_block[1648];
  wire _65924 = _65922 ^ _65923;
  wire _65925 = _65924 ^ uncoded_block[1652];
  wire _65926 = _65921 ^ _65925;
  wire _65927 = _65916 ^ _65926;
  wire _65928 = _65904 ^ _65927;
  wire _65929 = uncoded_block[24] ^ uncoded_block[82];
  wire _65930 = _3995 ^ _65929;
  wire _65931 = _50735 ^ _2497;
  wire _65932 = _65930 ^ _65931;
  wire _65933 = uncoded_block[155] ^ uncoded_block[189];
  wire _65934 = _65933 ^ _956;
  wire _65935 = uncoded_block[225] ^ uncoded_block[267];
  wire _65936 = uncoded_block[278] ^ uncoded_block[325];
  wire _65937 = _65935 ^ _65936;
  wire _65938 = _65934 ^ _65937;
  wire _65939 = _65932 ^ _65938;
  wire _65940 = _1819 ^ _1826;
  wire _65941 = uncoded_block[345] ^ uncoded_block[435];
  wire _65942 = _65941 ^ _9275;
  wire _65943 = _65940 ^ _65942;
  wire _65944 = uncoded_block[454] ^ uncoded_block[503];
  wire _65945 = uncoded_block[504] ^ uncoded_block[535];
  wire _65946 = _65944 ^ _65945;
  wire _65947 = uncoded_block[536] ^ uncoded_block[556];
  wire _65948 = _65947 ^ _4234;
  wire _65949 = _65946 ^ _65948;
  wire _65950 = _65943 ^ _65949;
  wire _65951 = _65939 ^ _65950;
  wire _65952 = uncoded_block[603] ^ uncoded_block[623];
  wire _65953 = _65952 ^ _1161;
  wire _65954 = uncoded_block[688] ^ uncoded_block[709];
  wire _65955 = uncoded_block[710] ^ uncoded_block[735];
  wire _65956 = _65954 ^ _65955;
  wire _65957 = _65953 ^ _65956;
  wire _65958 = uncoded_block[736] ^ uncoded_block[744];
  wire _65959 = uncoded_block[790] ^ uncoded_block[815];
  wire _65960 = _65958 ^ _65959;
  wire _65961 = uncoded_block[816] ^ uncoded_block[842];
  wire _65962 = _65961 ^ _1257;
  wire _65963 = _65960 ^ _65962;
  wire _65964 = _65957 ^ _65963;
  wire _65965 = uncoded_block[887] ^ uncoded_block[908];
  wire _65966 = uncoded_block[909] ^ uncoded_block[934];
  wire _65967 = _65965 ^ _65966;
  wire _65968 = uncoded_block[977] ^ uncoded_block[1005];
  wire _65969 = _3657 ^ _65968;
  wire _65970 = _65967 ^ _65969;
  wire _65971 = _3708 ^ _14380;
  wire _65972 = uncoded_block[1148] ^ uncoded_block[1164];
  wire _65973 = uncoded_block[1165] ^ uncoded_block[1172];
  wire _65974 = _65972 ^ _65973;
  wire _65975 = _65971 ^ _65974;
  wire _65976 = _65970 ^ _65975;
  wire _65977 = _65964 ^ _65976;
  wire _65978 = _65951 ^ _65977;
  wire _65979 = uncoded_block[1173] ^ uncoded_block[1192];
  wire _65980 = _65979 ^ _62755;
  wire _65981 = uncoded_block[1261] ^ uncoded_block[1293];
  wire _65982 = uncoded_block[1294] ^ uncoded_block[1333];
  wire _65983 = _65981 ^ _65982;
  wire _65984 = _65980 ^ _65983;
  wire _65985 = uncoded_block[1364] ^ uncoded_block[1395];
  wire _65986 = _1497 ^ _65985;
  wire _65987 = uncoded_block[1458] ^ uncoded_block[1494];
  wire _65988 = _2318 ^ _65987;
  wire _65989 = _65986 ^ _65988;
  wire _65990 = _65984 ^ _65989;
  wire _65991 = uncoded_block[1495] ^ uncoded_block[1507];
  wire _65992 = uncoded_block[1589] ^ uncoded_block[1606];
  wire _65993 = _65991 ^ _65992;
  wire _65994 = uncoded_block[1643] ^ uncoded_block[1659];
  wire _65995 = _14525 ^ _65994;
  wire _65996 = _65993 ^ _65995;
  wire _65997 = _65996 ^ uncoded_block[1704];
  wire _65998 = _65990 ^ _65997;
  wire _65999 = _65978 ^ _65998;
  wire _66000 = _3224 ^ _43266;
  wire _66001 = uncoded_block[70] ^ uncoded_block[82];
  wire _66002 = _66001 ^ _54;
  wire _66003 = _66000 ^ _66002;
  wire _66004 = uncoded_block[165] ^ uncoded_block[172];
  wire _66005 = uncoded_block[173] ^ uncoded_block[201];
  wire _66006 = _66004 ^ _66005;
  wire _66007 = uncoded_block[255] ^ uncoded_block[272];
  wire _66008 = uncoded_block[277] ^ uncoded_block[286];
  wire _66009 = _66007 ^ _66008;
  wire _66010 = _66006 ^ _66009;
  wire _66011 = _66003 ^ _66010;
  wire _66012 = uncoded_block[334] ^ uncoded_block[355];
  wire _66013 = _12515 ^ _66012;
  wire _66014 = uncoded_block[373] ^ uncoded_block[403];
  wire _66015 = _66014 ^ _15709;
  wire _66016 = _66013 ^ _66015;
  wire _66017 = uncoded_block[494] ^ uncoded_block[524];
  wire _66018 = _39197 ^ _66017;
  wire _66019 = uncoded_block[567] ^ uncoded_block[578];
  wire _66020 = _2687 ^ _66019;
  wire _66021 = _66018 ^ _66020;
  wire _66022 = _66016 ^ _66021;
  wire _66023 = _66011 ^ _66022;
  wire _66024 = uncoded_block[597] ^ uncoded_block[644];
  wire _66025 = uncoded_block[649] ^ uncoded_block[658];
  wire _66026 = _66024 ^ _66025;
  wire _66027 = uncoded_block[674] ^ uncoded_block[697];
  wire _66028 = uncoded_block[721] ^ uncoded_block[739];
  wire _66029 = _66027 ^ _66028;
  wire _66030 = _66026 ^ _66029;
  wire _66031 = uncoded_block[753] ^ uncoded_block[780];
  wire _66032 = uncoded_block[825] ^ uncoded_block[829];
  wire _66033 = _66031 ^ _66032;
  wire _66034 = uncoded_block[858] ^ uncoded_block[886];
  wire _66035 = uncoded_block[901] ^ uncoded_block[906];
  wire _66036 = _66034 ^ _66035;
  wire _66037 = _66033 ^ _66036;
  wire _66038 = _66030 ^ _66037;
  wire _66039 = uncoded_block[940] ^ uncoded_block[949];
  wire _66040 = uncoded_block[955] ^ uncoded_block[966];
  wire _66041 = _66039 ^ _66040;
  wire _66042 = uncoded_block[1081] ^ uncoded_block[1106];
  wire _66043 = _25768 ^ _66042;
  wire _66044 = _66041 ^ _66043;
  wire _66045 = uncoded_block[1139] ^ uncoded_block[1178];
  wire _66046 = _57147 ^ _66045;
  wire _66047 = uncoded_block[1179] ^ uncoded_block[1210];
  wire _66048 = uncoded_block[1221] ^ uncoded_block[1232];
  wire _66049 = _66047 ^ _66048;
  wire _66050 = _66046 ^ _66049;
  wire _66051 = _66044 ^ _66050;
  wire _66052 = _66038 ^ _66051;
  wire _66053 = _66023 ^ _66052;
  wire _66054 = uncoded_block[1240] ^ uncoded_block[1255];
  wire _66055 = uncoded_block[1281] ^ uncoded_block[1288];
  wire _66056 = _66054 ^ _66055;
  wire _66057 = uncoded_block[1292] ^ uncoded_block[1322];
  wire _66058 = uncoded_block[1364] ^ uncoded_block[1372];
  wire _66059 = _66057 ^ _66058;
  wire _66060 = _66056 ^ _66059;
  wire _66061 = _56893 ^ _59612;
  wire _66062 = uncoded_block[1421] ^ uncoded_block[1430];
  wire _66063 = uncoded_block[1465] ^ uncoded_block[1474];
  wire _66064 = _66062 ^ _66063;
  wire _66065 = _66061 ^ _66064;
  wire _66066 = _66060 ^ _66065;
  wire _66067 = uncoded_block[1506] ^ uncoded_block[1558];
  wire _66068 = _61949 ^ _66067;
  wire _66069 = uncoded_block[1587] ^ uncoded_block[1593];
  wire _66070 = uncoded_block[1618] ^ uncoded_block[1666];
  wire _66071 = _66069 ^ _66070;
  wire _66072 = _66068 ^ _66071;
  wire _66073 = _4698 ^ uncoded_block[1706];
  wire _66074 = _66072 ^ _66073;
  wire _66075 = _66066 ^ _66074;
  wire _66076 = _66053 ^ _66075;
  wire _66077 = uncoded_block[42] ^ uncoded_block[53];
  wire _66078 = uncoded_block[72] ^ uncoded_block[110];
  wire _66079 = _66077 ^ _66078;
  wire _66080 = uncoded_block[159] ^ uncoded_block[170];
  wire _66081 = uncoded_block[180] ^ uncoded_block[224];
  wire _66082 = _66080 ^ _66081;
  wire _66083 = _66079 ^ _66082;
  wire _66084 = uncoded_block[241] ^ uncoded_block[279];
  wire _66085 = uncoded_block[280] ^ uncoded_block[332];
  wire _66086 = _66084 ^ _66085;
  wire _66087 = uncoded_block[364] ^ uncoded_block[432];
  wire _66088 = uncoded_block[447] ^ uncoded_block[490];
  wire _66089 = _66087 ^ _66088;
  wire _66090 = _66086 ^ _66089;
  wire _66091 = _66083 ^ _66090;
  wire _66092 = uncoded_block[505] ^ uncoded_block[549];
  wire _66093 = uncoded_block[562] ^ uncoded_block[616];
  wire _66094 = _66092 ^ _66093;
  wire _66095 = uncoded_block[654] ^ uncoded_block[668];
  wire _66096 = uncoded_block[677] ^ uncoded_block[794];
  wire _66097 = _66095 ^ _66096;
  wire _66098 = _66094 ^ _66097;
  wire _66099 = uncoded_block[866] ^ uncoded_block[932];
  wire _66100 = uncoded_block[954] ^ uncoded_block[1026];
  wire _66101 = _66099 ^ _66100;
  wire _66102 = uncoded_block[1101] ^ uncoded_block[1158];
  wire _66103 = uncoded_block[1212] ^ uncoded_block[1272];
  wire _66104 = _66102 ^ _66103;
  wire _66105 = _66101 ^ _66104;
  wire _66106 = _66098 ^ _66105;
  wire _66107 = _66091 ^ _66106;
  wire _66108 = uncoded_block[1390] ^ uncoded_block[1421];
  wire _66109 = _65004 ^ _66108;
  wire _66110 = _66109 ^ _7257;
  wire _66111 = uncoded_block[1505] ^ uncoded_block[1509];
  wire _66112 = uncoded_block[1514] ^ uncoded_block[1519];
  wire _66113 = _66111 ^ _66112;
  wire _66114 = _36650 ^ _66113;
  wire _66115 = _66110 ^ _66114;
  wire _66116 = uncoded_block[1525] ^ uncoded_block[1532];
  wire _66117 = uncoded_block[1536] ^ uncoded_block[1552];
  wire _66118 = _66116 ^ _66117;
  wire _66119 = uncoded_block[1575] ^ uncoded_block[1601];
  wire _66120 = uncoded_block[1607] ^ uncoded_block[1628];
  wire _66121 = _66119 ^ _66120;
  wire _66122 = _66118 ^ _66121;
  wire _66123 = uncoded_block[1648] ^ uncoded_block[1677];
  wire _66124 = _66123 ^ _8526;
  wire _66125 = _66124 ^ uncoded_block[1718];
  wire _66126 = _66122 ^ _66125;
  wire _66127 = _66115 ^ _66126;
  wire _66128 = _66107 ^ _66127;
  wire _66129 = uncoded_block[7] ^ uncoded_block[27];
  wire _66130 = _66129 ^ _10234;
  wire _66131 = uncoded_block[54] ^ uncoded_block[70];
  wire _66132 = uncoded_block[73] ^ uncoded_block[98];
  wire _66133 = _66131 ^ _66132;
  wire _66134 = _66130 ^ _66133;
  wire _66135 = _64007 ^ _64009;
  wire _66136 = uncoded_block[185] ^ uncoded_block[199];
  wire _66137 = _66136 ^ _60761;
  wire _66138 = _66135 ^ _66137;
  wire _66139 = _66134 ^ _66138;
  wire _66140 = uncoded_block[242] ^ uncoded_block[256];
  wire _66141 = _40706 ^ _66140;
  wire _66142 = uncoded_block[305] ^ uncoded_block[328];
  wire _66143 = _4817 ^ _66142;
  wire _66144 = _66141 ^ _66143;
  wire _66145 = uncoded_block[337] ^ uncoded_block[349];
  wire _66146 = uncoded_block[369] ^ uncoded_block[382];
  wire _66147 = _66145 ^ _66146;
  wire _66148 = _10340 ^ _59717;
  wire _66149 = _66147 ^ _66148;
  wire _66150 = _66144 ^ _66149;
  wire _66151 = _66139 ^ _66150;
  wire _66152 = uncoded_block[476] ^ uncoded_block[495];
  wire _66153 = _66152 ^ _2667;
  wire _66154 = uncoded_block[523] ^ uncoded_block[572];
  wire _66155 = _17702 ^ _66154;
  wire _66156 = _66153 ^ _66155;
  wire _66157 = uncoded_block[600] ^ uncoded_block[625];
  wire _66158 = _64048 ^ _66157;
  wire _66159 = _302 ^ _3516;
  wire _66160 = _66158 ^ _66159;
  wire _66161 = _66156 ^ _66160;
  wire _66162 = uncoded_block[672] ^ uncoded_block[680];
  wire _66163 = uncoded_block[704] ^ uncoded_block[745];
  wire _66164 = _66162 ^ _66163;
  wire _66165 = uncoded_block[761] ^ uncoded_block[783];
  wire _66166 = _12663 ^ _66165;
  wire _66167 = _66164 ^ _66166;
  wire _66168 = uncoded_block[796] ^ uncoded_block[832];
  wire _66169 = _43031 ^ _66168;
  wire _66170 = uncoded_block[834] ^ uncoded_block[858];
  wire _66171 = uncoded_block[882] ^ uncoded_block[896];
  wire _66172 = _66170 ^ _66171;
  wire _66173 = _66169 ^ _66172;
  wire _66174 = _66167 ^ _66173;
  wire _66175 = _66161 ^ _66174;
  wire _66176 = _66151 ^ _66175;
  wire _66177 = uncoded_block[908] ^ uncoded_block[939];
  wire _66178 = _66177 ^ _64079;
  wire _66179 = uncoded_block[959] ^ uncoded_block[979];
  wire _66180 = uncoded_block[999] ^ uncoded_block[1012];
  wire _66181 = _66179 ^ _66180;
  wire _66182 = _66178 ^ _66181;
  wire _66183 = uncoded_block[1028] ^ uncoded_block[1042];
  wire _66184 = _66183 ^ _64093;
  wire _66185 = uncoded_block[1066] ^ uncoded_block[1077];
  wire _66186 = _66185 ^ _5166;
  wire _66187 = _66184 ^ _66186;
  wire _66188 = _66182 ^ _66187;
  wire _66189 = uncoded_block[1121] ^ uncoded_block[1149];
  wire _66190 = uncoded_block[1157] ^ uncoded_block[1186];
  wire _66191 = _66189 ^ _66190;
  wire _66192 = uncoded_block[1202] ^ uncoded_block[1227];
  wire _66193 = _66192 ^ _60875;
  wire _66194 = _66191 ^ _66193;
  wire _66195 = uncoded_block[1297] ^ uncoded_block[1321];
  wire _66196 = _64112 ^ _66195;
  wire _66197 = _63345 ^ _14447;
  wire _66198 = _66196 ^ _66197;
  wire _66199 = _66194 ^ _66198;
  wire _66200 = _66188 ^ _66199;
  wire _66201 = uncoded_block[1362] ^ uncoded_block[1387];
  wire _66202 = uncoded_block[1398] ^ uncoded_block[1436];
  wire _66203 = _66201 ^ _66202;
  wire _66204 = _60900 ^ _34623;
  wire _66205 = _66203 ^ _66204;
  wire _66206 = _50331 ^ _14492;
  wire _66207 = _58311 ^ _10176;
  wire _66208 = _66206 ^ _66207;
  wire _66209 = _66205 ^ _66208;
  wire _66210 = uncoded_block[1607] ^ uncoded_block[1617];
  wire _66211 = uncoded_block[1640] ^ uncoded_block[1666];
  wire _66212 = _66210 ^ _66211;
  wire _66213 = uncoded_block[1667] ^ uncoded_block[1693];
  wire _66214 = uncoded_block[1698] ^ uncoded_block[1710];
  wire _66215 = _66213 ^ _66214;
  wire _66216 = _66212 ^ _66215;
  wire _66217 = _66216 ^ uncoded_block[1718];
  wire _66218 = _66209 ^ _66217;
  wire _66219 = _66200 ^ _66218;
  wire _66220 = _66176 ^ _66219;
  wire _66221 = uncoded_block[14] ^ uncoded_block[47];
  wire _66222 = _66221 ^ _7374;
  wire _66223 = uncoded_block[116] ^ uncoded_block[149];
  wire _66224 = uncoded_block[174] ^ uncoded_block[212];
  wire _66225 = _66223 ^ _66224;
  wire _66226 = _66222 ^ _66225;
  wire _66227 = uncoded_block[248] ^ uncoded_block[292];
  wire _66228 = uncoded_block[319] ^ uncoded_block[345];
  wire _66229 = _66227 ^ _66228;
  wire _66230 = uncoded_block[362] ^ uncoded_block[392];
  wire _66231 = uncoded_block[440] ^ uncoded_block[488];
  wire _66232 = _66230 ^ _66231;
  wire _66233 = _66229 ^ _66232;
  wire _66234 = _66226 ^ _66233;
  wire _66235 = uncoded_block[503] ^ uncoded_block[522];
  wire _66236 = uncoded_block[537] ^ uncoded_block[575];
  wire _66237 = _66235 ^ _66236;
  wire _66238 = uncoded_block[613] ^ uncoded_block[627];
  wire _66239 = uncoded_block[635] ^ uncoded_block[689];
  wire _66240 = _66238 ^ _66239;
  wire _66241 = _66237 ^ _66240;
  wire _66242 = uncoded_block[702] ^ uncoded_block[731];
  wire _66243 = uncoded_block[767] ^ uncoded_block[779];
  wire _66244 = _66242 ^ _66243;
  wire _66245 = uncoded_block[871] ^ uncoded_block[912];
  wire _66246 = _26160 ^ _66245;
  wire _66247 = _66244 ^ _66246;
  wire _66248 = _66241 ^ _66247;
  wire _66249 = _66234 ^ _66248;
  wire _66250 = uncoded_block[980] ^ uncoded_block[1039];
  wire _66251 = _64965 ^ _66250;
  wire _66252 = uncoded_block[1046] ^ uncoded_block[1067];
  wire _66253 = uncoded_block[1068] ^ uncoded_block[1152];
  wire _66254 = _66252 ^ _66253;
  wire _66255 = _66251 ^ _66254;
  wire _66256 = uncoded_block[1159] ^ uncoded_block[1168];
  wire _66257 = uncoded_block[1183] ^ uncoded_block[1239];
  wire _66258 = _66256 ^ _66257;
  wire _66259 = uncoded_block[1245] ^ uncoded_block[1298];
  wire _66260 = uncoded_block[1311] ^ uncoded_block[1350];
  wire _66261 = _66259 ^ _66260;
  wire _66262 = _66258 ^ _66261;
  wire _66263 = _66255 ^ _66262;
  wire _66264 = uncoded_block[1402] ^ uncoded_block[1414];
  wire _66265 = uncoded_block[1438] ^ uncoded_block[1480];
  wire _66266 = _66264 ^ _66265;
  wire _66267 = uncoded_block[1500] ^ uncoded_block[1519];
  wire _66268 = uncoded_block[1534] ^ uncoded_block[1559];
  wire _66269 = _66267 ^ _66268;
  wire _66270 = _66266 ^ _66269;
  wire _66271 = uncoded_block[1599] ^ uncoded_block[1625];
  wire _66272 = uncoded_block[1633] ^ uncoded_block[1698];
  wire _66273 = _66271 ^ _66272;
  wire _66274 = _66273 ^ uncoded_block[1700];
  wire _66275 = _66270 ^ _66274;
  wire _66276 = _66263 ^ _66275;
  wire _66277 = _66249 ^ _66276;
  wire _66278 = uncoded_block[80] ^ uncoded_block[90];
  wire _66279 = uncoded_block[113] ^ uncoded_block[121];
  wire _66280 = _66278 ^ _66279;
  wire _66281 = uncoded_block[240] ^ uncoded_block[279];
  wire _66282 = _64644 ^ _66281;
  wire _66283 = _66280 ^ _66282;
  wire _66284 = uncoded_block[283] ^ uncoded_block[326];
  wire _66285 = _66284 ^ _31863;
  wire _66286 = _64660 ^ _58440;
  wire _66287 = _66285 ^ _66286;
  wire _66288 = _66283 ^ _66287;
  wire _66289 = uncoded_block[510] ^ uncoded_block[550];
  wire _66290 = uncoded_block[567] ^ uncoded_block[606];
  wire _66291 = _66289 ^ _66290;
  wire _66292 = uncoded_block[685] ^ uncoded_block[714];
  wire _66293 = _6968 ^ _66292;
  wire _66294 = _66291 ^ _66293;
  wire _66295 = uncoded_block[743] ^ uncoded_block[767];
  wire _66296 = uncoded_block[778] ^ uncoded_block[814];
  wire _66297 = _66295 ^ _66296;
  wire _66298 = uncoded_block[897] ^ uncoded_block[912];
  wire _66299 = _64702 ^ _66298;
  wire _66300 = _66297 ^ _66299;
  wire _66301 = _66294 ^ _66300;
  wire _66302 = _66288 ^ _66301;
  wire _66303 = uncoded_block[1007] ^ uncoded_block[1035];
  wire _66304 = _57704 ^ _66303;
  wire _66305 = uncoded_block[1060] ^ uncoded_block[1094];
  wire _66306 = uncoded_block[1114] ^ uncoded_block[1127];
  wire _66307 = _66305 ^ _66306;
  wire _66308 = _66304 ^ _66307;
  wire _66309 = uncoded_block[1181] ^ uncoded_block[1211];
  wire _66310 = uncoded_block[1255] ^ uncoded_block[1263];
  wire _66311 = _66309 ^ _66310;
  wire _66312 = uncoded_block[1296] ^ uncoded_block[1327];
  wire _66313 = uncoded_block[1342] ^ uncoded_block[1378];
  wire _66314 = _66312 ^ _66313;
  wire _66315 = _66311 ^ _66314;
  wire _66316 = _66308 ^ _66315;
  wire _66317 = uncoded_block[1399] ^ uncoded_block[1541];
  wire _66318 = _66317 ^ _57775;
  wire _66319 = uncoded_block[1599] ^ uncoded_block[1629];
  wire _66320 = _64760 ^ _66319;
  wire _66321 = _66318 ^ _66320;
  wire _66322 = uncoded_block[1635] ^ uncoded_block[1672];
  wire _66323 = uncoded_block[1681] ^ uncoded_block[1719];
  wire _66324 = _66322 ^ _66323;
  wire _66325 = _66324 ^ uncoded_block[1722];
  wire _66326 = _66321 ^ _66325;
  wire _66327 = _66316 ^ _66326;
  wire _66328 = _66302 ^ _66327;
  wire _66329 = uncoded_block[41] ^ uncoded_block[57];
  wire _66330 = _874 ^ _66329;
  wire _66331 = _62460 ^ _61576;
  wire _66332 = _66330 ^ _66331;
  wire _66333 = uncoded_block[143] ^ uncoded_block[174];
  wire _66334 = _59257 ^ _66333;
  wire _66335 = uncoded_block[218] ^ uncoded_block[238];
  wire _66336 = _8018 ^ _66335;
  wire _66337 = _66334 ^ _66336;
  wire _66338 = _66332 ^ _66337;
  wire _66339 = uncoded_block[239] ^ uncoded_block[270];
  wire _66340 = uncoded_block[272] ^ uncoded_block[286];
  wire _66341 = _66339 ^ _66340;
  wire _66342 = uncoded_block[307] ^ uncoded_block[325];
  wire _66343 = _66342 ^ _2587;
  wire _66344 = _66341 ^ _66343;
  wire _66345 = uncoded_block[373] ^ uncoded_block[408];
  wire _66346 = _61604 ^ _66345;
  wire _66347 = _24711 ^ _4882;
  wire _66348 = _66346 ^ _66347;
  wire _66349 = _66344 ^ _66348;
  wire _66350 = _66338 ^ _66349;
  wire _66351 = uncoded_block[453] ^ uncoded_block[473];
  wire _66352 = _66351 ^ _65494;
  wire _66353 = uncoded_block[514] ^ uncoded_block[549];
  wire _66354 = uncoded_block[550] ^ uncoded_block[578];
  wire _66355 = _66353 ^ _66354;
  wire _66356 = _66352 ^ _66355;
  wire _66357 = uncoded_block[588] ^ uncoded_block[605];
  wire _66358 = _66357 ^ _61635;
  wire _66359 = uncoded_block[635] ^ uncoded_block[649];
  wire _66360 = _66359 ^ _63070;
  wire _66361 = _66358 ^ _66360;
  wire _66362 = _66356 ^ _66361;
  wire _66363 = uncoded_block[684] ^ uncoded_block[699];
  wire _66364 = _66363 ^ _66028;
  wire _66365 = uncoded_block[766] ^ uncoded_block[805];
  wire _66366 = _13761 ^ _66365;
  wire _66367 = _66364 ^ _66366;
  wire _66368 = _11029 ^ _6402;
  wire _66369 = _26164 ^ _61482;
  wire _66370 = _66368 ^ _66369;
  wire _66371 = _66367 ^ _66370;
  wire _66372 = _66362 ^ _66371;
  wire _66373 = _66350 ^ _66372;
  wire _66374 = uncoded_block[906] ^ uncoded_block[912];
  wire _66375 = uncoded_block[938] ^ uncoded_block[960];
  wire _66376 = _66374 ^ _66375;
  wire _66377 = uncoded_block[997] ^ uncoded_block[1034];
  wire _66378 = _8282 ^ _66377;
  wire _66379 = _66376 ^ _66378;
  wire _66380 = uncoded_block[1041] ^ uncoded_block[1053];
  wire _66381 = uncoded_block[1058] ^ uncoded_block[1086];
  wire _66382 = _66380 ^ _66381;
  wire _66383 = _537 ^ _59567;
  wire _66384 = _66382 ^ _66383;
  wire _66385 = _66379 ^ _66384;
  wire _66386 = uncoded_block[1143] ^ uncoded_block[1179];
  wire _66387 = _558 ^ _66386;
  wire _66388 = uncoded_block[1180] ^ uncoded_block[1188];
  wire _66389 = uncoded_block[1207] ^ uncoded_block[1255];
  wire _66390 = _66388 ^ _66389;
  wire _66391 = _66387 ^ _66390;
  wire _66392 = uncoded_block[1272] ^ uncoded_block[1286];
  wire _66393 = _61711 ^ _66392;
  wire _66394 = uncoded_block[1293] ^ uncoded_block[1322];
  wire _66395 = uncoded_block[1326] ^ uncoded_block[1351];
  wire _66396 = _66394 ^ _66395;
  wire _66397 = _66393 ^ _66396;
  wire _66398 = _66391 ^ _66397;
  wire _66399 = _66385 ^ _66398;
  wire _66400 = _2283 ^ _61726;
  wire _66401 = uncoded_block[1400] ^ uncoded_block[1421];
  wire _66402 = uncoded_block[1451] ^ uncoded_block[1459];
  wire _66403 = _66401 ^ _66402;
  wire _66404 = _66400 ^ _66403;
  wire _66405 = uncoded_block[1470] ^ uncoded_block[1475];
  wire _66406 = _25416 ^ _66405;
  wire _66407 = uncoded_block[1547] ^ uncoded_block[1558];
  wire _66408 = uncoded_block[1563] ^ uncoded_block[1589];
  wire _66409 = _66407 ^ _66408;
  wire _66410 = _66406 ^ _66409;
  wire _66411 = _66404 ^ _66410;
  wire _66412 = uncoded_block[1609] ^ uncoded_block[1621];
  wire _66413 = uncoded_block[1653] ^ uncoded_block[1666];
  wire _66414 = _66412 ^ _66413;
  wire _66415 = _41009 ^ uncoded_block[1721];
  wire _66416 = _66414 ^ _66415;
  wire _66417 = _66411 ^ _66416;
  wire _66418 = _66399 ^ _66417;
  wire _66419 = _66373 ^ _66418;
  wire _66420 = uncoded_block[23] ^ uncoded_block[62];
  wire _66421 = uncoded_block[101] ^ uncoded_block[142];
  wire _66422 = _66420 ^ _66421;
  wire _66423 = uncoded_block[159] ^ uncoded_block[193];
  wire _66424 = uncoded_block[215] ^ uncoded_block[240];
  wire _66425 = _66423 ^ _66424;
  wire _66426 = _66422 ^ _66425;
  wire _66427 = uncoded_block[289] ^ uncoded_block[322];
  wire _66428 = uncoded_block[348] ^ uncoded_block[375];
  wire _66429 = _66427 ^ _66428;
  wire _66430 = uncoded_block[409] ^ uncoded_block[429];
  wire _66431 = _66430 ^ _62020;
  wire _66432 = _66429 ^ _66431;
  wire _66433 = _66426 ^ _66432;
  wire _66434 = uncoded_block[564] ^ uncoded_block[610];
  wire _66435 = _62021 ^ _66434;
  wire _66436 = uncoded_block[626] ^ uncoded_block[643];
  wire _66437 = uncoded_block[716] ^ uncoded_block[721];
  wire _66438 = _66436 ^ _66437;
  wire _66439 = _66435 ^ _66438;
  wire _66440 = uncoded_block[765] ^ uncoded_block[784];
  wire _66441 = _1987 ^ _66440;
  wire _66442 = uncoded_block[817] ^ uncoded_block[884];
  wire _66443 = _66442 ^ _7066;
  wire _66444 = _66441 ^ _66443;
  wire _66445 = _66439 ^ _66444;
  wire _66446 = _66433 ^ _66445;
  wire _66447 = uncoded_block[957] ^ uncoded_block[981];
  wire _66448 = uncoded_block[1015] ^ uncoded_block[1028];
  wire _66449 = _66447 ^ _66448;
  wire _66450 = uncoded_block[1068] ^ uncoded_block[1081];
  wire _66451 = uncoded_block[1121] ^ uncoded_block[1135];
  wire _66452 = _66450 ^ _66451;
  wire _66453 = _66449 ^ _66452;
  wire _66454 = uncoded_block[1221] ^ uncoded_block[1247];
  wire _66455 = _2200 ^ _66454;
  wire _66456 = uncoded_block[1267] ^ uncoded_block[1294];
  wire _66457 = uncoded_block[1296] ^ uncoded_block[1334];
  wire _66458 = _66456 ^ _66457;
  wire _66459 = _66455 ^ _66458;
  wire _66460 = _66453 ^ _66459;
  wire _66461 = uncoded_block[1346] ^ uncoded_block[1366];
  wire _66462 = uncoded_block[1409] ^ uncoded_block[1476];
  wire _66463 = _66461 ^ _66462;
  wire _66464 = uncoded_block[1477] ^ uncoded_block[1501];
  wire _66465 = uncoded_block[1551] ^ uncoded_block[1570];
  wire _66466 = _66464 ^ _66465;
  wire _66467 = _66463 ^ _66466;
  wire _66468 = uncoded_block[1611] ^ uncoded_block[1644];
  wire _66469 = uncoded_block[1665] ^ uncoded_block[1687];
  wire _66470 = _66468 ^ _66469;
  wire _66471 = _66470 ^ uncoded_block[1722];
  wire _66472 = _66467 ^ _66471;
  wire _66473 = _66460 ^ _66472;
  wire _66474 = _66446 ^ _66473;
  wire _66475 = uncoded_block[1] ^ uncoded_block[52];
  wire _66476 = uncoded_block[57] ^ uncoded_block[109];
  wire _66477 = _66475 ^ _66476;
  wire _66478 = uncoded_block[117] ^ uncoded_block[168];
  wire _66479 = uncoded_block[173] ^ uncoded_block[194];
  wire _66480 = _66478 ^ _66479;
  wire _66481 = _66477 ^ _66480;
  wire _66482 = uncoded_block[247] ^ uncoded_block[277];
  wire _66483 = uncoded_block[306] ^ uncoded_block[327];
  wire _66484 = _66482 ^ _66483;
  wire _66485 = uncoded_block[349] ^ uncoded_block[373];
  wire _66486 = uncoded_block[403] ^ uncoded_block[424];
  wire _66487 = _66485 ^ _66486;
  wire _66488 = _66484 ^ _66487;
  wire _66489 = _66481 ^ _66488;
  wire _66490 = uncoded_block[453] ^ uncoded_block[494];
  wire _66491 = uncoded_block[531] ^ uncoded_block[548];
  wire _66492 = _66490 ^ _66491;
  wire _66493 = _57661 ^ _3505;
  wire _66494 = _66492 ^ _66493;
  wire _66495 = uncoded_block[677] ^ uncoded_block[697];
  wire _66496 = uncoded_block[771] ^ uncoded_block[825];
  wire _66497 = _66495 ^ _66496;
  wire _66498 = uncoded_block[828] ^ uncoded_block[839];
  wire _66499 = uncoded_block[858] ^ uncoded_block[928];
  wire _66500 = _66498 ^ _66499;
  wire _66501 = _66497 ^ _66500;
  wire _66502 = _66494 ^ _66501;
  wire _66503 = _66489 ^ _66502;
  wire _66504 = uncoded_block[940] ^ uncoded_block[955];
  wire _66505 = uncoded_block[980] ^ uncoded_block[1014];
  wire _66506 = _66504 ^ _66505;
  wire _66507 = uncoded_block[1054] ^ uncoded_block[1091];
  wire _66508 = uncoded_block[1120] ^ uncoded_block[1133];
  wire _66509 = _66507 ^ _66508;
  wire _66510 = _66506 ^ _66509;
  wire _66511 = uncoded_block[1183] ^ uncoded_block[1210];
  wire _66512 = uncoded_block[1221] ^ uncoded_block[1240];
  wire _66513 = _66511 ^ _66512;
  wire _66514 = uncoded_block[1271] ^ uncoded_block[1292];
  wire _66515 = uncoded_block[1323] ^ uncoded_block[1333];
  wire _66516 = _66514 ^ _66515;
  wire _66517 = _66513 ^ _66516;
  wire _66518 = _66510 ^ _66517;
  wire _66519 = uncoded_block[1343] ^ uncoded_block[1372];
  wire _66520 = uncoded_block[1414] ^ uncoded_block[1430];
  wire _66521 = _66519 ^ _66520;
  wire _66522 = uncoded_block[1447] ^ uncoded_block[1483];
  wire _66523 = uncoded_block[1499] ^ uncoded_block[1506];
  wire _66524 = _66522 ^ _66523;
  wire _66525 = _66521 ^ _66524;
  wire _66526 = uncoded_block[1587] ^ uncoded_block[1618];
  wire _66527 = uncoded_block[1646] ^ uncoded_block[1699];
  wire _66528 = _66526 ^ _66527;
  wire _66529 = _66528 ^ uncoded_block[1706];
  wire _66530 = _66525 ^ _66529;
  wire _66531 = _66518 ^ _66530;
  wire _66532 = _66503 ^ _66531;
  wire _66533 = uncoded_block[3] ^ uncoded_block[37];
  wire _66534 = _66533 ^ _65059;
  wire _66535 = uncoded_block[181] ^ uncoded_block[207];
  wire _66536 = _10828 ^ _66535;
  wire _66537 = _66534 ^ _66536;
  wire _66538 = uncoded_block[247] ^ uncoded_block[262];
  wire _66539 = uncoded_block[313] ^ uncoded_block[331];
  wire _66540 = _66538 ^ _66539;
  wire _66541 = uncoded_block[336] ^ uncoded_block[370];
  wire _66542 = uncoded_block[396] ^ uncoded_block[431];
  wire _66543 = _66541 ^ _66542;
  wire _66544 = _66540 ^ _66543;
  wire _66545 = _66537 ^ _66544;
  wire _66546 = uncoded_block[463] ^ uncoded_block[471];
  wire _66547 = uncoded_block[535] ^ uncoded_block[548];
  wire _66548 = _66546 ^ _66547;
  wire _66549 = uncoded_block[562] ^ uncoded_block[599];
  wire _66550 = uncoded_block[631] ^ uncoded_block[672];
  wire _66551 = _66549 ^ _66550;
  wire _66552 = _66548 ^ _66551;
  wire _66553 = uncoded_block[686] ^ uncoded_block[732];
  wire _66554 = uncoded_block[769] ^ uncoded_block[787];
  wire _66555 = _66553 ^ _66554;
  wire _66556 = uncoded_block[819] ^ uncoded_block[862];
  wire _66557 = uncoded_block[868] ^ uncoded_block[918];
  wire _66558 = _66556 ^ _66557;
  wire _66559 = _66555 ^ _66558;
  wire _66560 = _66552 ^ _66559;
  wire _66561 = _66545 ^ _66560;
  wire _66562 = uncoded_block[925] ^ uncoded_block[960];
  wire _66563 = uncoded_block[991] ^ uncoded_block[1024];
  wire _66564 = _66562 ^ _66563;
  wire _66565 = uncoded_block[1037] ^ uncoded_block[1071];
  wire _66566 = _66565 ^ _51674;
  wire _66567 = _66564 ^ _66566;
  wire _66568 = uncoded_block[1117] ^ uncoded_block[1165];
  wire _66569 = _66568 ^ _63116;
  wire _66570 = uncoded_block[1220] ^ uncoded_block[1227];
  wire _66571 = uncoded_block[1254] ^ uncoded_block[1288];
  wire _66572 = _66570 ^ _66571;
  wire _66573 = _66569 ^ _66572;
  wire _66574 = _66567 ^ _66573;
  wire _66575 = uncoded_block[1409] ^ uncoded_block[1418];
  wire _66576 = _66313 ^ _66575;
  wire _66577 = uncoded_block[1467] ^ uncoded_block[1492];
  wire _66578 = _65015 ^ _66577;
  wire _66579 = _66576 ^ _66578;
  wire _66580 = uncoded_block[1528] ^ uncoded_block[1603];
  wire _66581 = uncoded_block[1637] ^ uncoded_block[1653];
  wire _66582 = _66580 ^ _66581;
  wire _66583 = _66582 ^ uncoded_block[1669];
  wire _66584 = _66579 ^ _66583;
  wire _66585 = _66574 ^ _66584;
  wire _66586 = _66561 ^ _66585;
  wire _66587 = uncoded_block[5] ^ uncoded_block[51];
  wire _66588 = uncoded_block[85] ^ uncoded_block[108];
  wire _66589 = _66587 ^ _66588;
  wire _66590 = uncoded_block[146] ^ uncoded_block[166];
  wire _66591 = uncoded_block[194] ^ uncoded_block[203];
  wire _66592 = _66590 ^ _66591;
  wire _66593 = _66589 ^ _66592;
  wire _66594 = uncoded_block[303] ^ uncoded_block[317];
  wire _66595 = _1775 ^ _66594;
  wire _66596 = uncoded_block[396] ^ uncoded_block[428];
  wire _66597 = _40360 ^ _66596;
  wire _66598 = _66595 ^ _66597;
  wire _66599 = _66593 ^ _66598;
  wire _66600 = uncoded_block[463] ^ uncoded_block[495];
  wire _66601 = uncoded_block[511] ^ uncoded_block[536];
  wire _66602 = _66600 ^ _66601;
  wire _66603 = uncoded_block[575] ^ uncoded_block[593];
  wire _66604 = uncoded_block[624] ^ uncoded_block[650];
  wire _66605 = _66603 ^ _66604;
  wire _66606 = _66602 ^ _66605;
  wire _66607 = uncoded_block[671] ^ uncoded_block[720];
  wire _66608 = _66607 ^ _40817;
  wire _66609 = uncoded_block[786] ^ uncoded_block[798];
  wire _66610 = uncoded_block[835] ^ uncoded_block[880];
  wire _66611 = _66609 ^ _66610;
  wire _66612 = _66608 ^ _66611;
  wire _66613 = _66606 ^ _66612;
  wire _66614 = _66599 ^ _66613;
  wire _66615 = uncoded_block[894] ^ uncoded_block[933];
  wire _66616 = _66615 ^ _6457;
  wire _66617 = uncoded_block[1026] ^ uncoded_block[1076];
  wire _66618 = _61887 ^ _66617;
  wire _66619 = _66616 ^ _66618;
  wire _66620 = uncoded_block[1092] ^ uncoded_block[1108];
  wire _66621 = uncoded_block[1155] ^ uncoded_block[1162];
  wire _66622 = _66620 ^ _66621;
  wire _66623 = uncoded_block[1213] ^ uncoded_block[1240];
  wire _66624 = uncoded_block[1303] ^ uncoded_block[1319];
  wire _66625 = _66623 ^ _66624;
  wire _66626 = _66622 ^ _66625;
  wire _66627 = _66619 ^ _66626;
  wire _66628 = uncoded_block[1338] ^ uncoded_block[1354];
  wire _66629 = uncoded_block[1431] ^ uncoded_block[1464];
  wire _66630 = _66628 ^ _66629;
  wire _66631 = uncoded_block[1471] ^ uncoded_block[1484];
  wire _66632 = uncoded_block[1522] ^ uncoded_block[1596];
  wire _66633 = _66631 ^ _66632;
  wire _66634 = _66630 ^ _66633;
  wire _66635 = uncoded_block[1638] ^ uncoded_block[1652];
  wire _66636 = uncoded_block[1666] ^ uncoded_block[1690];
  wire _66637 = _66635 ^ _66636;
  wire _66638 = _66637 ^ uncoded_block[1696];
  wire _66639 = _66634 ^ _66638;
  wire _66640 = _66627 ^ _66639;
  wire _66641 = _66614 ^ _66640;
  wire _66642 = uncoded_block[73] ^ uncoded_block[81];
  wire _66643 = _66129 ^ _66642;
  wire _66644 = uncoded_block[199] ^ uncoded_block[210];
  wire _66645 = _59257 ^ _66644;
  wire _66646 = _66643 ^ _66645;
  wire _66647 = uncoded_block[225] ^ uncoded_block[277];
  wire _66648 = _66647 ^ _32682;
  wire _66649 = uncoded_block[337] ^ uncoded_block[343];
  wire _66650 = uncoded_block[412] ^ uncoded_block[444];
  wire _66651 = _66649 ^ _66650;
  wire _66652 = _66648 ^ _66651;
  wire _66653 = _66646 ^ _66652;
  wire _66654 = uncoded_block[523] ^ uncoded_block[534];
  wire _66655 = _20592 ^ _66654;
  wire _66656 = uncoded_block[572] ^ uncoded_block[589];
  wire _66657 = uncoded_block[625] ^ uncoded_block[637];
  wire _66658 = _66656 ^ _66657;
  wire _66659 = _66655 ^ _66658;
  wire _66660 = uncoded_block[680] ^ uncoded_block[708];
  wire _66661 = uncoded_block[734] ^ uncoded_block[745];
  wire _66662 = _66660 ^ _66661;
  wire _66663 = uncoded_block[845] ^ uncoded_block[858];
  wire _66664 = _64385 ^ _66663;
  wire _66665 = _66662 ^ _66664;
  wire _66666 = _66659 ^ _66665;
  wire _66667 = _66653 ^ _66666;
  wire _66668 = uncoded_block[907] ^ uncoded_block[939];
  wire _66669 = uncoded_block[959] ^ uncoded_block[975];
  wire _66670 = _66668 ^ _66669;
  wire _66671 = uncoded_block[1042] ^ uncoded_block[1077];
  wire _66672 = uncoded_block[1105] ^ uncoded_block[1113];
  wire _66673 = _66671 ^ _66672;
  wire _66674 = _66670 ^ _66673;
  wire _66675 = uncoded_block[1121] ^ uncoded_block[1134];
  wire _66676 = uncoded_block[1171] ^ uncoded_block[1202];
  wire _66677 = _66675 ^ _66676;
  wire _66678 = uncoded_block[1259] ^ uncoded_block[1264];
  wire _66679 = uncoded_block[1297] ^ uncoded_block[1330];
  wire _66680 = _66678 ^ _66679;
  wire _66681 = _66677 ^ _66680;
  wire _66682 = _66674 ^ _66681;
  wire _66683 = uncoded_block[1339] ^ uncoded_block[1360];
  wire _66684 = _66683 ^ _60085;
  wire _66685 = uncoded_block[1437] ^ uncoded_block[1505];
  wire _66686 = uncoded_block[1540] ^ uncoded_block[1604];
  wire _66687 = _66685 ^ _66686;
  wire _66688 = _66684 ^ _66687;
  wire _66689 = uncoded_block[1605] ^ uncoded_block[1666];
  wire _66690 = uncoded_block[1686] ^ uncoded_block[1703];
  wire _66691 = _66689 ^ _66690;
  wire _66692 = _66691 ^ uncoded_block[1710];
  wire _66693 = _66688 ^ _66692;
  wire _66694 = _66682 ^ _66693;
  wire _66695 = _66667 ^ _66694;
  wire _66696 = uncoded_block[10] ^ uncoded_block[38];
  wire _66697 = uncoded_block[94] ^ uncoded_block[110];
  wire _66698 = _66696 ^ _66697;
  wire _66699 = uncoded_block[184] ^ uncoded_block[228];
  wire _66700 = _60486 ^ _66699;
  wire _66701 = _66698 ^ _66700;
  wire _66702 = uncoded_block[322] ^ uncoded_block[334];
  wire _66703 = _65353 ^ _66702;
  wire _66704 = uncoded_block[380] ^ uncoded_block[399];
  wire _66705 = uncoded_block[420] ^ uncoded_block[467];
  wire _66706 = _66704 ^ _66705;
  wire _66707 = _66703 ^ _66706;
  wire _66708 = _66701 ^ _66707;
  wire _66709 = uncoded_block[522] ^ uncoded_block[565];
  wire _66710 = _65363 ^ _66709;
  wire _66711 = uncoded_block[584] ^ uncoded_block[621];
  wire _66712 = uncoded_block[654] ^ uncoded_block[680];
  wire _66713 = _66711 ^ _66712;
  wire _66714 = _66710 ^ _66713;
  wire _66715 = uncoded_block[715] ^ uncoded_block[726];
  wire _66716 = uncoded_block[729] ^ uncoded_block[795];
  wire _66717 = _66715 ^ _66716;
  wire _66718 = uncoded_block[800] ^ uncoded_block[863];
  wire _66719 = _66718 ^ _60543;
  wire _66720 = _66717 ^ _66719;
  wire _66721 = _66714 ^ _66720;
  wire _66722 = _66708 ^ _66721;
  wire _66723 = uncoded_block[905] ^ uncoded_block[947];
  wire _66724 = uncoded_block[984] ^ uncoded_block[1012];
  wire _66725 = _66723 ^ _66724;
  wire _66726 = uncoded_block[1052] ^ uncoded_block[1086];
  wire _66727 = uncoded_block[1088] ^ uncoded_block[1127];
  wire _66728 = _66726 ^ _66727;
  wire _66729 = _66725 ^ _66728;
  wire _66730 = uncoded_block[1151] ^ uncoded_block[1175];
  wire _66731 = uncoded_block[1200] ^ uncoded_block[1242];
  wire _66732 = _66730 ^ _66731;
  wire _66733 = uncoded_block[1260] ^ uncoded_block[1301];
  wire _66734 = uncoded_block[1313] ^ uncoded_block[1346];
  wire _66735 = _66733 ^ _66734;
  wire _66736 = _66732 ^ _66735;
  wire _66737 = _66729 ^ _66736;
  wire _66738 = uncoded_block[1382] ^ uncoded_block[1406];
  wire _66739 = uncoded_block[1413] ^ uncoded_block[1433];
  wire _66740 = _66738 ^ _66739;
  wire _66741 = uncoded_block[1574] ^ uncoded_block[1612];
  wire _66742 = _65403 ^ _66741;
  wire _66743 = _66740 ^ _66742;
  wire _66744 = uncoded_block[1621] ^ uncoded_block[1650];
  wire _66745 = _66744 ^ _60610;
  wire _66746 = _66745 ^ uncoded_block[1706];
  wire _66747 = _66743 ^ _66746;
  wire _66748 = _66737 ^ _66747;
  wire _66749 = _66722 ^ _66748;
  wire _66750 = uncoded_block[29] ^ uncoded_block[54];
  wire _66751 = _32609 ^ _66750;
  wire _66752 = uncoded_block[77] ^ uncoded_block[84];
  wire _66753 = uncoded_block[90] ^ uncoded_block[118];
  wire _66754 = _66752 ^ _66753;
  wire _66755 = _66751 ^ _66754;
  wire _66756 = uncoded_block[131] ^ uncoded_block[148];
  wire _66757 = uncoded_block[163] ^ uncoded_block[177];
  wire _66758 = _66756 ^ _66757;
  wire _66759 = uncoded_block[205] ^ uncoded_block[233];
  wire _66760 = uncoded_block[236] ^ uncoded_block[265];
  wire _66761 = _66759 ^ _66760;
  wire _66762 = _66758 ^ _66761;
  wire _66763 = _66755 ^ _66762;
  wire _66764 = uncoded_block[270] ^ uncoded_block[298];
  wire _66765 = _66764 ^ _59030;
  wire _66766 = uncoded_block[317] ^ uncoded_block[340];
  wire _66767 = uncoded_block[356] ^ uncoded_block[369];
  wire _66768 = _66766 ^ _66767;
  wire _66769 = _66765 ^ _66768;
  wire _66770 = uncoded_block[386] ^ uncoded_block[394];
  wire _66771 = uncoded_block[422] ^ uncoded_block[449];
  wire _66772 = _66770 ^ _66771;
  wire _66773 = uncoded_block[463] ^ uncoded_block[497];
  wire _66774 = uncoded_block[498] ^ uncoded_block[512];
  wire _66775 = _66773 ^ _66774;
  wire _66776 = _66772 ^ _66775;
  wire _66777 = _66769 ^ _66776;
  wire _66778 = _66763 ^ _66777;
  wire _66779 = uncoded_block[513] ^ uncoded_block[528];
  wire _66780 = uncoded_block[557] ^ uncoded_block[569];
  wire _66781 = _66779 ^ _66780;
  wire _66782 = uncoded_block[603] ^ uncoded_block[638];
  wire _66783 = _12057 ^ _66782;
  wire _66784 = _66781 ^ _66783;
  wire _66785 = uncoded_block[652] ^ uncoded_block[669];
  wire _66786 = _19177 ^ _66785;
  wire _66787 = uncoded_block[677] ^ uncoded_block[700];
  wire _66788 = uncoded_block[742] ^ uncoded_block[755];
  wire _66789 = _66787 ^ _66788;
  wire _66790 = _66786 ^ _66789;
  wire _66791 = _66784 ^ _66790;
  wire _66792 = uncoded_block[788] ^ uncoded_block[799];
  wire _66793 = _9917 ^ _66792;
  wire _66794 = uncoded_block[852] ^ uncoded_block[875];
  wire _66795 = _59316 ^ _66794;
  wire _66796 = _66793 ^ _66795;
  wire _66797 = uncoded_block[896] ^ uncoded_block[923];
  wire _66798 = _55042 ^ _66797;
  wire _66799 = uncoded_block[950] ^ uncoded_block[968];
  wire _66800 = _13809 ^ _66799;
  wire _66801 = _66798 ^ _66800;
  wire _66802 = _66796 ^ _66801;
  wire _66803 = _66791 ^ _66802;
  wire _66804 = _66778 ^ _66803;
  wire _66805 = uncoded_block[976] ^ uncoded_block[999];
  wire _66806 = _66805 ^ _48255;
  wire _66807 = _62068 ^ _14366;
  wire _66808 = _66806 ^ _66807;
  wire _66809 = uncoded_block[1120] ^ uncoded_block[1147];
  wire _66810 = uncoded_block[1157] ^ uncoded_block[1171];
  wire _66811 = _66809 ^ _66810;
  wire _66812 = uncoded_block[1190] ^ uncoded_block[1202];
  wire _66813 = uncoded_block[1237] ^ uncoded_block[1248];
  wire _66814 = _66812 ^ _66813;
  wire _66815 = _66811 ^ _66814;
  wire _66816 = _66808 ^ _66815;
  wire _66817 = uncoded_block[1272] ^ uncoded_block[1308];
  wire _66818 = _66817 ^ _653;
  wire _66819 = uncoded_block[1321] ^ uncoded_block[1340];
  wire _66820 = _66819 ^ _673;
  wire _66821 = _66818 ^ _66820;
  wire _66822 = uncoded_block[1383] ^ uncoded_block[1403];
  wire _66823 = _66822 ^ _58003;
  wire _66824 = uncoded_block[1478] ^ uncoded_block[1498];
  wire _66825 = _35423 ^ _66824;
  wire _66826 = _66823 ^ _66825;
  wire _66827 = _66821 ^ _66826;
  wire _66828 = _66816 ^ _66827;
  wire _66829 = _23624 ^ _50331;
  wire _66830 = uncoded_block[1545] ^ uncoded_block[1559];
  wire _66831 = uncoded_block[1560] ^ uncoded_block[1587];
  wire _66832 = _66830 ^ _66831;
  wire _66833 = _66829 ^ _66832;
  wire _66834 = uncoded_block[1591] ^ uncoded_block[1598];
  wire _66835 = uncoded_block[1617] ^ uncoded_block[1640];
  wire _66836 = _66834 ^ _66835;
  wire _66837 = uncoded_block[1667] ^ uncoded_block[1674];
  wire _66838 = _48771 ^ _66837;
  wire _66839 = _66836 ^ _66838;
  wire _66840 = _66833 ^ _66839;
  wire _66841 = uncoded_block[1698] ^ uncoded_block[1713];
  wire _66842 = _66841 ^ uncoded_block[1721];
  wire _66843 = _66840 ^ _66842;
  wire _66844 = _66828 ^ _66843;
  wire _66845 = _66804 ^ _66844;
  wire _66846 = uncoded_block[15] ^ uncoded_block[35];
  wire _66847 = uncoded_block[56] ^ uncoded_block[96];
  wire _66848 = _66846 ^ _66847;
  wire _66849 = uncoded_block[163] ^ uncoded_block[209];
  wire _66850 = uncoded_block[216] ^ uncoded_block[247];
  wire _66851 = _66849 ^ _66850;
  wire _66852 = _66848 ^ _66851;
  wire _66853 = uncoded_block[272] ^ uncoded_block[287];
  wire _66854 = uncoded_block[322] ^ uncoded_block[344];
  wire _66855 = _66853 ^ _66854;
  wire _66856 = uncoded_block[389] ^ uncoded_block[418];
  wire _66857 = uncoded_block[426] ^ uncoded_block[459];
  wire _66858 = _66856 ^ _66857;
  wire _66859 = _66855 ^ _66858;
  wire _66860 = _66852 ^ _66859;
  wire _66861 = uncoded_block[482] ^ uncoded_block[516];
  wire _66862 = uncoded_block[550] ^ uncoded_block[600];
  wire _66863 = _66861 ^ _66862;
  wire _66864 = uncoded_block[602] ^ uncoded_block[660];
  wire _66865 = uncoded_block[666] ^ uncoded_block[682];
  wire _66866 = _66864 ^ _66865;
  wire _66867 = _66863 ^ _66866;
  wire _66868 = uncoded_block[738] ^ uncoded_block[776];
  wire _66869 = _1200 ^ _66868;
  wire _66870 = uncoded_block[791] ^ uncoded_block[821];
  wire _66871 = _66870 ^ _52862;
  wire _66872 = _66869 ^ _66871;
  wire _66873 = _66867 ^ _66872;
  wire _66874 = _66860 ^ _66873;
  wire _66875 = uncoded_block[898] ^ uncoded_block[943];
  wire _66876 = uncoded_block[952] ^ uncoded_block[1002];
  wire _66877 = _66875 ^ _66876;
  wire _66878 = uncoded_block[1006] ^ uncoded_block[1032];
  wire _66879 = uncoded_block[1100] ^ uncoded_block[1162];
  wire _66880 = _66878 ^ _66879;
  wire _66881 = _66877 ^ _66880;
  wire _66882 = uncoded_block[1163] ^ uncoded_block[1203];
  wire _66883 = uncoded_block[1217] ^ uncoded_block[1274];
  wire _66884 = _66882 ^ _66883;
  wire _66885 = uncoded_block[1281] ^ uncoded_block[1299];
  wire _66886 = uncoded_block[1308] ^ uncoded_block[1355];
  wire _66887 = _66885 ^ _66886;
  wire _66888 = _66884 ^ _66887;
  wire _66889 = _66881 ^ _66888;
  wire _66890 = uncoded_block[1368] ^ uncoded_block[1397];
  wire _66891 = uncoded_block[1414] ^ uncoded_block[1470];
  wire _66892 = _66890 ^ _66891;
  wire _66893 = uncoded_block[1507] ^ uncoded_block[1525];
  wire _66894 = uncoded_block[1563] ^ uncoded_block[1578];
  wire _66895 = _66893 ^ _66894;
  wire _66896 = _66892 ^ _66895;
  wire _66897 = uncoded_block[1580] ^ uncoded_block[1640];
  wire _66898 = _66897 ^ _6691;
  wire _66899 = _66898 ^ uncoded_block[1672];
  wire _66900 = _66896 ^ _66899;
  wire _66901 = _66889 ^ _66900;
  wire _66902 = _66874 ^ _66901;
  wire _66903 = uncoded_block[27] ^ uncoded_block[41];
  wire _66904 = uncoded_block[49] ^ uncoded_block[80];
  wire _66905 = _66903 ^ _66904;
  wire _66906 = uncoded_block[113] ^ uncoded_block[138];
  wire _66907 = _58997 ^ _66906;
  wire _66908 = _66905 ^ _66907;
  wire _66909 = uncoded_block[170] ^ uncoded_block[182];
  wire _66910 = uncoded_block[191] ^ uncoded_block[223];
  wire _66911 = _66909 ^ _66910;
  wire _66912 = uncoded_block[293] ^ uncoded_block[302];
  wire _66913 = _9222 ^ _66912;
  wire _66914 = _66911 ^ _66913;
  wire _66915 = _66908 ^ _66914;
  wire _66916 = uncoded_block[321] ^ uncoded_block[346];
  wire _66917 = uncoded_block[354] ^ uncoded_block[369];
  wire _66918 = _66916 ^ _66917;
  wire _66919 = uncoded_block[400] ^ uncoded_block[435];
  wire _66920 = uncoded_block[437] ^ uncoded_block[467];
  wire _66921 = _66919 ^ _66920;
  wire _66922 = _66918 ^ _66921;
  wire _66923 = _9832 ^ _19638;
  wire _66924 = uncoded_block[544] ^ uncoded_block[573];
  wire _66925 = uncoded_block[593] ^ uncoded_block[614];
  wire _66926 = _66924 ^ _66925;
  wire _66927 = _66923 ^ _66926;
  wire _66928 = _66922 ^ _66927;
  wire _66929 = _66915 ^ _66928;
  wire _66930 = uncoded_block[663] ^ uncoded_block[681];
  wire _66931 = _62205 ^ _66930;
  wire _66932 = uncoded_block[739] ^ uncoded_block[750];
  wire _66933 = _51599 ^ _66932;
  wire _66934 = _66931 ^ _66933;
  wire _66935 = uncoded_block[821] ^ uncoded_block[855];
  wire _66936 = _8793 ^ _66935;
  wire _66937 = uncoded_block[902] ^ uncoded_block[929];
  wire _66938 = _59108 ^ _66937;
  wire _66939 = _66936 ^ _66938;
  wire _66940 = _66934 ^ _66939;
  wire _66941 = uncoded_block[936] ^ uncoded_block[951];
  wire _66942 = uncoded_block[962] ^ uncoded_block[992];
  wire _66943 = _66941 ^ _66942;
  wire _66944 = uncoded_block[1019] ^ uncoded_block[1050];
  wire _66945 = uncoded_block[1089] ^ uncoded_block[1101];
  wire _66946 = _66944 ^ _66945;
  wire _66947 = _66943 ^ _66946;
  wire _66948 = uncoded_block[1104] ^ uncoded_block[1116];
  wire _66949 = uncoded_block[1129] ^ uncoded_block[1154];
  wire _66950 = _66948 ^ _66949;
  wire _66951 = uncoded_block[1182] ^ uncoded_block[1206];
  wire _66952 = _37388 ^ _66951;
  wire _66953 = _66950 ^ _66952;
  wire _66954 = _66947 ^ _66953;
  wire _66955 = _66940 ^ _66954;
  wire _66956 = _66929 ^ _66955;
  wire _66957 = uncoded_block[1212] ^ uncoded_block[1237];
  wire _66958 = uncoded_block[1253] ^ uncoded_block[1261];
  wire _66959 = _66957 ^ _66958;
  wire _66960 = uncoded_block[1278] ^ uncoded_block[1287];
  wire _66961 = _66960 ^ _34168;
  wire _66962 = _66959 ^ _66961;
  wire _66963 = _38205 ^ _49438;
  wire _66964 = uncoded_block[1467] ^ uncoded_block[1499];
  wire _66965 = _65248 ^ _66964;
  wire _66966 = _66963 ^ _66965;
  wire _66967 = _66962 ^ _66966;
  wire _66968 = uncoded_block[1504] ^ uncoded_block[1533];
  wire _66969 = uncoded_block[1544] ^ uncoded_block[1580];
  wire _66970 = _66968 ^ _66969;
  wire _66971 = uncoded_block[1641] ^ uncoded_block[1653];
  wire _66972 = _16031 ^ _66971;
  wire _66973 = _66970 ^ _66972;
  wire _66974 = _3976 ^ uncoded_block[1708];
  wire _66975 = _66973 ^ _66974;
  wire _66976 = _66967 ^ _66975;
  wire _66977 = _66956 ^ _66976;
  wire _66978 = uncoded_block[11] ^ uncoded_block[35];
  wire _66979 = uncoded_block[40] ^ uncoded_block[70];
  wire _66980 = _66978 ^ _66979;
  wire _66981 = uncoded_block[84] ^ uncoded_block[108];
  wire _66982 = uncoded_block[127] ^ uncoded_block[158];
  wire _66983 = _66981 ^ _66982;
  wire _66984 = _66980 ^ _66983;
  wire _66985 = uncoded_block[159] ^ uncoded_block[187];
  wire _66986 = uncoded_block[193] ^ uncoded_block[206];
  wire _66987 = _66985 ^ _66986;
  wire _66988 = uncoded_block[256] ^ uncoded_block[260];
  wire _66989 = uncoded_block[274] ^ uncoded_block[288];
  wire _66990 = _66988 ^ _66989;
  wire _66991 = _66987 ^ _66990;
  wire _66992 = _66984 ^ _66991;
  wire _66993 = uncoded_block[298] ^ uncoded_block[325];
  wire _66994 = _66993 ^ _4141;
  wire _66995 = uncoded_block[408] ^ uncoded_block[426];
  wire _66996 = _16671 ^ _66995;
  wire _66997 = _66994 ^ _66996;
  wire _66998 = uncoded_block[496] ^ uncoded_block[532];
  wire _66999 = _12578 ^ _66998;
  wire _67000 = uncoded_block[544] ^ uncoded_block[553];
  wire _67001 = _67000 ^ _9319;
  wire _67002 = _66999 ^ _67001;
  wire _67003 = _66997 ^ _67002;
  wire _67004 = _66992 ^ _67003;
  wire _67005 = uncoded_block[590] ^ uncoded_block[631];
  wire _67006 = uncoded_block[662] ^ uncoded_block[672];
  wire _67007 = _67005 ^ _67006;
  wire _67008 = uncoded_block[724] ^ uncoded_block[772];
  wire _67009 = _50516 ^ _67008;
  wire _67010 = _67007 ^ _67009;
  wire _67011 = uncoded_block[774] ^ uncoded_block[802];
  wire _67012 = uncoded_block[814] ^ uncoded_block[827];
  wire _67013 = _67011 ^ _67012;
  wire _67014 = uncoded_block[844] ^ uncoded_block[863];
  wire _67015 = uncoded_block[869] ^ uncoded_block[888];
  wire _67016 = _67014 ^ _67015;
  wire _67017 = _67013 ^ _67016;
  wire _67018 = _67010 ^ _67017;
  wire _67019 = uncoded_block[913] ^ uncoded_block[930];
  wire _67020 = uncoded_block[949] ^ uncoded_block[965];
  wire _67021 = _67019 ^ _67020;
  wire _67022 = uncoded_block[970] ^ uncoded_block[1009];
  wire _67023 = uncoded_block[1010] ^ uncoded_block[1040];
  wire _67024 = _67022 ^ _67023;
  wire _67025 = _67021 ^ _67024;
  wire _67026 = uncoded_block[1076] ^ uncoded_block[1091];
  wire _67027 = uncoded_block[1094] ^ uncoded_block[1146];
  wire _67028 = _67026 ^ _67027;
  wire _67029 = uncoded_block[1156] ^ uncoded_block[1167];
  wire _67030 = uncoded_block[1192] ^ uncoded_block[1200];
  wire _67031 = _67029 ^ _67030;
  wire _67032 = _67028 ^ _67031;
  wire _67033 = _67025 ^ _67032;
  wire _67034 = _67018 ^ _67033;
  wire _67035 = _67004 ^ _67034;
  wire _67036 = uncoded_block[1217] ^ uncoded_block[1240];
  wire _67037 = uncoded_block[1253] ^ uncoded_block[1265];
  wire _67038 = _67036 ^ _67037;
  wire _67039 = uncoded_block[1276] ^ uncoded_block[1300];
  wire _67040 = uncoded_block[1306] ^ uncoded_block[1315];
  wire _67041 = _67039 ^ _67040;
  wire _67042 = _67038 ^ _67041;
  wire _67043 = uncoded_block[1349] ^ uncoded_block[1361];
  wire _67044 = uncoded_block[1392] ^ uncoded_block[1405];
  wire _67045 = _67043 ^ _67044;
  wire _67046 = uncoded_block[1437] ^ uncoded_block[1496];
  wire _67047 = uncoded_block[1513] ^ uncoded_block[1534];
  wire _67048 = _67046 ^ _67047;
  wire _67049 = _67045 ^ _67048;
  wire _67050 = _67042 ^ _67049;
  wire _67051 = uncoded_block[1544] ^ uncoded_block[1559];
  wire _67052 = uncoded_block[1565] ^ uncoded_block[1579];
  wire _67053 = _67051 ^ _67052;
  wire _67054 = _60917 ^ _17020;
  wire _67055 = _67053 ^ _67054;
  wire _67056 = uncoded_block[1645] ^ uncoded_block[1680];
  wire _67057 = _67056 ^ uncoded_block[1714];
  wire _67058 = _67055 ^ _67057;
  wire _67059 = _67050 ^ _67058;
  wire _67060 = _67035 ^ _67059;
  wire _67061 = _64628 ^ _20453;
  wire _67062 = uncoded_block[41] ^ uncoded_block[68];
  wire _67063 = _67062 ^ _10246;
  wire _67064 = _67061 ^ _67063;
  wire _67065 = uncoded_block[118] ^ uncoded_block[123];
  wire _67066 = _67065 ^ _57605;
  wire _67067 = uncoded_block[189] ^ uncoded_block[212];
  wire _67068 = _59935 ^ _67067;
  wire _67069 = _67066 ^ _67068;
  wire _67070 = _67064 ^ _67069;
  wire _67071 = uncoded_block[233] ^ uncoded_block[251];
  wire _67072 = uncoded_block[257] ^ uncoded_block[288];
  wire _67073 = _67071 ^ _67072;
  wire _67074 = _964 ^ _67073;
  wire _67075 = uncoded_block[313] ^ uncoded_block[326];
  wire _67076 = _57627 ^ _67075;
  wire _67077 = _52744 ^ _59962;
  wire _67078 = _67076 ^ _67077;
  wire _67079 = _67074 ^ _67078;
  wire _67080 = _67070 ^ _67079;
  wire _67081 = uncoded_block[382] ^ uncoded_block[413];
  wire _67082 = uncoded_block[416] ^ uncoded_block[425];
  wire _67083 = _67081 ^ _67082;
  wire _67084 = _4174 ^ _59466;
  wire _67085 = _67083 ^ _67084;
  wire _67086 = uncoded_block[471] ^ uncoded_block[499];
  wire _67087 = uncoded_block[504] ^ uncoded_block[530];
  wire _67088 = _67086 ^ _67087;
  wire _67089 = uncoded_block[536] ^ uncoded_block[545];
  wire _67090 = _67089 ^ _44134;
  wire _67091 = _67088 ^ _67090;
  wire _67092 = _67085 ^ _67091;
  wire _67093 = uncoded_block[592] ^ uncoded_block[600];
  wire _67094 = _49541 ^ _67093;
  wire _67095 = _59988 ^ _21575;
  wire _67096 = _67094 ^ _67095;
  wire _67097 = uncoded_block[647] ^ uncoded_block[656];
  wire _67098 = uncoded_block[677] ^ uncoded_block[690];
  wire _67099 = _67097 ^ _67098;
  wire _67100 = uncoded_block[710] ^ uncoded_block[731];
  wire _67101 = _41180 ^ _67100;
  wire _67102 = _67099 ^ _67101;
  wire _67103 = _67096 ^ _67102;
  wire _67104 = _67092 ^ _67103;
  wire _67105 = _67080 ^ _67104;
  wire _67106 = _6377 ^ _364;
  wire _67107 = uncoded_block[790] ^ uncoded_block[806];
  wire _67108 = _67107 ^ _1239;
  wire _67109 = _67106 ^ _67108;
  wire _67110 = uncoded_block[826] ^ uncoded_block[847];
  wire _67111 = uncoded_block[848] ^ uncoded_block[873];
  wire _67112 = _67110 ^ _67111;
  wire _67113 = uncoded_block[874] ^ uncoded_block[883];
  wire _67114 = uncoded_block[897] ^ uncoded_block[909];
  wire _67115 = _67113 ^ _67114;
  wire _67116 = _67112 ^ _67115;
  wire _67117 = _67109 ^ _67116;
  wire _67118 = uncoded_block[919] ^ uncoded_block[931];
  wire _67119 = uncoded_block[936] ^ uncoded_block[967];
  wire _67120 = _67118 ^ _67119;
  wire _67121 = uncoded_block[977] ^ uncoded_block[985];
  wire _67122 = _67121 ^ _28985;
  wire _67123 = _67120 ^ _67122;
  wire _67124 = uncoded_block[1021] ^ uncoded_block[1030];
  wire _67125 = _8868 ^ _67124;
  wire _67126 = uncoded_block[1064] ^ uncoded_block[1071];
  wire _67127 = uncoded_block[1074] ^ uncoded_block[1107];
  wire _67128 = _67126 ^ _67127;
  wire _67129 = _67125 ^ _67128;
  wire _67130 = _67123 ^ _67129;
  wire _67131 = _67117 ^ _67130;
  wire _67132 = uncoded_block[1109] ^ uncoded_block[1122];
  wire _67133 = _67132 ^ _7737;
  wire _67134 = uncoded_block[1165] ^ uncoded_block[1173];
  wire _67135 = _45022 ^ _67134;
  wire _67136 = _67133 ^ _67135;
  wire _67137 = uncoded_block[1175] ^ uncoded_block[1197];
  wire _67138 = _67137 ^ _49584;
  wire _67139 = uncoded_block[1226] ^ uncoded_block[1249];
  wire _67140 = uncoded_block[1252] ^ uncoded_block[1261];
  wire _67141 = _67139 ^ _67140;
  wire _67142 = _67138 ^ _67141;
  wire _67143 = _67136 ^ _67142;
  wire _67144 = uncoded_block[1266] ^ uncoded_block[1294];
  wire _67145 = _67144 ^ _60071;
  wire _67146 = uncoded_block[1327] ^ uncoded_block[1341];
  wire _67147 = uncoded_block[1365] ^ uncoded_block[1385];
  wire _67148 = _67146 ^ _67147;
  wire _67149 = _67145 ^ _67148;
  wire _67150 = _10678 ^ _20355;
  wire _67151 = _2329 ^ _64604;
  wire _67152 = _67150 ^ _67151;
  wire _67153 = _67149 ^ _67152;
  wire _67154 = _67143 ^ _67153;
  wire _67155 = _67131 ^ _67154;
  wire _67156 = _67105 ^ _67155;
  wire _67157 = uncoded_block[1552] ^ uncoded_block[1565];
  wire _67158 = _60098 ^ _67157;
  wire _67159 = _67158 ^ _44378;
  wire _67160 = uncoded_block[1594] ^ uncoded_block[1628];
  wire _67161 = _67160 ^ _3166;
  wire _67162 = uncoded_block[1663] ^ uncoded_block[1683];
  wire _67163 = _36687 ^ _67162;
  wire _67164 = _67161 ^ _67163;
  wire _67165 = _67159 ^ _67164;
  wire _67166 = _3976 ^ uncoded_block[1715];
  wire _67167 = _67165 ^ _67166;
  wire _67168 = _67156 ^ _67167;
  wire _67169 = uncoded_block[7] ^ uncoded_block[19];
  wire _67170 = uncoded_block[46] ^ uncoded_block[76];
  wire _67171 = _67169 ^ _67170;
  wire _67172 = uncoded_block[89] ^ uncoded_block[99];
  wire _67173 = _67172 ^ _60487;
  wire _67174 = _67171 ^ _67173;
  wire _67175 = uncoded_block[137] ^ uncoded_block[176];
  wire _67176 = _67175 ^ _60493;
  wire _67177 = uncoded_block[251] ^ uncoded_block[257];
  wire _67178 = uncoded_block[261] ^ uncoded_block[282];
  wire _67179 = _67177 ^ _67178;
  wire _67180 = _67176 ^ _67179;
  wire _67181 = _67174 ^ _67180;
  wire _67182 = uncoded_block[350] ^ uncoded_block[356];
  wire _67183 = _8632 ^ _67182;
  wire _67184 = uncoded_block[376] ^ uncoded_block[402];
  wire _67185 = uncoded_block[404] ^ uncoded_block[422];
  wire _67186 = _67184 ^ _67185;
  wire _67187 = _67183 ^ _67186;
  wire _67188 = uncoded_block[450] ^ uncoded_block[467];
  wire _67189 = uncoded_block[496] ^ uncoded_block[517];
  wire _67190 = _67188 ^ _67189;
  wire _67191 = uncoded_block[533] ^ uncoded_block[540];
  wire _67192 = uncoded_block[566] ^ uncoded_block[601];
  wire _67193 = _67191 ^ _67192;
  wire _67194 = _67190 ^ _67193;
  wire _67195 = _67187 ^ _67194;
  wire _67196 = _67181 ^ _67195;
  wire _67197 = uncoded_block[612] ^ uncoded_block[635];
  wire _67198 = _67197 ^ _9885;
  wire _67199 = uncoded_block[673] ^ uncoded_block[686];
  wire _67200 = uncoded_block[715] ^ uncoded_block[746];
  wire _67201 = _67199 ^ _67200;
  wire _67202 = _67198 ^ _67201;
  wire _67203 = _60534 ^ _56506;
  wire _67204 = uncoded_block[835] ^ uncoded_block[867];
  wire _67205 = _60540 ^ _67204;
  wire _67206 = _67203 ^ _67205;
  wire _67207 = _67202 ^ _67206;
  wire _67208 = uncoded_block[925] ^ uncoded_block[949];
  wire _67209 = _6428 ^ _67208;
  wire _67210 = uncoded_block[968] ^ uncoded_block[993];
  wire _67211 = _67210 ^ _35710;
  wire _67212 = _67209 ^ _67211;
  wire _67213 = uncoded_block[1049] ^ uncoded_block[1067];
  wire _67214 = _67213 ^ _36955;
  wire _67215 = uncoded_block[1140] ^ uncoded_block[1150];
  wire _67216 = _67215 ^ _60567;
  wire _67217 = _67214 ^ _67216;
  wire _67218 = _67212 ^ _67217;
  wire _67219 = _67207 ^ _67218;
  wire _67220 = _67196 ^ _67219;
  wire _67221 = uncoded_block[1202] ^ uncoded_block[1238];
  wire _67222 = uncoded_block[1246] ^ uncoded_block[1270];
  wire _67223 = _67221 ^ _67222;
  wire _67224 = uncoded_block[1290] ^ uncoded_block[1313];
  wire _67225 = _2248 ^ _67224;
  wire _67226 = _67223 ^ _67225;
  wire _67227 = _54498 ^ _60586;
  wire _67228 = uncoded_block[1464] ^ uncoded_block[1536];
  wire _67229 = _67228 ^ _60596;
  wire _67230 = _67227 ^ _67229;
  wire _67231 = _67226 ^ _67230;
  wire _67232 = uncoded_block[1564] ^ uncoded_block[1592];
  wire _67233 = _57554 ^ _67232;
  wire _67234 = uncoded_block[1607] ^ uncoded_block[1625];
  wire _67235 = _67234 ^ _12947;
  wire _67236 = _67233 ^ _67235;
  wire _67237 = _67236 ^ uncoded_block[1649];
  wire _67238 = _67231 ^ _67237;
  wire _67239 = _67220 ^ _67238;
  wire _67240 = uncoded_block[1] ^ uncoded_block[44];
  wire _67241 = _67240 ^ _17067;
  wire _67242 = uncoded_block[59] ^ uncoded_block[64];
  wire _67243 = _67242 ^ _63558;
  wire _67244 = _67241 ^ _67243;
  wire _67245 = uncoded_block[148] ^ uncoded_block[153];
  wire _67246 = _48814 ^ _67245;
  wire _67247 = _65752 ^ _52383;
  wire _67248 = _67246 ^ _67247;
  wire _67249 = _67244 ^ _67248;
  wire _67250 = uncoded_block[248] ^ uncoded_block[270];
  wire _67251 = _60765 ^ _67250;
  wire _67252 = uncoded_block[280] ^ uncoded_block[300];
  wire _67253 = _67252 ^ _57843;
  wire _67254 = _67251 ^ _67253;
  wire _67255 = uncoded_block[350] ^ uncoded_block[365];
  wire _67256 = _67255 ^ _6879;
  wire _67257 = uncoded_block[416] ^ uncoded_block[468];
  wire _67258 = _5559 ^ _67257;
  wire _67259 = _67256 ^ _67258;
  wire _67260 = _67254 ^ _67259;
  wire _67261 = _67249 ^ _67260;
  wire _67262 = uncoded_block[486] ^ uncoded_block[509];
  wire _67263 = _28866 ^ _67262;
  wire _67264 = uncoded_block[522] ^ uncoded_block[529];
  wire _67265 = uncoded_block[554] ^ uncoded_block[591];
  wire _67266 = _67264 ^ _67265;
  wire _67267 = _67263 ^ _67266;
  wire _67268 = uncoded_block[592] ^ uncoded_block[607];
  wire _67269 = uncoded_block[624] ^ uncoded_block[659];
  wire _67270 = _67268 ^ _67269;
  wire _67271 = uncoded_block[681] ^ uncoded_block[697];
  wire _67272 = _308 ^ _67271;
  wire _67273 = _67270 ^ _67272;
  wire _67274 = _67267 ^ _67273;
  wire _67275 = uncoded_block[699] ^ uncoded_block[719];
  wire _67276 = _67275 ^ _49300;
  wire _67277 = uncoded_block[757] ^ uncoded_block[769];
  wire _67278 = uncoded_block[778] ^ uncoded_block[790];
  wire _67279 = _67277 ^ _67278;
  wire _67280 = _67276 ^ _67279;
  wire _67281 = uncoded_block[791] ^ uncoded_block[804];
  wire _67282 = uncoded_block[830] ^ uncoded_block[846];
  wire _67283 = _67281 ^ _67282;
  wire _67284 = uncoded_block[869] ^ uncoded_block[889];
  wire _67285 = _6410 ^ _67284;
  wire _67286 = _67283 ^ _67285;
  wire _67287 = _67280 ^ _67286;
  wire _67288 = _67274 ^ _67287;
  wire _67289 = _67261 ^ _67288;
  wire _67290 = uncoded_block[921] ^ uncoded_block[931];
  wire _67291 = uncoded_block[934] ^ uncoded_block[970];
  wire _67292 = _67290 ^ _67291;
  wire _67293 = uncoded_block[971] ^ uncoded_block[982];
  wire _67294 = uncoded_block[998] ^ uncoded_block[1009];
  wire _67295 = _67293 ^ _67294;
  wire _67296 = _67292 ^ _67295;
  wire _67297 = uncoded_block[1016] ^ uncoded_block[1030];
  wire _67298 = uncoded_block[1043] ^ uncoded_block[1063];
  wire _67299 = _67297 ^ _67298;
  wire _67300 = uncoded_block[1069] ^ uncoded_block[1078];
  wire _67301 = uncoded_block[1083] ^ uncoded_block[1130];
  wire _67302 = _67300 ^ _67301;
  wire _67303 = _67299 ^ _67302;
  wire _67304 = _67296 ^ _67303;
  wire _67305 = uncoded_block[1161] ^ uncoded_block[1167];
  wire _67306 = _7743 ^ _67305;
  wire _67307 = uncoded_block[1209] ^ uncoded_block[1217];
  wire _67308 = _61017 ^ _67307;
  wire _67309 = _67306 ^ _67308;
  wire _67310 = uncoded_block[1224] ^ uncoded_block[1231];
  wire _67311 = uncoded_block[1236] ^ uncoded_block[1263];
  wire _67312 = _67310 ^ _67311;
  wire _67313 = uncoded_block[1271] ^ uncoded_block[1285];
  wire _67314 = uncoded_block[1299] ^ uncoded_block[1320];
  wire _67315 = _67313 ^ _67314;
  wire _67316 = _67312 ^ _67315;
  wire _67317 = _67309 ^ _67316;
  wire _67318 = _67304 ^ _67317;
  wire _67319 = uncoded_block[1322] ^ uncoded_block[1333];
  wire _67320 = uncoded_block[1338] ^ uncoded_block[1376];
  wire _67321 = _67319 ^ _67320;
  wire _67322 = uncoded_block[1395] ^ uncoded_block[1435];
  wire _67323 = _3058 ^ _67322;
  wire _67324 = _67321 ^ _67323;
  wire _67325 = uncoded_block[1474] ^ uncoded_block[1494];
  wire _67326 = uncoded_block[1543] ^ uncoded_block[1548];
  wire _67327 = _67325 ^ _67326;
  wire _67328 = uncoded_block[1550] ^ uncoded_block[1571];
  wire _67329 = _67328 ^ _34240;
  wire _67330 = _67327 ^ _67329;
  wire _67331 = _67324 ^ _67330;
  wire _67332 = uncoded_block[1591] ^ uncoded_block[1604];
  wire _67333 = uncoded_block[1634] ^ uncoded_block[1642];
  wire _67334 = _67332 ^ _67333;
  wire _67335 = uncoded_block[1684] ^ uncoded_block[1703];
  wire _67336 = _8522 ^ _67335;
  wire _67337 = _67334 ^ _67336;
  wire _67338 = _67337 ^ uncoded_block[1710];
  wire _67339 = _67331 ^ _67338;
  wire _67340 = _67318 ^ _67339;
  wire _67341 = _67289 ^ _67340;
  wire _67342 = uncoded_block[26] ^ uncoded_block[50];
  wire _67343 = uncoded_block[55] ^ uncoded_block[100];
  wire _67344 = _67342 ^ _67343;
  wire _67345 = uncoded_block[115] ^ uncoded_block[137];
  wire _67346 = uncoded_block[171] ^ uncoded_block[181];
  wire _67347 = _67345 ^ _67346;
  wire _67348 = _67344 ^ _67347;
  wire _67349 = uncoded_block[245] ^ uncoded_block[275];
  wire _67350 = uncoded_block[304] ^ uncoded_block[320];
  wire _67351 = _67349 ^ _67350;
  wire _67352 = uncoded_block[353] ^ uncoded_block[371];
  wire _67353 = uncoded_block[401] ^ uncoded_block[436];
  wire _67354 = _67352 ^ _67353;
  wire _67355 = _67351 ^ _67354;
  wire _67356 = _67348 ^ _67355;
  wire _67357 = uncoded_block[517] ^ uncoded_block[546];
  wire _67358 = _9291 ^ _67357;
  wire _67359 = uncoded_block[572] ^ uncoded_block[595];
  wire _67360 = uncoded_block[642] ^ uncoded_block[662];
  wire _67361 = _67359 ^ _67360;
  wire _67362 = _67358 ^ _67361;
  wire _67363 = uncoded_block[749] ^ uncoded_block[803];
  wire _67364 = _27413 ^ _67363;
  wire _67365 = uncoded_block[823] ^ uncoded_block[881];
  wire _67366 = uncoded_block[928] ^ uncoded_block[938];
  wire _67367 = _67365 ^ _67366;
  wire _67368 = _67364 ^ _67367;
  wire _67369 = _67362 ^ _67368;
  wire _67370 = _67356 ^ _67369;
  wire _67371 = uncoded_block[1018] ^ uncoded_block[1052];
  wire _67372 = _65705 ^ _67371;
  wire _67373 = uncoded_block[1088] ^ uncoded_block[1106];
  wire _67374 = uncoded_block[1118] ^ uncoded_block[1128];
  wire _67375 = _67373 ^ _67374;
  wire _67376 = _67372 ^ _67375;
  wire _67377 = uncoded_block[1164] ^ uncoded_block[1208];
  wire _67378 = _67377 ^ _57736;
  wire _67379 = _64577 ^ _1468;
  wire _67380 = _67378 ^ _67379;
  wire _67381 = _67376 ^ _67380;
  wire _67382 = uncoded_block[1412] ^ uncoded_block[1418];
  wire _67383 = _40945 ^ _67382;
  wire _67384 = uncoded_block[1499] ^ uncoded_block[1583];
  wire _67385 = _58934 ^ _67384;
  wire _67386 = _67383 ^ _67385;
  wire _67387 = uncoded_block[1585] ^ uncoded_block[1616];
  wire _67388 = uncoded_block[1640] ^ uncoded_block[1654];
  wire _67389 = _67387 ^ _67388;
  wire _67390 = _67389 ^ uncoded_block[1684];
  wire _67391 = _67386 ^ _67390;
  wire _67392 = _67381 ^ _67391;
  wire _67393 = _67370 ^ _67392;
  wire _67394 = uncoded_block[19] ^ uncoded_block[40];
  wire _67395 = _67394 ^ _61254;
  wire _67396 = uncoded_block[79] ^ uncoded_block[107];
  wire _67397 = uncoded_block[128] ^ uncoded_block[167];
  wire _67398 = _67396 ^ _67397;
  wire _67399 = _67395 ^ _67398;
  wire _67400 = uncoded_block[170] ^ uncoded_block[190];
  wire _67401 = _67400 ^ _6800;
  wire _67402 = uncoded_block[243] ^ uncoded_block[265];
  wire _67403 = _67402 ^ _61268;
  wire _67404 = _67401 ^ _67403;
  wire _67405 = _67399 ^ _67404;
  wire _67406 = _35929 ^ _11987;
  wire _67407 = uncoded_block[385] ^ uncoded_block[433];
  wire _67408 = uncoded_block[435] ^ uncoded_block[440];
  wire _67409 = _67407 ^ _67408;
  wire _67410 = _67406 ^ _67409;
  wire _67411 = uncoded_block[456] ^ uncoded_block[466];
  wire _67412 = uncoded_block[501] ^ uncoded_block[518];
  wire _67413 = _67411 ^ _67412;
  wire _67414 = _61289 ^ _6310;
  wire _67415 = _67413 ^ _67414;
  wire _67416 = _67410 ^ _67415;
  wire _67417 = _67405 ^ _67416;
  wire _67418 = uncoded_block[612] ^ uncoded_block[639];
  wire _67419 = _67418 ^ _65621;
  wire _67420 = uncoded_block[680] ^ uncoded_block[709];
  wire _67421 = _67420 ^ _61308;
  wire _67422 = _67419 ^ _67421;
  wire _67423 = uncoded_block[737] ^ uncoded_block[761];
  wire _67424 = uncoded_block[794] ^ uncoded_block[805];
  wire _67425 = _67423 ^ _67424;
  wire _67426 = uncoded_block[822] ^ uncoded_block[857];
  wire _67427 = uncoded_block[869] ^ uncoded_block[877];
  wire _67428 = _67426 ^ _67427;
  wire _67429 = _67425 ^ _67428;
  wire _67430 = _67422 ^ _67429;
  wire _67431 = uncoded_block[900] ^ uncoded_block[958];
  wire _67432 = _56807 ^ _67431;
  wire _67433 = uncoded_block[991] ^ uncoded_block[1001];
  wire _67434 = uncoded_block[1036] ^ uncoded_block[1049];
  wire _67435 = _67433 ^ _67434;
  wire _67436 = _67432 ^ _67435;
  wire _67437 = uncoded_block[1057] ^ uncoded_block[1072];
  wire _67438 = _67437 ^ _5846;
  wire _67439 = _6507 ^ _11163;
  wire _67440 = _67438 ^ _67439;
  wire _67441 = _67436 ^ _67440;
  wire _67442 = _67430 ^ _67441;
  wire _67443 = _67417 ^ _67442;
  wire _67444 = uncoded_block[1259] ^ uncoded_block[1277];
  wire _67445 = _620 ^ _67444;
  wire _67446 = _61357 ^ _61359;
  wire _67447 = _67445 ^ _67446;
  wire _67448 = uncoded_block[1415] ^ uncoded_block[1442];
  wire _67449 = _61366 ^ _67448;
  wire _67450 = uncoded_block[1455] ^ uncoded_block[1485];
  wire _67451 = uncoded_block[1510] ^ uncoded_block[1518];
  wire _67452 = _67450 ^ _67451;
  wire _67453 = _67449 ^ _67452;
  wire _67454 = _67447 ^ _67453;
  wire _67455 = uncoded_block[1542] ^ uncoded_block[1579];
  wire _67456 = uncoded_block[1580] ^ uncoded_block[1605];
  wire _67457 = _67455 ^ _67456;
  wire _67458 = uncoded_block[1609] ^ uncoded_block[1623];
  wire _67459 = _67458 ^ _12960;
  wire _67460 = _67457 ^ _67459;
  wire _67461 = uncoded_block[1683] ^ uncoded_block[1689];
  wire _67462 = _67461 ^ uncoded_block[1707];
  wire _67463 = _67460 ^ _67462;
  wire _67464 = _67454 ^ _67463;
  wire _67465 = _67443 ^ _67464;
  wire _67466 = uncoded_block[1] ^ uncoded_block[19];
  wire _67467 = uncoded_block[23] ^ uncoded_block[68];
  wire _67468 = _67466 ^ _67467;
  wire _67469 = uncoded_block[76] ^ uncoded_block[100];
  wire _67470 = uncoded_block[101] ^ uncoded_block[126];
  wire _67471 = _67469 ^ _67470;
  wire _67472 = _67468 ^ _67471;
  wire _67473 = uncoded_block[152] ^ uncoded_block[178];
  wire _67474 = _58371 ^ _67473;
  wire _67475 = uncoded_block[193] ^ uncoded_block[198];
  wire _67476 = uncoded_block[223] ^ uncoded_block[239];
  wire _67477 = _67475 ^ _67476;
  wire _67478 = _67474 ^ _67477;
  wire _67479 = _67472 ^ _67478;
  wire _67480 = uncoded_block[240] ^ uncoded_block[248];
  wire _67481 = _67480 ^ _49516;
  wire _67482 = uncoded_block[291] ^ uncoded_block[315];
  wire _67483 = uncoded_block[322] ^ uncoded_block[363];
  wire _67484 = _67482 ^ _67483;
  wire _67485 = _67481 ^ _67484;
  wire _67486 = uncoded_block[365] ^ uncoded_block[375];
  wire _67487 = _67486 ^ _67184;
  wire _67488 = uncoded_block[429] ^ uncoded_block[467];
  wire _67489 = _14682 ^ _67488;
  wire _67490 = _67487 ^ _67489;
  wire _67491 = _67485 ^ _67490;
  wire _67492 = _67479 ^ _67491;
  wire _67493 = uncoded_block[486] ^ uncoded_block[514];
  wire _67494 = _59726 ^ _67493;
  wire _67495 = uncoded_block[541] ^ uncoded_block[587];
  wire _67496 = _60517 ^ _67495;
  wire _67497 = _67494 ^ _67496;
  wire _67498 = _14739 ^ _61829;
  wire _67499 = uncoded_block[643] ^ uncoded_block[697];
  wire _67500 = _290 ^ _67499;
  wire _67501 = _67498 ^ _67500;
  wire _67502 = _67497 ^ _67501;
  wire _67503 = uncoded_block[716] ^ uncoded_block[722];
  wire _67504 = _19201 ^ _67503;
  wire _67505 = uncoded_block[724] ^ uncoded_block[736];
  wire _67506 = uncoded_block[750] ^ uncoded_block[769];
  wire _67507 = _67505 ^ _67506;
  wire _67508 = _67504 ^ _67507;
  wire _67509 = _56506 ^ _12679;
  wire _67510 = uncoded_block[834] ^ uncoded_block[861];
  wire _67511 = _67510 ^ _423;
  wire _67512 = _67509 ^ _67511;
  wire _67513 = _67508 ^ _67512;
  wire _67514 = _67502 ^ _67513;
  wire _67515 = _67492 ^ _67514;
  wire _67516 = uncoded_block[925] ^ uncoded_block[934];
  wire _67517 = _12159 ^ _67516;
  wire _67518 = uncoded_block[968] ^ uncoded_block[980];
  wire _67519 = uncoded_block[981] ^ uncoded_block[998];
  wire _67520 = _67518 ^ _67519;
  wire _67521 = _67517 ^ _67520;
  wire _67522 = uncoded_block[1030] ^ uncoded_block[1048];
  wire _67523 = _18801 ^ _67522;
  wire _67524 = uncoded_block[1068] ^ uncoded_block[1083];
  wire _67525 = uncoded_block[1096] ^ uncoded_block[1121];
  wire _67526 = _67524 ^ _67525;
  wire _67527 = _67523 ^ _67526;
  wire _67528 = _67521 ^ _67527;
  wire _67529 = uncoded_block[1132] ^ uncoded_block[1140];
  wire _67530 = uncoded_block[1146] ^ uncoded_block[1167];
  wire _67531 = _67529 ^ _67530;
  wire _67532 = uncoded_block[1188] ^ uncoded_block[1209];
  wire _67533 = _67532 ^ _1440;
  wire _67534 = _67531 ^ _67533;
  wire _67535 = uncoded_block[1238] ^ uncoded_block[1267];
  wire _67536 = uncoded_block[1290] ^ uncoded_block[1296];
  wire _67537 = _67535 ^ _67536;
  wire _67538 = uncoded_block[1299] ^ uncoded_block[1307];
  wire _67539 = _67538 ^ _1495;
  wire _67540 = _67537 ^ _67539;
  wire _67541 = _67534 ^ _67540;
  wire _67542 = _67528 ^ _67541;
  wire _67543 = uncoded_block[1355] ^ uncoded_block[1366];
  wire _67544 = uncoded_block[1418] ^ uncoded_block[1444];
  wire _67545 = _67543 ^ _67544;
  wire _67546 = uncoded_block[1494] ^ uncoded_block[1506];
  wire _67547 = _5316 ^ _67546;
  wire _67548 = _67545 ^ _67547;
  wire _67549 = _65262 ^ _55416;
  wire _67550 = uncoded_block[1596] ^ uncoded_block[1611];
  wire _67551 = _3146 ^ _67550;
  wire _67552 = _67549 ^ _67551;
  wire _67553 = _67548 ^ _67552;
  wire _67554 = uncoded_block[1626] ^ uncoded_block[1649];
  wire _67555 = uncoded_block[1662] ^ uncoded_block[1687];
  wire _67556 = _67554 ^ _67555;
  wire _67557 = uncoded_block[1691] ^ uncoded_block[1710];
  wire _67558 = _67557 ^ uncoded_block[1719];
  wire _67559 = _67556 ^ _67558;
  wire _67560 = _67553 ^ _67559;
  wire _67561 = _67542 ^ _67560;
  wire _67562 = _67515 ^ _67561;
  wire _67563 = uncoded_block[2] ^ uncoded_block[45];
  wire _67564 = uncoded_block[54] ^ uncoded_block[102];
  wire _67565 = _67563 ^ _67564;
  wire _67566 = uncoded_block[134] ^ uncoded_block[169];
  wire _67567 = uncoded_block[195] ^ uncoded_block[204];
  wire _67568 = _67566 ^ _67567;
  wire _67569 = _67565 ^ _67568;
  wire _67570 = uncoded_block[300] ^ uncoded_block[328];
  wire _67571 = _5505 ^ _67570;
  wire _67572 = uncoded_block[350] ^ uncoded_block[387];
  wire _67573 = uncoded_block[406] ^ uncoded_block[425];
  wire _67574 = _67572 ^ _67573;
  wire _67575 = _67571 ^ _67574;
  wire _67576 = _67569 ^ _67575;
  wire _67577 = uncoded_block[532] ^ uncoded_block[554];
  wire _67578 = _60643 ^ _67577;
  wire _67579 = uncoded_block[570] ^ uncoded_block[582];
  wire _67580 = uncoded_block[628] ^ uncoded_block[647];
  wire _67581 = _67579 ^ _67580;
  wire _67582 = _67578 ^ _67581;
  wire _67583 = uncoded_block[678] ^ uncoded_block[711];
  wire _67584 = uncoded_block[760] ^ uncoded_block[772];
  wire _67585 = _67583 ^ _67584;
  wire _67586 = uncoded_block[820] ^ uncoded_block[829];
  wire _67587 = uncoded_block[840] ^ uncoded_block[856];
  wire _67588 = _67586 ^ _67587;
  wire _67589 = _67585 ^ _67588;
  wire _67590 = _67582 ^ _67589;
  wire _67591 = _67576 ^ _67590;
  wire _67592 = uncoded_block[919] ^ uncoded_block[929];
  wire _67593 = uncoded_block[946] ^ uncoded_block[1015];
  wire _67594 = _67592 ^ _67593;
  wire _67595 = uncoded_block[1024] ^ uncoded_block[1061];
  wire _67596 = uncoded_block[1092] ^ uncoded_block[1134];
  wire _67597 = _67595 ^ _67596;
  wire _67598 = _67594 ^ _67597;
  wire _67599 = uncoded_block[1139] ^ uncoded_block[1184];
  wire _67600 = uncoded_block[1210] ^ uncoded_block[1241];
  wire _67601 = _67599 ^ _67600;
  wire _67602 = uncoded_block[1272] ^ uncoded_block[1324];
  wire _67603 = _67602 ^ _60708;
  wire _67604 = _67601 ^ _67603;
  wire _67605 = _67598 ^ _67604;
  wire _67606 = uncoded_block[1356] ^ uncoded_block[1386];
  wire _67607 = _67606 ^ _8450;
  wire _67608 = uncoded_block[1486] ^ uncoded_block[1532];
  wire _67609 = uncoded_block[1576] ^ uncoded_block[1613];
  wire _67610 = _67608 ^ _67609;
  wire _67611 = _67607 ^ _67610;
  wire _67612 = uncoded_block[1647] ^ uncoded_block[1656];
  wire _67613 = uncoded_block[1685] ^ uncoded_block[1700];
  wire _67614 = _67612 ^ _67613;
  wire _67615 = _67614 ^ uncoded_block[1707];
  wire _67616 = _67611 ^ _67615;
  wire _67617 = _67605 ^ _67616;
  wire _67618 = _67591 ^ _67617;
  wire _67619 = uncoded_block[63] ^ uncoded_block[70];
  wire _67620 = _62454 ^ _67619;
  wire _67621 = uncoded_block[162] ^ uncoded_block[169];
  wire _67622 = _67621 ^ _60756;
  wire _67623 = _67620 ^ _67622;
  wire _67624 = uncoded_block[227] ^ uncoded_block[267];
  wire _67625 = uncoded_block[282] ^ uncoded_block[303];
  wire _67626 = _67624 ^ _67625;
  wire _67627 = _10907 ^ _4169;
  wire _67628 = _67626 ^ _67627;
  wire _67629 = _67623 ^ _67628;
  wire _67630 = uncoded_block[482] ^ uncoded_block[503];
  wire _67631 = uncoded_block[513] ^ uncoded_block[543];
  wire _67632 = _67630 ^ _67631;
  wire _67633 = uncoded_block[619] ^ uncoded_block[642];
  wire _67634 = _62506 ^ _67633;
  wire _67635 = _67632 ^ _67634;
  wire _67636 = uncoded_block[733] ^ uncoded_block[816];
  wire _67637 = _60818 ^ _67636;
  wire _67638 = uncoded_block[824] ^ uncoded_block[864];
  wire _67639 = uncoded_block[879] ^ uncoded_block[899];
  wire _67640 = _67638 ^ _67639;
  wire _67641 = _67637 ^ _67640;
  wire _67642 = _67635 ^ _67641;
  wire _67643 = _67629 ^ _67642;
  wire _67644 = uncoded_block[904] ^ uncoded_block[960];
  wire _67645 = uncoded_block[973] ^ uncoded_block[1036];
  wire _67646 = _67644 ^ _67645;
  wire _67647 = uncoded_block[1051] ^ uncoded_block[1066];
  wire _67648 = uncoded_block[1100] ^ uncoded_block[1159];
  wire _67649 = _67647 ^ _67648;
  wire _67650 = _67646 ^ _67649;
  wire _67651 = uncoded_block[1174] ^ uncoded_block[1195];
  wire _67652 = _67651 ^ _8958;
  wire _67653 = uncoded_block[1249] ^ uncoded_block[1312];
  wire _67654 = uncoded_block[1315] ^ uncoded_block[1332];
  wire _67655 = _67653 ^ _67654;
  wire _67656 = _67652 ^ _67655;
  wire _67657 = _67650 ^ _67656;
  wire _67658 = uncoded_block[1346] ^ uncoded_block[1358];
  wire _67659 = uncoded_block[1385] ^ uncoded_block[1415];
  wire _67660 = _67658 ^ _67659;
  wire _67661 = uncoded_block[1512] ^ uncoded_block[1541];
  wire _67662 = _62583 ^ _67661;
  wire _67663 = _67660 ^ _67662;
  wire _67664 = uncoded_block[1574] ^ uncoded_block[1625];
  wire _67665 = uncoded_block[1631] ^ uncoded_block[1690];
  wire _67666 = _67664 ^ _67665;
  wire _67667 = _67666 ^ uncoded_block[1710];
  wire _67668 = _67663 ^ _67667;
  wire _67669 = _67657 ^ _67668;
  wire _67670 = _67643 ^ _67669;
  wire _67671 = uncoded_block[4] ^ uncoded_block[47];
  wire _67672 = uncoded_block[87] ^ uncoded_block[105];
  wire _67673 = _67671 ^ _67672;
  wire _67674 = uncoded_block[111] ^ uncoded_block[148];
  wire _67675 = uncoded_block[208] ^ uncoded_block[215];
  wire _67676 = _67674 ^ _67675;
  wire _67677 = _67673 ^ _67676;
  wire _67678 = uncoded_block[254] ^ uncoded_block[267];
  wire _67679 = _67678 ^ _64891;
  wire _67680 = uncoded_block[415] ^ uncoded_block[438];
  wire _67681 = _57854 ^ _67680;
  wire _67682 = _67679 ^ _67681;
  wire _67683 = _67677 ^ _67682;
  wire _67684 = uncoded_block[526] ^ uncoded_block[552];
  wire _67685 = _60965 ^ _67684;
  wire _67686 = uncoded_block[573] ^ uncoded_block[599];
  wire _67687 = uncoded_block[625] ^ uncoded_block[666];
  wire _67688 = _67686 ^ _67687;
  wire _67689 = _67685 ^ _67688;
  wire _67690 = uncoded_block[692] ^ uncoded_block[711];
  wire _67691 = _67690 ^ _20156;
  wire _67692 = uncoded_block[780] ^ uncoded_block[789];
  wire _67693 = uncoded_block[841] ^ uncoded_block[859];
  wire _67694 = _67692 ^ _67693;
  wire _67695 = _67691 ^ _67694;
  wire _67696 = _67689 ^ _67695;
  wire _67697 = _67683 ^ _67696;
  wire _67698 = uncoded_block[977] ^ uncoded_block[997];
  wire _67699 = _45738 ^ _67698;
  wire _67700 = uncoded_block[1017] ^ uncoded_block[1057];
  wire _67701 = uncoded_block[1098] ^ uncoded_block[1114];
  wire _67702 = _67700 ^ _67701;
  wire _67703 = _67699 ^ _67702;
  wire _67704 = uncoded_block[1146] ^ uncoded_block[1179];
  wire _67705 = uncoded_block[1193] ^ uncoded_block[1258];
  wire _67706 = _67704 ^ _67705;
  wire _67707 = uncoded_block[1270] ^ uncoded_block[1306];
  wire _67708 = uncoded_block[1348] ^ uncoded_block[1372];
  wire _67709 = _67707 ^ _67708;
  wire _67710 = _67706 ^ _67709;
  wire _67711 = _67703 ^ _67710;
  wire _67712 = uncoded_block[1440] ^ uncoded_block[1483];
  wire _67713 = _65013 ^ _67712;
  wire _67714 = uncoded_block[1509] ^ uncoded_block[1527];
  wire _67715 = _27184 ^ _67714;
  wire _67716 = _67713 ^ _67715;
  wire _67717 = uncoded_block[1610] ^ uncoded_block[1670];
  wire _67718 = uncoded_block[1674] ^ uncoded_block[1689];
  wire _67719 = _67717 ^ _67718;
  wire _67720 = _67719 ^ uncoded_block[1717];
  wire _67721 = _67716 ^ _67720;
  wire _67722 = _67711 ^ _67721;
  wire _67723 = _67697 ^ _67722;
  wire _67724 = uncoded_block[29] ^ uncoded_block[41];
  wire _67725 = _67724 ^ _10246;
  wire _67726 = uncoded_block[129] ^ uncoded_block[155];
  wire _67727 = uncoded_block[203] ^ uncoded_block[213];
  wire _67728 = _67726 ^ _67727;
  wire _67729 = _67725 ^ _67728;
  wire _67730 = uncoded_block[231] ^ uncoded_block[262];
  wire _67731 = _67730 ^ _3332;
  wire _67732 = uncoded_block[347] ^ uncoded_block[376];
  wire _67733 = uncoded_block[399] ^ uncoded_block[433];
  wire _67734 = _67732 ^ _67733;
  wire _67735 = _67731 ^ _67734;
  wire _67736 = _67729 ^ _67735;
  wire _67737 = uncoded_block[466] ^ uncoded_block[507];
  wire _67738 = uncoded_block[509] ^ uncoded_block[590];
  wire _67739 = _67737 ^ _67738;
  wire _67740 = uncoded_block[616] ^ uncoded_block[652];
  wire _67741 = uncoded_block[660] ^ uncoded_block[679];
  wire _67742 = _67740 ^ _67741;
  wire _67743 = _67739 ^ _67742;
  wire _67744 = uncoded_block[694] ^ uncoded_block[751];
  wire _67745 = uncoded_block[758] ^ uncoded_block[788];
  wire _67746 = _67744 ^ _67745;
  wire _67747 = uncoded_block[812] ^ uncoded_block[843];
  wire _67748 = uncoded_block[872] ^ uncoded_block[916];
  wire _67749 = _67747 ^ _67748;
  wire _67750 = _67746 ^ _67749;
  wire _67751 = _67743 ^ _67750;
  wire _67752 = _67736 ^ _67751;
  wire _67753 = uncoded_block[918] ^ uncoded_block[957];
  wire _67754 = uncoded_block[980] ^ uncoded_block[1067];
  wire _67755 = _67753 ^ _67754;
  wire _67756 = uncoded_block[1077] ^ uncoded_block[1128];
  wire _67757 = uncoded_block[1149] ^ uncoded_block[1178];
  wire _67758 = _67756 ^ _67757;
  wire _67759 = _67755 ^ _67758;
  wire _67760 = uncoded_block[1192] ^ uncoded_block[1226];
  wire _67761 = uncoded_block[1268] ^ uncoded_block[1284];
  wire _67762 = _67760 ^ _67761;
  wire _67763 = uncoded_block[1314] ^ uncoded_block[1353];
  wire _67764 = uncoded_block[1377] ^ uncoded_block[1398];
  wire _67765 = _67763 ^ _67764;
  wire _67766 = _67762 ^ _67765;
  wire _67767 = _67759 ^ _67766;
  wire _67768 = uncoded_block[1453] ^ uncoded_block[1484];
  wire _67769 = _10690 ^ _67768;
  wire _67770 = uncoded_block[1487] ^ uncoded_block[1540];
  wire _67771 = uncoded_block[1553] ^ uncoded_block[1587];
  wire _67772 = _67770 ^ _67771;
  wire _67773 = _67769 ^ _67772;
  wire _67774 = uncoded_block[1639] ^ uncoded_block[1651];
  wire _67775 = uncoded_block[1672] ^ uncoded_block[1699];
  wire _67776 = _67774 ^ _67775;
  wire _67777 = _67776 ^ uncoded_block[1703];
  wire _67778 = _67773 ^ _67777;
  wire _67779 = _67767 ^ _67778;
  wire _67780 = _67752 ^ _67779;
  wire _67781 = uncoded_block[48] ^ uncoded_block[70];
  wire _67782 = _63165 ^ _67781;
  wire _67783 = uncoded_block[76] ^ uncoded_block[106];
  wire _67784 = _67783 ^ _3256;
  wire _67785 = _67782 ^ _67784;
  wire _67786 = uncoded_block[137] ^ uncoded_block[174];
  wire _67787 = uncoded_block[185] ^ uncoded_block[202];
  wire _67788 = _67786 ^ _67787;
  wire _67789 = uncoded_block[228] ^ uncoded_block[242];
  wire _67790 = uncoded_block[270] ^ uncoded_block[284];
  wire _67791 = _67789 ^ _67790;
  wire _67792 = _67788 ^ _67791;
  wire _67793 = _67785 ^ _67792;
  wire _67794 = _4125 ^ _37591;
  wire _67795 = uncoded_block[382] ^ uncoded_block[395];
  wire _67796 = uncoded_block[408] ^ uncoded_block[415];
  wire _67797 = _67795 ^ _67796;
  wire _67798 = _67794 ^ _67797;
  wire _67799 = uncoded_block[502] ^ uncoded_block[509];
  wire _67800 = _51559 ^ _67799;
  wire _67801 = uncoded_block[575] ^ uncoded_block[583];
  wire _67802 = _63228 ^ _67801;
  wire _67803 = _67800 ^ _67802;
  wire _67804 = _67798 ^ _67803;
  wire _67805 = _67793 ^ _67804;
  wire _67806 = uncoded_block[628] ^ uncoded_block[653];
  wire _67807 = _65501 ^ _67806;
  wire _67808 = uncoded_block[682] ^ uncoded_block[699];
  wire _67809 = uncoded_block[704] ^ uncoded_block[748];
  wire _67810 = _67808 ^ _67809;
  wire _67811 = _67807 ^ _67810;
  wire _67812 = uncoded_block[753] ^ uncoded_block[761];
  wire _67813 = uncoded_block[784] ^ uncoded_block[798];
  wire _67814 = _67812 ^ _67813;
  wire _67815 = uncoded_block[810] ^ uncoded_block[832];
  wire _67816 = uncoded_block[835] ^ uncoded_block[861];
  wire _67817 = _67815 ^ _67816;
  wire _67818 = _67814 ^ _67817;
  wire _67819 = _67811 ^ _67818;
  wire _67820 = uncoded_block[912] ^ uncoded_block[940];
  wire _67821 = uncoded_block[942] ^ uncoded_block[962];
  wire _67822 = _67820 ^ _67821;
  wire _67823 = uncoded_block[979] ^ uncoded_block[997];
  wire _67824 = uncoded_block[1012] ^ uncoded_block[1041];
  wire _67825 = _67823 ^ _67824;
  wire _67826 = _67822 ^ _67825;
  wire _67827 = uncoded_block[1045] ^ uncoded_block[1079];
  wire _67828 = _67827 ^ _61337;
  wire _67829 = uncoded_block[1123] ^ uncoded_block[1143];
  wire _67830 = _67829 ^ _9508;
  wire _67831 = _67828 ^ _67830;
  wire _67832 = _67826 ^ _67831;
  wire _67833 = _67819 ^ _67832;
  wire _67834 = _67805 ^ _67833;
  wire _67835 = uncoded_block[1205] ^ uncoded_block[1227];
  wire _67836 = uncoded_block[1257] ^ uncoded_block[1267];
  wire _67837 = _67835 ^ _67836;
  wire _67838 = uncoded_block[1300] ^ uncoded_block[1357];
  wire _67839 = _18417 ^ _67838;
  wire _67840 = _67837 ^ _67839;
  wire _67841 = uncoded_block[1390] ^ uncoded_block[1398];
  wire _67842 = _7211 ^ _67841;
  wire _67843 = uncoded_block[1436] ^ uncoded_block[1458];
  wire _67844 = _67843 ^ _3093;
  wire _67845 = _67842 ^ _67844;
  wire _67846 = _67840 ^ _67845;
  wire _67847 = uncoded_block[1475] ^ uncoded_block[1512];
  wire _67848 = _67847 ^ _30437;
  wire _67849 = uncoded_block[1554] ^ uncoded_block[1609];
  wire _67850 = uncoded_block[1617] ^ uncoded_block[1653];
  wire _67851 = _67849 ^ _67850;
  wire _67852 = _67848 ^ _67851;
  wire _67853 = uncoded_block[1694] ^ uncoded_block[1711];
  wire _67854 = _67853 ^ uncoded_block[1718];
  wire _67855 = _67852 ^ _67854;
  wire _67856 = _67846 ^ _67855;
  wire _67857 = _67834 ^ _67856;
  wire _67858 = uncoded_block[33] ^ uncoded_block[47];
  wire _67859 = uncoded_block[60] ^ uncoded_block[88];
  wire _67860 = _67858 ^ _67859;
  wire _67861 = uncoded_block[135] ^ uncoded_block[146];
  wire _67862 = _67861 ^ _20013;
  wire _67863 = _67860 ^ _67862;
  wire _67864 = _4084 ^ _59702;
  wire _67865 = uncoded_block[352] ^ uncoded_block[370];
  wire _67866 = uncoded_block[404] ^ uncoded_block[446];
  wire _67867 = _67865 ^ _67866;
  wire _67868 = _67864 ^ _67867;
  wire _67869 = _67863 ^ _67868;
  wire _67870 = uncoded_block[452] ^ uncoded_block[471];
  wire _67871 = _67870 ^ _49253;
  wire _67872 = uncoded_block[561] ^ uncoded_block[595];
  wire _67873 = _67872 ^ _2742;
  wire _67874 = _67871 ^ _67873;
  wire _67875 = uncoded_block[675] ^ uncoded_block[684];
  wire _67876 = uncoded_block[757] ^ uncoded_block[765];
  wire _67877 = _67875 ^ _67876;
  wire _67878 = uncoded_block[777] ^ uncoded_block[793];
  wire _67879 = uncoded_block[807] ^ uncoded_block[849];
  wire _67880 = _67878 ^ _67879;
  wire _67881 = _67877 ^ _67880;
  wire _67882 = _67874 ^ _67881;
  wire _67883 = _67869 ^ _67882;
  wire _67884 = uncoded_block[853] ^ uncoded_block[923];
  wire _67885 = uncoded_block[941] ^ uncoded_block[974];
  wire _67886 = _67884 ^ _67885;
  wire _67887 = uncoded_block[985] ^ uncoded_block[1019];
  wire _67888 = uncoded_block[1056] ^ uncoded_block[1072];
  wire _67889 = _67887 ^ _67888;
  wire _67890 = _67886 ^ _67889;
  wire _67891 = uncoded_block[1096] ^ uncoded_block[1131];
  wire _67892 = uncoded_block[1133] ^ uncoded_block[1196];
  wire _67893 = _67891 ^ _67892;
  wire _67894 = uncoded_block[1210] ^ uncoded_block[1274];
  wire _67895 = uncoded_block[1275] ^ uncoded_block[1287];
  wire _67896 = _67894 ^ _67895;
  wire _67897 = _67893 ^ _67896;
  wire _67898 = _67890 ^ _67897;
  wire _67899 = uncoded_block[1296] ^ uncoded_block[1354];
  wire _67900 = uncoded_block[1382] ^ uncoded_block[1403];
  wire _67901 = _67899 ^ _67900;
  wire _67902 = uncoded_block[1438] ^ uncoded_block[1454];
  wire _67903 = _67902 ^ _60900;
  wire _67904 = _67901 ^ _67903;
  wire _67905 = uncoded_block[1546] ^ uncoded_block[1581];
  wire _67906 = uncoded_block[1624] ^ uncoded_block[1644];
  wire _67907 = _67905 ^ _67906;
  wire _67908 = _67907 ^ uncoded_block[1706];
  wire _67909 = _67904 ^ _67908;
  wire _67910 = _67898 ^ _67909;
  wire _67911 = _67883 ^ _67910;
  wire _67912 = uncoded_block[34] ^ uncoded_block[44];
  wire _67913 = uncoded_block[72] ^ uncoded_block[97];
  wire _67914 = _67912 ^ _67913;
  wire _67915 = uncoded_block[131] ^ uncoded_block[143];
  wire _67916 = _67915 ^ _30082;
  wire _67917 = _67914 ^ _67916;
  wire _67918 = uncoded_block[231] ^ uncoded_block[255];
  wire _67919 = uncoded_block[280] ^ uncoded_block[329];
  wire _67920 = _67918 ^ _67919;
  wire _67921 = uncoded_block[348] ^ uncoded_block[390];
  wire _67922 = _67921 ^ _24707;
  wire _67923 = _67920 ^ _67922;
  wire _67924 = _67917 ^ _67923;
  wire _67925 = uncoded_block[494] ^ uncoded_block[504];
  wire _67926 = uncoded_block[510] ^ uncoded_block[516];
  wire _67927 = _67925 ^ _67926;
  wire _67928 = uncoded_block[584] ^ uncoded_block[599];
  wire _67929 = uncoded_block[632] ^ uncoded_block[665];
  wire _67930 = _67928 ^ _67929;
  wire _67931 = _67927 ^ _67930;
  wire _67932 = uncoded_block[671] ^ uncoded_block[690];
  wire _67933 = uncoded_block[760] ^ uncoded_block[768];
  wire _67934 = _67932 ^ _67933;
  wire _67935 = uncoded_block[782] ^ uncoded_block[820];
  wire _67936 = uncoded_block[833] ^ uncoded_block[849];
  wire _67937 = _67935 ^ _67936;
  wire _67938 = _67934 ^ _67937;
  wire _67939 = _67931 ^ _67938;
  wire _67940 = _67924 ^ _67939;
  wire _67941 = uncoded_block[907] ^ uncoded_block[917];
  wire _67942 = uncoded_block[947] ^ uncoded_block[988];
  wire _67943 = _67941 ^ _67942;
  wire _67944 = uncoded_block[1065] ^ uncoded_block[1104];
  wire _67945 = _1356 ^ _67944;
  wire _67946 = _67943 ^ _67945;
  wire _67947 = uncoded_block[1148] ^ uncoded_block[1198];
  wire _67948 = uncoded_block[1238] ^ uncoded_block[1268];
  wire _67949 = _67947 ^ _67948;
  wire _67950 = uncoded_block[1278] ^ uncoded_block[1308];
  wire _67951 = _67950 ^ _2269;
  wire _67952 = _67949 ^ _67951;
  wire _67953 = _67946 ^ _67952;
  wire _67954 = uncoded_block[1361] ^ uncoded_block[1424];
  wire _67955 = uncoded_block[1435] ^ uncoded_block[1510];
  wire _67956 = _67954 ^ _67955;
  wire _67957 = uncoded_block[1515] ^ uncoded_block[1530];
  wire _67958 = uncoded_block[1538] ^ uncoded_block[1560];
  wire _67959 = _67957 ^ _67958;
  wire _67960 = _67956 ^ _67959;
  wire _67961 = uncoded_block[1589] ^ uncoded_block[1607];
  wire _67962 = uncoded_block[1626] ^ uncoded_block[1640];
  wire _67963 = _67961 ^ _67962;
  wire _67964 = _67963 ^ uncoded_block[1667];
  wire _67965 = _67960 ^ _67964;
  wire _67966 = _67953 ^ _67965;
  wire _67967 = _67940 ^ _67966;
  wire _67968 = uncoded_block[14] ^ uncoded_block[35];
  wire _67969 = _46913 ^ _67968;
  wire _67970 = uncoded_block[66] ^ uncoded_block[83];
  wire _67971 = _67970 ^ _64464;
  wire _67972 = _67969 ^ _67971;
  wire _67973 = uncoded_block[153] ^ uncoded_block[164];
  wire _67974 = _33056 ^ _67973;
  wire _67975 = uncoded_block[187] ^ uncoded_block[212];
  wire _67976 = _61781 ^ _67975;
  wire _67977 = _67974 ^ _67976;
  wire _67978 = _67972 ^ _67977;
  wire _67979 = uncoded_block[225] ^ uncoded_block[248];
  wire _67980 = _67979 ^ _4803;
  wire _67981 = _35929 ^ _48476;
  wire _67982 = _67980 ^ _67981;
  wire _67983 = uncoded_block[335] ^ uncoded_block[371];
  wire _67984 = uncoded_block[406] ^ uncoded_block[422];
  wire _67985 = _67983 ^ _67984;
  wire _67986 = _42300 ^ _2660;
  wire _67987 = _67985 ^ _67986;
  wire _67988 = _67982 ^ _67987;
  wire _67989 = _67978 ^ _67988;
  wire _67990 = uncoded_block[488] ^ uncoded_block[504];
  wire _67991 = uncoded_block[527] ^ uncoded_block[536];
  wire _67992 = _67990 ^ _67991;
  wire _67993 = _64508 ^ _67801;
  wire _67994 = _67992 ^ _67993;
  wire _67995 = uncoded_block[591] ^ uncoded_block[612];
  wire _67996 = _67995 ^ _2720;
  wire _67997 = _65691 ^ _64521;
  wire _67998 = _67996 ^ _67997;
  wire _67999 = _67994 ^ _67998;
  wire _68000 = uncoded_block[722] ^ uncoded_block[736];
  wire _68001 = _64523 ^ _68000;
  wire _68002 = uncoded_block[737] ^ uncoded_block[767];
  wire _68003 = _68002 ^ _36469;
  wire _68004 = _68001 ^ _68003;
  wire _68005 = uncoded_block[828] ^ uncoded_block[836];
  wire _68006 = _61859 ^ _68005;
  wire _68007 = uncoded_block[866] ^ uncoded_block[909];
  wire _68008 = _46711 ^ _68007;
  wire _68009 = _68006 ^ _68008;
  wire _68010 = _68004 ^ _68009;
  wire _68011 = _67999 ^ _68010;
  wire _68012 = _67989 ^ _68011;
  wire _68013 = uncoded_block[915] ^ uncoded_block[937];
  wire _68014 = _68013 ^ _1300;
  wire _68015 = _32427 ^ _64557;
  wire _68016 = _68014 ^ _68015;
  wire _68017 = uncoded_block[1046] ^ uncoded_block[1068];
  wire _68018 = uncoded_block[1081] ^ uncoded_block[1088];
  wire _68019 = _68017 ^ _68018;
  wire _68020 = uncoded_block[1107] ^ uncoded_block[1118];
  wire _68021 = uncoded_block[1136] ^ uncoded_block[1152];
  wire _68022 = _68020 ^ _68021;
  wire _68023 = _68019 ^ _68022;
  wire _68024 = _68016 ^ _68023;
  wire _68025 = _63324 ^ _2965;
  wire _68026 = _2982 ^ _62416;
  wire _68027 = _68025 ^ _68026;
  wire _68028 = uncoded_block[1239] ^ uncoded_block[1261];
  wire _68029 = uncoded_block[1268] ^ uncoded_block[1285];
  wire _68030 = _68028 ^ _68029;
  wire _68031 = uncoded_block[1303] ^ uncoded_block[1341];
  wire _68032 = _26274 ^ _68031;
  wire _68033 = _68030 ^ _68032;
  wire _68034 = _68027 ^ _68033;
  wire _68035 = _68024 ^ _68034;
  wire _68036 = uncoded_block[1344] ^ uncoded_block[1373];
  wire _68037 = _68036 ^ _64595;
  wire _68038 = _2318 ^ _64603;
  wire _68039 = _68037 ^ _68038;
  wire _68040 = _64604 ^ _64607;
  wire _68041 = _39834 ^ _63974;
  wire _68042 = _68040 ^ _68041;
  wire _68043 = _68039 ^ _68042;
  wire _68044 = _64613 ^ _14006;
  wire _68045 = uncoded_block[1651] ^ uncoded_block[1698];
  wire _68046 = _68045 ^ uncoded_block[1704];
  wire _68047 = _68044 ^ _68046;
  wire _68048 = _68043 ^ _68047;
  wire _68049 = _68035 ^ _68048;
  wire _68050 = _68012 ^ _68049;
  wire _68051 = uncoded_block[0] ^ uncoded_block[38];
  wire _68052 = uncoded_block[87] ^ uncoded_block[98];
  wire _68053 = _68051 ^ _68052;
  wire _68054 = uncoded_block[151] ^ uncoded_block[166];
  wire _68055 = uncoded_block[189] ^ uncoded_block[219];
  wire _68056 = _68054 ^ _68055;
  wire _68057 = _68053 ^ _68056;
  wire _68058 = uncoded_block[280] ^ uncoded_block[324];
  wire _68059 = _7432 ^ _68058;
  wire _68060 = uncoded_block[333] ^ uncoded_block[357];
  wire _68061 = uncoded_block[404] ^ uncoded_block[429];
  wire _68062 = _68060 ^ _68061;
  wire _68063 = _68059 ^ _68062;
  wire _68064 = _68057 ^ _68063;
  wire _68065 = uncoded_block[462] ^ uncoded_block[497];
  wire _68066 = uncoded_block[553] ^ uncoded_block[559];
  wire _68067 = _68065 ^ _68066;
  wire _68068 = uncoded_block[592] ^ uncoded_block[602];
  wire _68069 = uncoded_block[643] ^ uncoded_block[663];
  wire _68070 = _68068 ^ _68069;
  wire _68071 = _68067 ^ _68070;
  wire _68072 = uncoded_block[729] ^ uncoded_block[741];
  wire _68073 = _38450 ^ _68072;
  wire _68074 = uncoded_block[831] ^ uncoded_block[876];
  wire _68075 = _58182 ^ _68074;
  wire _68076 = _68073 ^ _68075;
  wire _68077 = _68071 ^ _68076;
  wire _68078 = _68064 ^ _68077;
  wire _68079 = uncoded_block[901] ^ uncoded_block[920];
  wire _68080 = uncoded_block[946] ^ uncoded_block[1002];
  wire _68081 = _68079 ^ _68080;
  wire _68082 = uncoded_block[1034] ^ uncoded_block[1051];
  wire _68083 = _68082 ^ _19794;
  wire _68084 = _68081 ^ _68083;
  wire _68085 = uncoded_block[1154] ^ uncoded_block[1199];
  wire _68086 = uncoded_block[1206] ^ uncoded_block[1257];
  wire _68087 = _68085 ^ _68086;
  wire _68088 = uncoded_block[1279] ^ uncoded_block[1301];
  wire _68089 = uncoded_block[1330] ^ uncoded_block[1370];
  wire _68090 = _68088 ^ _68089;
  wire _68091 = _68087 ^ _68090;
  wire _68092 = _68084 ^ _68091;
  wire _68093 = uncoded_block[1377] ^ uncoded_block[1400];
  wire _68094 = uncoded_block[1401] ^ uncoded_block[1431];
  wire _68095 = _68093 ^ _68094;
  wire _68096 = uncoded_block[1490] ^ uncoded_block[1511];
  wire _68097 = uncoded_block[1520] ^ uncoded_block[1529];
  wire _68098 = _68096 ^ _68097;
  wire _68099 = _68095 ^ _68098;
  wire _68100 = uncoded_block[1566] ^ uncoded_block[1583];
  wire _68101 = uncoded_block[1597] ^ uncoded_block[1643];
  wire _68102 = _68100 ^ _68101;
  wire _68103 = _68102 ^ uncoded_block[1658];
  wire _68104 = _68099 ^ _68103;
  wire _68105 = _68092 ^ _68104;
  wire _68106 = _68078 ^ _68105;
  wire _68107 = uncoded_block[43] ^ uncoded_block[55];
  wire _68108 = _1691 ^ _68107;
  wire _68109 = uncoded_block[75] ^ uncoded_block[103];
  wire _68110 = uncoded_block[120] ^ uncoded_block[145];
  wire _68111 = _68109 ^ _68110;
  wire _68112 = _68108 ^ _68111;
  wire _68113 = uncoded_block[161] ^ uncoded_block[195];
  wire _68114 = _68113 ^ _39928;
  wire _68115 = uncoded_block[268] ^ uncoded_block[308];
  wire _68116 = _67789 ^ _68115;
  wire _68117 = _68114 ^ _68116;
  wire _68118 = _68112 ^ _68117;
  wire _68119 = uncoded_block[337] ^ uncoded_block[362];
  wire _68120 = _8058 ^ _68119;
  wire _68121 = uncoded_block[378] ^ uncoded_block[410];
  wire _68122 = uncoded_block[414] ^ uncoded_block[432];
  wire _68123 = _68121 ^ _68122;
  wire _68124 = _68120 ^ _68123;
  wire _68125 = uncoded_block[489] ^ uncoded_block[506];
  wire _68126 = _3416 ^ _68125;
  wire _68127 = uncoded_block[516] ^ uncoded_block[542];
  wire _68128 = uncoded_block[572] ^ uncoded_block[578];
  wire _68129 = _68127 ^ _68128;
  wire _68130 = _68126 ^ _68129;
  wire _68131 = _68124 ^ _68130;
  wire _68132 = _68118 ^ _68131;
  wire _68133 = uncoded_block[613] ^ uncoded_block[644];
  wire _68134 = uncoded_block[646] ^ uncoded_block[653];
  wire _68135 = _68133 ^ _68134;
  wire _68136 = uncoded_block[695] ^ uncoded_block[707];
  wire _68137 = uncoded_block[718] ^ uncoded_block[726];
  wire _68138 = _68136 ^ _68137;
  wire _68139 = _68135 ^ _68138;
  wire _68140 = uncoded_block[763] ^ uncoded_block[776];
  wire _68141 = _68140 ^ _1224;
  wire _68142 = uncoded_block[794] ^ uncoded_block[831];
  wire _68143 = _68142 ^ _54762;
  wire _68144 = _68141 ^ _68143;
  wire _68145 = _68139 ^ _68144;
  wire _68146 = uncoded_block[887] ^ uncoded_block[906];
  wire _68147 = _68146 ^ _32411;
  wire _68148 = uncoded_block[964] ^ uncoded_block[984];
  wire _68149 = uncoded_block[989] ^ uncoded_block[1010];
  wire _68150 = _68148 ^ _68149;
  wire _68151 = _68147 ^ _68150;
  wire _68152 = uncoded_block[1061] ^ uncoded_block[1070];
  wire _68153 = _4417 ^ _68152;
  wire _68154 = uncoded_block[1074] ^ uncoded_block[1115];
  wire _68155 = uncoded_block[1123] ^ uncoded_block[1135];
  wire _68156 = _68154 ^ _68155;
  wire _68157 = _68153 ^ _68156;
  wire _68158 = _68151 ^ _68157;
  wire _68159 = _68145 ^ _68158;
  wire _68160 = _68132 ^ _68159;
  wire _68161 = uncoded_block[1168] ^ uncoded_block[1177];
  wire _68162 = uncoded_block[1191] ^ uncoded_block[1206];
  wire _68163 = _68161 ^ _68162;
  wire _68164 = uncoded_block[1298] ^ uncoded_block[1310];
  wire _68165 = _57498 ^ _68164;
  wire _68166 = _68163 ^ _68165;
  wire _68167 = uncoded_block[1324] ^ uncoded_block[1369];
  wire _68168 = uncoded_block[1385] ^ uncoded_block[1405];
  wire _68169 = _68167 ^ _68168;
  wire _68170 = uncoded_block[1431] ^ uncoded_block[1450];
  wire _68171 = uncoded_block[1461] ^ uncoded_block[1473];
  wire _68172 = _68170 ^ _68171;
  wire _68173 = _68169 ^ _68172;
  wire _68174 = _68166 ^ _68173;
  wire _68175 = uncoded_block[1478] ^ uncoded_block[1487];
  wire _68176 = uncoded_block[1613] ^ uncoded_block[1618];
  wire _68177 = _68175 ^ _68176;
  wire _68178 = uncoded_block[1619] ^ uncoded_block[1658];
  wire _68179 = _68178 ^ _62121;
  wire _68180 = _68177 ^ _68179;
  wire _68181 = uncoded_block[1697] ^ uncoded_block[1712];
  wire _68182 = _68181 ^ uncoded_block[1713];
  wire _68183 = _68180 ^ _68182;
  wire _68184 = _68174 ^ _68183;
  wire _68185 = _68160 ^ _68184;
  wire _68186 = uncoded_block[26] ^ uncoded_block[65];
  wire _68187 = uncoded_block[100] ^ uncoded_block[137];
  wire _68188 = _68186 ^ _68187;
  wire _68189 = uncoded_block[154] ^ uncoded_block[181];
  wire _68190 = uncoded_block[206] ^ uncoded_block[243];
  wire _68191 = _68189 ^ _68190;
  wire _68192 = _68188 ^ _68191;
  wire _68193 = uncoded_block[245] ^ uncoded_block[307];
  wire _68194 = uncoded_block[320] ^ uncoded_block[334];
  wire _68195 = _68193 ^ _68194;
  wire _68196 = uncoded_block[353] ^ uncoded_block[403];
  wire _68197 = uncoded_block[436] ^ uncoded_block[479];
  wire _68198 = _68196 ^ _68197;
  wire _68199 = _68195 ^ _68198;
  wire _68200 = _68192 ^ _68199;
  wire _68201 = uncoded_block[488] ^ uncoded_block[517];
  wire _68202 = uncoded_block[530] ^ uncoded_block[572];
  wire _68203 = _68201 ^ _68202;
  wire _68204 = uncoded_block[608] ^ uncoded_block[662];
  wire _68205 = uncoded_block[665] ^ uncoded_block[700];
  wire _68206 = _68204 ^ _68205;
  wire _68207 = _68203 ^ _68206;
  wire _68208 = uncoded_block[701] ^ uncoded_block[749];
  wire _68209 = uncoded_block[750] ^ uncoded_block[791];
  wire _68210 = _68208 ^ _68209;
  wire _68211 = uncoded_block[803] ^ uncoded_block[870];
  wire _68212 = uncoded_block[881] ^ uncoded_block[887];
  wire _68213 = _68211 ^ _68212;
  wire _68214 = _68210 ^ _68213;
  wire _68215 = _68207 ^ _68214;
  wire _68216 = _68200 ^ _68215;
  wire _68217 = uncoded_block[928] ^ uncoded_block[932];
  wire _68218 = uncoded_block[961] ^ uncoded_block[972];
  wire _68219 = _68217 ^ _68218;
  wire _68220 = uncoded_block[1018] ^ uncoded_block[1044];
  wire _68221 = uncoded_block[1064] ^ uncoded_block[1088];
  wire _68222 = _68220 ^ _68221;
  wire _68223 = _68219 ^ _68222;
  wire _68224 = uncoded_block[1128] ^ uncoded_block[1143];
  wire _68225 = uncoded_block[1164] ^ uncoded_block[1173];
  wire _68226 = _68224 ^ _68225;
  wire _68227 = uncoded_block[1211] ^ uncoded_block[1252];
  wire _68228 = uncoded_block[1264] ^ uncoded_block[1291];
  wire _68229 = _68227 ^ _68228;
  wire _68230 = _68226 ^ _68229;
  wire _68231 = _68223 ^ _68230;
  wire _68232 = uncoded_block[1321] ^ uncoded_block[1374];
  wire _68233 = uncoded_block[1377] ^ uncoded_block[1418];
  wire _68234 = _68232 ^ _68233;
  wire _68235 = uncoded_block[1432] ^ uncoded_block[1551];
  wire _68236 = uncoded_block[1572] ^ uncoded_block[1583];
  wire _68237 = _68235 ^ _68236;
  wire _68238 = _68234 ^ _68237;
  wire _68239 = uncoded_block[1640] ^ uncoded_block[1674];
  wire _68240 = _11849 ^ _68239;
  wire _68241 = _68240 ^ uncoded_block[1684];
  wire _68242 = _68238 ^ _68241;
  wire _68243 = _68231 ^ _68242;
  wire _68244 = _68216 ^ _68243;
  wire _68245 = uncoded_block[129] ^ uncoded_block[140];
  wire _68246 = _68245 ^ _33494;
  wire _68247 = _64632 ^ _68246;
  wire _68248 = uncoded_block[285] ^ uncoded_block[330];
  wire _68249 = _8616 ^ _68248;
  wire _68250 = uncoded_block[335] ^ uncoded_block[385];
  wire _68251 = _68250 ^ _10340;
  wire _68252 = _68249 ^ _68251;
  wire _68253 = _68247 ^ _68252;
  wire _68254 = uncoded_block[462] ^ uncoded_block[477];
  wire _68255 = uncoded_block[520] ^ uncoded_block[547];
  wire _68256 = _68254 ^ _68255;
  wire _68257 = uncoded_block[630] ^ uncoded_block[654];
  wire _68258 = _64677 ^ _68257;
  wire _68259 = _68256 ^ _68258;
  wire _68260 = uncoded_block[671] ^ uncoded_block[706];
  wire _68261 = uncoded_block[731] ^ uncoded_block[756];
  wire _68262 = _68260 ^ _68261;
  wire _68263 = uncoded_block[786] ^ uncoded_block[818];
  wire _68264 = _68263 ^ _67204;
  wire _68265 = _68262 ^ _68264;
  wire _68266 = _68259 ^ _68265;
  wire _68267 = _68253 ^ _68266;
  wire _68268 = uncoded_block[924] ^ uncoded_block[959];
  wire _68269 = uncoded_block[981] ^ uncoded_block[1014];
  wire _68270 = _68268 ^ _68269;
  wire _68271 = uncoded_block[1023] ^ uncoded_block[1070];
  wire _68272 = uncoded_block[1099] ^ uncoded_block[1116];
  wire _68273 = _68271 ^ _68272;
  wire _68274 = _68270 ^ _68273;
  wire _68275 = uncoded_block[1164] ^ uncoded_block[1189];
  wire _68276 = uncoded_block[1190] ^ uncoded_block[1226];
  wire _68277 = _68275 ^ _68276;
  wire _68278 = uncoded_block[1230] ^ uncoded_block[1287];
  wire _68279 = uncoded_block[1292] ^ uncoded_block[1341];
  wire _68280 = _68278 ^ _68279;
  wire _68281 = _68277 ^ _68280;
  wire _68282 = _68274 ^ _68281;
  wire _68283 = uncoded_block[1359] ^ uncoded_block[1401];
  wire _68284 = uncoded_block[1408] ^ uncoded_block[1439];
  wire _68285 = _68283 ^ _68284;
  wire _68286 = uncoded_block[1441] ^ uncoded_block[1459];
  wire _68287 = uncoded_block[1465] ^ uncoded_block[1491];
  wire _68288 = _68286 ^ _68287;
  wire _68289 = _68285 ^ _68288;
  wire _68290 = uncoded_block[1513] ^ uncoded_block[1556];
  wire _68291 = uncoded_block[1620] ^ uncoded_block[1694];
  wire _68292 = _68290 ^ _68291;
  wire _68293 = _68292 ^ uncoded_block[1718];
  wire _68294 = _68289 ^ _68293;
  wire _68295 = _68282 ^ _68294;
  wire _68296 = _68267 ^ _68295;
  wire _68297 = uncoded_block[19] ^ uncoded_block[53];
  wire _68298 = uncoded_block[63] ^ uncoded_block[108];
  wire _68299 = _68297 ^ _68298;
  wire _68300 = uncoded_block[178] ^ uncoded_block[198];
  wire _68301 = _68245 ^ _68300;
  wire _68302 = _68299 ^ _68301;
  wire _68303 = uncoded_block[244] ^ uncoded_block[258];
  wire _68304 = uncoded_block[298] ^ uncoded_block[314];
  wire _68305 = _68303 ^ _68304;
  wire _68306 = uncoded_block[341] ^ uncoded_block[368];
  wire _68307 = uncoded_block[391] ^ uncoded_block[417];
  wire _68308 = _68306 ^ _68307;
  wire _68309 = _68305 ^ _68308;
  wire _68310 = _68302 ^ _68309;
  wire _68311 = uncoded_block[441] ^ uncoded_block[454];
  wire _68312 = uncoded_block[457] ^ uncoded_block[534];
  wire _68313 = _68311 ^ _68312;
  wire _68314 = uncoded_block[555] ^ uncoded_block[579];
  wire _68315 = uncoded_block[593] ^ uncoded_block[634];
  wire _68316 = _68314 ^ _68315;
  wire _68317 = _68313 ^ _68316;
  wire _68318 = uncoded_block[640] ^ uncoded_block[691];
  wire _68319 = uncoded_block[710] ^ uncoded_block[746];
  wire _68320 = _68318 ^ _68319;
  wire _68321 = uncoded_block[762] ^ uncoded_block[795];
  wire _68322 = uncoded_block[807] ^ uncoded_block[858];
  wire _68323 = _68321 ^ _68322;
  wire _68324 = _68320 ^ _68323;
  wire _68325 = _68317 ^ _68324;
  wire _68326 = _68310 ^ _68325;
  wire _68327 = uncoded_block[874] ^ uncoded_block[893];
  wire _68328 = uncoded_block[898] ^ uncoded_block[986];
  wire _68329 = _68327 ^ _68328;
  wire _68330 = uncoded_block[1002] ^ uncoded_block[1018];
  wire _68331 = uncoded_block[1037] ^ uncoded_block[1073];
  wire _68332 = _68330 ^ _68331;
  wire _68333 = _68329 ^ _68332;
  wire _68334 = uncoded_block[1075] ^ uncoded_block[1123];
  wire _68335 = uncoded_block[1157] ^ uncoded_block[1170];
  wire _68336 = _68334 ^ _68335;
  wire _68337 = uncoded_block[1198] ^ uncoded_block[1227];
  wire _68338 = uncoded_block[1244] ^ uncoded_block[1286];
  wire _68339 = _68337 ^ _68338;
  wire _68340 = _68336 ^ _68339;
  wire _68341 = _68333 ^ _68340;
  wire _68342 = uncoded_block[1322] ^ uncoded_block[1345];
  wire _68343 = uncoded_block[1366] ^ uncoded_block[1404];
  wire _68344 = _68342 ^ _68343;
  wire _68345 = uncoded_block[1445] ^ uncoded_block[1493];
  wire _68346 = _68345 ^ _13478;
  wire _68347 = _68344 ^ _68346;
  wire _68348 = uncoded_block[1631] ^ uncoded_block[1706];
  wire _68349 = _63381 ^ _68348;
  wire _68350 = _68349 ^ uncoded_block[1707];
  wire _68351 = _68347 ^ _68350;
  wire _68352 = _68341 ^ _68351;
  wire _68353 = _68326 ^ _68352;
  wire _68354 = uncoded_block[8] ^ uncoded_block[41];
  wire _68355 = uncoded_block[60] ^ uncoded_block[80];
  wire _68356 = _68354 ^ _68355;
  wire _68357 = uncoded_block[82] ^ uncoded_block[117];
  wire _68358 = uncoded_block[139] ^ uncoded_block[170];
  wire _68359 = _68357 ^ _68358;
  wire _68360 = _68356 ^ _68359;
  wire _68361 = uncoded_block[211] ^ uncoded_block[271];
  wire _68362 = _49666 ^ _68361;
  wire _68363 = uncoded_block[281] ^ uncoded_block[293];
  wire _68364 = _10303 ^ _68363;
  wire _68365 = _68362 ^ _68364;
  wire _68366 = _68360 ^ _68365;
  wire _68367 = uncoded_block[325] ^ uncoded_block[334];
  wire _68368 = _68367 ^ _4131;
  wire _68369 = uncoded_block[394] ^ uncoded_block[435];
  wire _68370 = uncoded_block[445] ^ uncoded_block[467];
  wire _68371 = _68369 ^ _68370;
  wire _68372 = _68368 ^ _68371;
  wire _68373 = uncoded_block[487] ^ uncoded_block[503];
  wire _68374 = uncoded_block[519] ^ uncoded_block[535];
  wire _68375 = _68373 ^ _68374;
  wire _68376 = uncoded_block[555] ^ uncoded_block[590];
  wire _68377 = uncoded_block[614] ^ uncoded_block[638];
  wire _68378 = _68376 ^ _68377;
  wire _68379 = _68375 ^ _68378;
  wire _68380 = _68372 ^ _68379;
  wire _68381 = _68366 ^ _68380;
  wire _68382 = uncoded_block[648] ^ uncoded_block[660];
  wire _68383 = uncoded_block[681] ^ uncoded_block[709];
  wire _68384 = _68382 ^ _68383;
  wire _68385 = uncoded_block[720] ^ uncoded_block[735];
  wire _68386 = uncoded_block[739] ^ uncoded_block[758];
  wire _68387 = _68385 ^ _68386;
  wire _68388 = _68384 ^ _68387;
  wire _68389 = uncoded_block[779] ^ uncoded_block[806];
  wire _68390 = uncoded_block[815] ^ uncoded_block[846];
  wire _68391 = _68389 ^ _68390;
  wire _68392 = uncoded_block[860] ^ uncoded_block[871];
  wire _68393 = uncoded_block[890] ^ uncoded_block[902];
  wire _68394 = _68392 ^ _68393;
  wire _68395 = _68391 ^ _68394;
  wire _68396 = _68388 ^ _68395;
  wire _68397 = uncoded_block[908] ^ uncoded_block[971];
  wire _68398 = uncoded_block[976] ^ uncoded_block[992];
  wire _68399 = _68397 ^ _68398;
  wire _68400 = uncoded_block[1010] ^ uncoded_block[1079];
  wire _68401 = _68400 ^ _16880;
  wire _68402 = _68399 ^ _68401;
  wire _68403 = uncoded_block[1135] ^ uncoded_block[1154];
  wire _68404 = _68403 ^ _3734;
  wire _68405 = uncoded_block[1172] ^ uncoded_block[1182];
  wire _68406 = uncoded_block[1237] ^ uncoded_block[1260];
  wire _68407 = _68405 ^ _68406;
  wire _68408 = _68404 ^ _68407;
  wire _68409 = _68402 ^ _68408;
  wire _68410 = _68396 ^ _68409;
  wire _68411 = _68381 ^ _68410;
  wire _68412 = uncoded_block[1261] ^ uncoded_block[1276];
  wire _68413 = _68412 ^ _66960;
  wire _68414 = uncoded_block[1293] ^ uncoded_block[1323];
  wire _68415 = _68414 ^ _64285;
  wire _68416 = _68413 ^ _68415;
  wire _68417 = uncoded_block[1381] ^ uncoded_block[1395];
  wire _68418 = uncoded_block[1438] ^ uncoded_block[1467];
  wire _68419 = _68417 ^ _68418;
  wire _68420 = uncoded_block[1495] ^ uncoded_block[1504];
  wire _68421 = _68420 ^ _64305;
  wire _68422 = _68419 ^ _68421;
  wire _68423 = _68416 ^ _68422;
  wire _68424 = uncoded_block[1533] ^ uncoded_block[1544];
  wire _68425 = uncoded_block[1549] ^ uncoded_block[1580];
  wire _68426 = _68424 ^ _68425;
  wire _68427 = uncoded_block[1586] ^ uncoded_block[1606];
  wire _68428 = uncoded_block[1611] ^ uncoded_block[1627];
  wire _68429 = _68427 ^ _68428;
  wire _68430 = _68426 ^ _68429;
  wire _68431 = uncoded_block[1635] ^ uncoded_block[1708];
  wire _68432 = _68431 ^ uncoded_block[1720];
  wire _68433 = _68430 ^ _68432;
  wire _68434 = _68423 ^ _68433;
  wire _68435 = _68411 ^ _68434;
  wire _68436 = _5423 ^ _53574;
  wire _68437 = _36287 ^ _68436;
  wire _68438 = _3220 ^ _13539;
  wire _68439 = _874 ^ _3225;
  wire _68440 = _68438 ^ _68439;
  wire _68441 = _68437 ^ _68440;
  wire _68442 = _3227 ^ _14047;
  wire _68443 = _68442 ^ _12426;
  wire _68444 = _17568 ^ _25;
  wire _68445 = _13552 ^ _1705;
  wire _68446 = _68444 ^ _68445;
  wire _68447 = _68443 ^ _68446;
  wire _68448 = _68441 ^ _68447;
  wire _68449 = _25510 ^ _63173;
  wire _68450 = _901 ^ _4735;
  wire _68451 = _13558 ^ _33894;
  wire _68452 = _68450 ^ _68451;
  wire _68453 = _68449 ^ _68452;
  wire _68454 = _46543 ^ _29608;
  wire _68455 = _5453 ^ _6763;
  wire _68456 = _23711 ^ _68455;
  wire _68457 = _68454 ^ _68456;
  wire _68458 = _68453 ^ _68457;
  wire _68459 = _68448 ^ _68458;
  wire _68460 = _2498 ^ _10821;
  wire _68461 = _32226 ^ _68460;
  wire _68462 = _10822 ^ _4754;
  wire _68463 = _46554 ^ _1736;
  wire _68464 = _68462 ^ _68463;
  wire _68465 = _68461 ^ _68464;
  wire _68466 = _7999 ^ _11383;
  wire _68467 = _3269 ^ _3271;
  wire _68468 = _68466 ^ _68467;
  wire _68469 = _13577 ^ _41854;
  wire _68470 = _68468 ^ _68469;
  wire _68471 = _68465 ^ _68470;
  wire _68472 = _14092 ^ _13583;
  wire _68473 = _30521 ^ _68472;
  wire _68474 = _26424 ^ _3285;
  wire _68475 = _68473 ^ _68474;
  wire _68476 = _4068 ^ _3289;
  wire _68477 = _6806 ^ _12483;
  wire _68478 = _68476 ^ _68477;
  wire _68479 = _3296 ^ _960;
  wire _68480 = _102 ^ _104;
  wire _68481 = _68479 ^ _68480;
  wire _68482 = _68478 ^ _68481;
  wire _68483 = _68475 ^ _68482;
  wire _68484 = _68471 ^ _68483;
  wire _68485 = _68459 ^ _68484;
  wire _68486 = _2545 ^ _4080;
  wire _68487 = _4081 ^ _35141;
  wire _68488 = _68486 ^ _68487;
  wire _68489 = _8616 ^ _2556;
  wire _68490 = _21466 ^ _68489;
  wire _68491 = _68488 ^ _68490;
  wire _68492 = _2557 ^ _1786;
  wire _68493 = _68492 ^ _978;
  wire _68494 = _984 ^ _3320;
  wire _68495 = _68494 ^ _11965;
  wire _68496 = _68493 ^ _68495;
  wire _68497 = _68491 ^ _68496;
  wire _68498 = _134 ^ _992;
  wire _68499 = _56685 ^ _68498;
  wire _68500 = _2577 ^ _31847;
  wire _68501 = _43685 ^ _68500;
  wire _68502 = _68499 ^ _68501;
  wire _68503 = _16648 ^ _6850;
  wire _68504 = _68503 ^ _30560;
  wire _68505 = _60196 ^ _15173;
  wire _68506 = _68505 ^ _13631;
  wire _68507 = _68504 ^ _68506;
  wire _68508 = _68502 ^ _68507;
  wire _68509 = _68497 ^ _68508;
  wire _68510 = _4132 ^ _2601;
  wire _68511 = _27734 ^ _68510;
  wire _68512 = _60205 ^ _22885;
  wire _68513 = _68511 ^ _68512;
  wire _68514 = _4140 ^ _8079;
  wire _68515 = _4854 ^ _2612;
  wire _68516 = _68514 ^ _68515;
  wire _68517 = uncoded_block[389] ^ uncoded_block[394];
  wire _68518 = _4149 ^ _68517;
  wire _68519 = _68518 ^ _30137;
  wire _68520 = _68516 ^ _68519;
  wire _68521 = _68513 ^ _68520;
  wire _68522 = _184 ^ _8091;
  wire _68523 = _2630 ^ _13112;
  wire _68524 = _68522 ^ _68523;
  wire _68525 = _2633 ^ _9816;
  wire _68526 = _14161 ^ _68525;
  wire _68527 = _68524 ^ _68526;
  wire _68528 = _1857 ^ _27350;
  wire _68529 = _34378 ^ _25607;
  wire _68530 = _68528 ^ _68529;
  wire _68531 = _4185 ^ _3416;
  wire _68532 = _55913 ^ _68531;
  wire _68533 = _68530 ^ _68532;
  wire _68534 = _68527 ^ _68533;
  wire _68535 = _68521 ^ _68534;
  wire _68536 = _68509 ^ _68535;
  wire _68537 = _68485 ^ _68536;
  wire _68538 = _21527 ^ _32308;
  wire _68539 = _13135 ^ _17198;
  wire _68540 = _4905 ^ _30604;
  wire _68541 = _68539 ^ _68540;
  wire _68542 = _68538 ^ _68541;
  wire _68543 = _5611 ^ _38397;
  wire _68544 = _23370 ^ _10947;
  wire _68545 = _68543 ^ _68544;
  wire _68546 = _16709 ^ _4922;
  wire _68547 = _68546 ^ _58455;
  wire _68548 = _68545 ^ _68547;
  wire _68549 = _68542 ^ _68548;
  wire _68550 = _3451 ^ _32324;
  wire _68551 = _23382 ^ _41932;
  wire _68552 = _68550 ^ _68551;
  wire _68553 = _3464 ^ _20110;
  wire _68554 = _6309 ^ _17221;
  wire _68555 = _68553 ^ _68554;
  wire _68556 = _68552 ^ _68555;
  wire _68557 = _28136 ^ _265;
  wire _68558 = _2696 ^ _19656;
  wire _68559 = _68557 ^ _68558;
  wire _68560 = _1938 ^ _17721;
  wire _68561 = _5646 ^ _8152;
  wire _68562 = _68560 ^ _68561;
  wire _68563 = _68559 ^ _68562;
  wire _68564 = _68556 ^ _68563;
  wire _68565 = _68549 ^ _68564;
  wire _68566 = _16734 ^ _13713;
  wire _68567 = _68566 ^ _60258;
  wire _68568 = _17238 ^ _43761;
  wire _68569 = _68568 ^ _46666;
  wire _68570 = _68567 ^ _68569;
  wire _68571 = _304 ^ _64518;
  wire _68572 = _16248 ^ _68571;
  wire _68573 = _7582 ^ _17742;
  wire _68574 = _68573 ^ _16254;
  wire _68575 = _68572 ^ _68574;
  wire _68576 = _68570 ^ _68575;
  wire _68577 = _33622 ^ _43008;
  wire _68578 = _13735 ^ _6985;
  wire _68579 = _8186 ^ _11562;
  wire _68580 = _68578 ^ _68579;
  wire _68581 = _68577 ^ _68580;
  wire _68582 = _14250 ^ _60273;
  wire _68583 = _68582 ^ _55603;
  wire _68584 = uncoded_block[732] ^ uncoded_block[739];
  wire _68585 = _4283 ^ _68584;
  wire _68586 = _342 ^ _68585;
  wire _68587 = _68583 ^ _68586;
  wire _68588 = _68581 ^ _68587;
  wire _68589 = _68576 ^ _68588;
  wire _68590 = _68565 ^ _68589;
  wire _68591 = _352 ^ _5702;
  wire _68592 = _68591 ^ _44571;
  wire _68593 = _5016 ^ _2778;
  wire _68594 = _68593 ^ _60288;
  wire _68595 = _68592 ^ _68594;
  wire _68596 = _3562 ^ _9382;
  wire _68597 = _15800 ^ _68596;
  wire _68598 = _2794 ^ _16786;
  wire _68599 = _68598 ^ _15806;
  wire _68600 = _68597 ^ _68599;
  wire _68601 = _68595 ^ _68600;
  wire _68602 = _36054 ^ _41215;
  wire _68603 = _2026 ^ _2808;
  wire _68604 = _55274 ^ _2812;
  wire _68605 = _68603 ^ _68604;
  wire _68606 = _68602 ^ _68605;
  wire _68607 = _400 ^ _1250;
  wire _68608 = _1253 ^ _47836;
  wire _68609 = _68607 ^ _68608;
  wire _68610 = uncoded_block[852] ^ uncoded_block[855];
  wire _68611 = _68610 ^ _14300;
  wire _68612 = _43048 ^ _68611;
  wire _68613 = _68609 ^ _68612;
  wire _68614 = _68606 ^ _68613;
  wire _68615 = _68601 ^ _68614;
  wire _68616 = _6410 ^ _14302;
  wire _68617 = _5071 ^ _12696;
  wire _68618 = _68616 ^ _68617;
  wire _68619 = _2831 ^ _5079;
  wire _68620 = _68619 ^ _48967;
  wire _68621 = _68618 ^ _68620;
  wire _68622 = _15343 ^ _3617;
  wire _68623 = _68622 ^ _25728;
  wire _68624 = uncoded_block[913] ^ uncoded_block[920];
  wire _68625 = _19252 ^ _68624;
  wire _68626 = _2076 ^ _448;
  wire _68627 = _68625 ^ _68626;
  wire _68628 = _68623 ^ _68627;
  wire _68629 = _68621 ^ _68628;
  wire _68630 = _4377 ^ _13266;
  wire _68631 = _38109 ^ _68630;
  wire _68632 = _7083 ^ _45753;
  wire _68633 = _68632 ^ _22568;
  wire _68634 = _68631 ^ _68633;
  wire _68635 = uncoded_block[973] ^ uncoded_block[978];
  wire _68636 = _467 ^ _68635;
  wire _68637 = _68636 ^ _50209;
  wire _68638 = _68637 ^ _58552;
  wire _68639 = _68634 ^ _68638;
  wire _68640 = _68629 ^ _68639;
  wire _68641 = _68615 ^ _68640;
  wire _68642 = _68590 ^ _68641;
  wire _68643 = _68537 ^ _68642;
  wire _68644 = _28241 ^ _2111;
  wire _68645 = _43085 ^ _13283;
  wire _68646 = _68644 ^ _68645;
  wire _68647 = _1334 ^ _19766;
  wire _68648 = _26211 ^ _68647;
  wire _68649 = _68646 ^ _68648;
  wire _68650 = _11668 ^ _502;
  wire _68651 = _10007 ^ _68650;
  wire _68652 = _512 ^ _2913;
  wire _68653 = _68652 ^ _60342;
  wire _68654 = _68651 ^ _68653;
  wire _68655 = _68649 ^ _68654;
  wire _68656 = _42044 ^ _25773;
  wire _68657 = _5158 ^ _8895;
  wire _68658 = _68656 ^ _68657;
  wire _68659 = _46374 ^ _20253;
  wire _68660 = _68659 ^ _19789;
  wire _68661 = _68658 ^ _68660;
  wire _68662 = _10026 ^ _5169;
  wire _68663 = _68662 ^ _58577;
  wire _68664 = _2165 ^ _7133;
  wire _68665 = _19313 ^ _9489;
  wire _68666 = _68664 ^ _68665;
  wire _68667 = _68663 ^ _68666;
  wire _68668 = _68661 ^ _68667;
  wire _68669 = _68655 ^ _68668;
  wire _68670 = _14886 ^ _58584;
  wire _68671 = _4462 ^ _7141;
  wire _68672 = _6505 ^ _577;
  wire _68673 = _68671 ^ _68672;
  wire _68674 = _68670 ^ _68673;
  wire _68675 = _27105 ^ _40539;
  wire _68676 = _2967 ^ _34961;
  wire _68677 = _68675 ^ _68676;
  wire _68678 = _31213 ^ _53831;
  wire _68679 = _68677 ^ _68678;
  wire _68680 = _68674 ^ _68679;
  wire _68681 = _15431 ^ _6529;
  wire _68682 = _60374 ^ _68681;
  wire _68683 = _2979 ^ _1428;
  wire _68684 = _68683 ^ _23106;
  wire _68685 = _68682 ^ _68684;
  wire _68686 = _4502 ^ _1436;
  wire _68687 = _18400 ^ _31228;
  wire _68688 = _68686 ^ _68687;
  wire _68689 = _13360 ^ _2230;
  wire _68690 = uncoded_block[1246] ^ uncoded_block[1249];
  wire _68691 = _68690 ^ _2235;
  wire _68692 = _68689 ^ _68691;
  wire _68693 = _68688 ^ _68692;
  wire _68694 = _68685 ^ _68693;
  wire _68695 = _68680 ^ _68694;
  wire _68696 = _68669 ^ _68695;
  wire _68697 = _5234 ^ _30361;
  wire _68698 = _68697 ^ _9534;
  wire _68699 = _49897 ^ _2247;
  wire _68700 = _68699 ^ _7794;
  wire _68701 = _68698 ^ _68700;
  wire _68702 = _4529 ^ _30797;
  wire _68703 = _17427 ^ _68702;
  wire _68704 = uncoded_block[1299] ^ uncoded_block[1304];
  wire _68705 = _19369 ^ _68704;
  wire _68706 = _1479 ^ _6572;
  wire _68707 = _68705 ^ _68706;
  wire _68708 = _68703 ^ _68707;
  wire _68709 = _68701 ^ _68708;
  wire _68710 = _8407 ^ _12287;
  wire _68711 = uncoded_block[1326] ^ uncoded_block[1333];
  wire _68712 = _37813 ^ _68711;
  wire _68713 = _68710 ^ _68712;
  wire _68714 = _1495 ^ _9564;
  wire _68715 = _11218 ^ _33363;
  wire _68716 = _68714 ^ _68715;
  wire _68717 = _68713 ^ _68716;
  wire _68718 = _12300 ^ _66058;
  wire _68719 = _8420 ^ _68718;
  wire _68720 = _3834 ^ _12311;
  wire _68721 = _5286 ^ _68720;
  wire _68722 = _68719 ^ _68721;
  wire _68723 = _68717 ^ _68722;
  wire _68724 = _68709 ^ _68723;
  wire _68725 = _691 ^ _28340;
  wire _68726 = _4572 ^ _63711;
  wire _68727 = _68725 ^ _68726;
  wire _68728 = _5962 ^ _8438;
  wire _68729 = _25408 ^ _68728;
  wire _68730 = _68727 ^ _68729;
  wire _68731 = _10683 ^ _1530;
  wire _68732 = _17961 ^ _68731;
  wire _68733 = _1534 ^ _29508;
  wire _68734 = uncoded_block[1443] ^ uncoded_block[1449];
  wire _68735 = _5304 ^ _68734;
  wire _68736 = _68733 ^ _68735;
  wire _68737 = _68732 ^ _68736;
  wire _68738 = _68730 ^ _68737;
  wire _68739 = _18465 ^ _11249;
  wire _68740 = _68739 ^ _9039;
  wire _68741 = _68740 ^ _60431;
  wire _68742 = _1571 ^ _39041;
  wire _68743 = _3115 ^ _7265;
  wire _68744 = _68742 ^ _68743;
  wire _68745 = uncoded_block[1519] ^ uncoded_block[1527];
  wire _68746 = _68745 ^ _9631;
  wire _68747 = _12914 ^ _6006;
  wire _68748 = _68746 ^ _68747;
  wire _68749 = _68744 ^ _68748;
  wire _68750 = _68741 ^ _68749;
  wire _68751 = _68738 ^ _68750;
  wire _68752 = _68724 ^ _68751;
  wire _68753 = _68696 ^ _68752;
  wire _68754 = uncoded_block[1541] ^ uncoded_block[1551];
  wire _68755 = _68754 ^ _6657;
  wire _68756 = _68755 ^ _60440;
  wire _68757 = _774 ^ _20392;
  wire _68758 = _9072 ^ _17007;
  wire _68759 = _68757 ^ _68758;
  wire _68760 = _68756 ^ _68759;
  wire _68761 = _3924 ^ _15538;
  wire _68762 = _6664 ^ _68761;
  wire _68763 = _6673 ^ _1620;
  wire _68764 = _1621 ^ _10742;
  wire _68765 = _68763 ^ _68764;
  wire _68766 = _68762 ^ _68765;
  wire _68767 = _68760 ^ _68766;
  wire _68768 = uncoded_block[1611] ^ uncoded_block[1620];
  wire _68769 = _3154 ^ _68768;
  wire _68770 = _27649 ^ _2404;
  wire _68771 = _68769 ^ _68770;
  wire _68772 = _42177 ^ _3948;
  wire _68773 = _2408 ^ _816;
  wire _68774 = _68772 ^ _68773;
  wire _68775 = _68771 ^ _68774;
  wire _68776 = _4674 ^ _10194;
  wire _68777 = _68776 ^ _27979;
  wire _68778 = _60462 ^ _27223;
  wire _68779 = _68777 ^ _68778;
  wire _68780 = _68775 ^ _68779;
  wire _68781 = _68767 ^ _68780;
  wire _68782 = _832 ^ _20427;
  wire _68783 = _4691 ^ _836;
  wire _68784 = _68782 ^ _68783;
  wire _68785 = uncoded_block[1688] ^ uncoded_block[1693];
  wire _68786 = _68785 ^ _840;
  wire _68787 = _10212 ^ _22773;
  wire _68788 = _68786 ^ _68787;
  wire _68789 = _68784 ^ _68788;
  wire _68790 = _2437 ^ _55813;
  wire _68791 = _1677 ^ uncoded_block[1722];
  wire _68792 = _68790 ^ _68791;
  wire _68793 = _68789 ^ _68792;
  wire _68794 = _68781 ^ _68793;
  wire _68795 = _68753 ^ _68794;
  wire _68796 = _68643 ^ _68795;
  wire _68797 = uncoded_block[5] ^ uncoded_block[15];
  wire _68798 = uncoded_block[57] ^ uncoded_block[87];
  wire _68799 = _68797 ^ _68798;
  wire _68800 = uncoded_block[88] ^ uncoded_block[111];
  wire _68801 = uncoded_block[149] ^ uncoded_block[163];
  wire _68802 = _68800 ^ _68801;
  wire _68803 = _68799 ^ _68802;
  wire _68804 = uncoded_block[191] ^ uncoded_block[198];
  wire _68805 = uncoded_block[216] ^ uncoded_block[237];
  wire _68806 = _68804 ^ _68805;
  wire _68807 = uncoded_block[309] ^ uncoded_block[323];
  wire _68808 = _37959 ^ _68807;
  wire _68809 = _68806 ^ _68808;
  wire _68810 = _68803 ^ _68809;
  wire _68811 = uncoded_block[329] ^ uncoded_block[371];
  wire _68812 = _68811 ^ _18632;
  wire _68813 = uncoded_block[439] ^ uncoded_block[461];
  wire _68814 = _17678 ^ _68813;
  wire _68815 = _68812 ^ _68814;
  wire _68816 = uncoded_block[471] ^ uncoded_block[497];
  wire _68817 = uncoded_block[537] ^ uncoded_block[547];
  wire _68818 = _68816 ^ _68817;
  wire _68819 = uncoded_block[553] ^ uncoded_block[567];
  wire _68820 = uncoded_block[574] ^ uncoded_block[603];
  wire _68821 = _68819 ^ _68820;
  wire _68822 = _68818 ^ _68821;
  wire _68823 = _68815 ^ _68822;
  wire _68824 = _68810 ^ _68823;
  wire _68825 = uncoded_block[667] ^ uncoded_block[682];
  wire _68826 = _12075 ^ _68825;
  wire _68827 = uncoded_block[728] ^ uncoded_block[743];
  wire _68828 = _2762 ^ _68827;
  wire _68829 = _68826 ^ _68828;
  wire _68830 = uncoded_block[764] ^ uncoded_block[781];
  wire _68831 = uncoded_block[811] ^ uncoded_block[819];
  wire _68832 = _68830 ^ _68831;
  wire _68833 = uncoded_block[842] ^ uncoded_block[851];
  wire _68834 = uncoded_block[874] ^ uncoded_block[892];
  wire _68835 = _68833 ^ _68834;
  wire _68836 = _68832 ^ _68835;
  wire _68837 = _68829 ^ _68836;
  wire _68838 = _5083 ^ _6441;
  wire _68839 = uncoded_block[998] ^ uncoded_block[1018];
  wire _68840 = uncoded_block[1033] ^ uncoded_block[1045];
  wire _68841 = _68839 ^ _68840;
  wire _68842 = _68838 ^ _68841;
  wire _68843 = uncoded_block[1099] ^ uncoded_block[1124];
  wire _68844 = _11689 ^ _68843;
  wire _68845 = uncoded_block[1161] ^ uncoded_block[1178];
  wire _68846 = uncoded_block[1180] ^ uncoded_block[1243];
  wire _68847 = _68845 ^ _68846;
  wire _68848 = _68844 ^ _68847;
  wire _68849 = _68842 ^ _68848;
  wire _68850 = _68837 ^ _68849;
  wire _68851 = _68824 ^ _68850;
  wire _68852 = uncoded_block[1260] ^ uncoded_block[1271];
  wire _68853 = uncoded_block[1280] ^ uncoded_block[1307];
  wire _68854 = _68852 ^ _68853;
  wire _68855 = uncoded_block[1331] ^ uncoded_block[1354];
  wire _68856 = _63934 ^ _68855;
  wire _68857 = _68854 ^ _68856;
  wire _68858 = uncoded_block[1396] ^ uncoded_block[1410];
  wire _68859 = _25849 ^ _68858;
  wire _68860 = uncoded_block[1422] ^ uncoded_block[1429];
  wire _68861 = uncoded_block[1486] ^ uncoded_block[1517];
  wire _68862 = _68860 ^ _68861;
  wire _68863 = _68859 ^ _68862;
  wire _68864 = _68857 ^ _68863;
  wire _68865 = uncoded_block[1570] ^ uncoded_block[1588];
  wire _68866 = _63966 ^ _68865;
  wire _68867 = uncoded_block[1602] ^ uncoded_block[1611];
  wire _68868 = uncoded_block[1619] ^ uncoded_block[1628];
  wire _68869 = _68867 ^ _68868;
  wire _68870 = _68866 ^ _68869;
  wire _68871 = uncoded_block[1657] ^ uncoded_block[1708];
  wire _68872 = _68871 ^ uncoded_block[1720];
  wire _68873 = _68870 ^ _68872;
  wire _68874 = _68864 ^ _68873;
  wire _68875 = _68851 ^ _68874;
  wire _68876 = uncoded_block[6] ^ uncoded_block[12];
  wire _68877 = uncoded_block[22] ^ uncoded_block[44];
  wire _68878 = _68876 ^ _68877;
  wire _68879 = uncoded_block[54] ^ uncoded_block[75];
  wire _68880 = uncoded_block[86] ^ uncoded_block[108];
  wire _68881 = _68879 ^ _68880;
  wire _68882 = _68878 ^ _68881;
  wire _68883 = uncoded_block[132] ^ uncoded_block[143];
  wire _68884 = _68883 ^ _21906;
  wire _68885 = uncoded_block[189] ^ uncoded_block[202];
  wire _68886 = _68885 ^ _48830;
  wire _68887 = _68884 ^ _68886;
  wire _68888 = _68882 ^ _68887;
  wire _68889 = uncoded_block[228] ^ uncoded_block[234];
  wire _68890 = _68889 ^ _19061;
  wire _68891 = uncoded_block[300] ^ uncoded_block[308];
  wire _68892 = uncoded_block[314] ^ uncoded_block[327];
  wire _68893 = _68891 ^ _68892;
  wire _68894 = _68890 ^ _68893;
  wire _68895 = uncoded_block[350] ^ uncoded_block[378];
  wire _68896 = _10323 ^ _68895;
  wire _68897 = uncoded_block[391] ^ uncoded_block[401];
  wire _68898 = uncoded_block[410] ^ uncoded_block[428];
  wire _68899 = _68897 ^ _68898;
  wire _68900 = _68896 ^ _68899;
  wire _68901 = _68894 ^ _68900;
  wire _68902 = _68888 ^ _68901;
  wire _68903 = uncoded_block[429] ^ uncoded_block[494];
  wire _68904 = uncoded_block[509] ^ uncoded_block[534];
  wire _68905 = _68903 ^ _68904;
  wire _68906 = uncoded_block[542] ^ uncoded_block[550];
  wire _68907 = _68906 ^ _15239;
  wire _68908 = _68905 ^ _68907;
  wire _68909 = uncoded_block[578] ^ uncoded_block[592];
  wire _68910 = uncoded_block[622] ^ uncoded_block[633];
  wire _68911 = _68909 ^ _68910;
  wire _68912 = uncoded_block[644] ^ uncoded_block[663];
  wire _68913 = uncoded_block[671] ^ uncoded_block[681];
  wire _68914 = _68912 ^ _68913;
  wire _68915 = _68911 ^ _68914;
  wire _68916 = _68908 ^ _68915;
  wire _68917 = uncoded_block[695] ^ uncoded_block[709];
  wire _68918 = _68917 ^ _34442;
  wire _68919 = uncoded_block[754] ^ uncoded_block[763];
  wire _68920 = _68919 ^ _38078;
  wire _68921 = _68918 ^ _68920;
  wire _68922 = _60831 ^ _11609;
  wire _68923 = uncoded_block[890] ^ uncoded_block[916];
  wire _68924 = _64074 ^ _68923;
  wire _68925 = _68922 ^ _68924;
  wire _68926 = _68921 ^ _68925;
  wire _68927 = _68916 ^ _68926;
  wire _68928 = _68902 ^ _68927;
  wire _68929 = uncoded_block[951] ^ uncoded_block[964];
  wire _68930 = _38500 ^ _68929;
  wire _68931 = uncoded_block[982] ^ uncoded_block[1010];
  wire _68932 = _68931 ^ _6462;
  wire _68933 = _68930 ^ _68932;
  wire _68934 = uncoded_block[1042] ^ uncoded_block[1061];
  wire _68935 = _68934 ^ _23969;
  wire _68936 = uncoded_block[1093] ^ uncoded_block[1130];
  wire _68937 = _68936 ^ _5856;
  wire _68938 = _68935 ^ _68937;
  wire _68939 = _68933 ^ _68938;
  wire _68940 = uncoded_block[1158] ^ uncoded_block[1168];
  wire _68941 = _68940 ^ _24910;
  wire _68942 = uncoded_block[1206] ^ uncoded_block[1241];
  wire _68943 = uncoded_block[1243] ^ uncoded_block[1263];
  wire _68944 = _68942 ^ _68943;
  wire _68945 = _68941 ^ _68944;
  wire _68946 = _67313 ^ _3025;
  wire _68947 = uncoded_block[1351] ^ uncoded_block[1379];
  wire _68948 = _26729 ^ _68947;
  wire _68949 = _68946 ^ _68948;
  wire _68950 = _68945 ^ _68949;
  wire _68951 = _68939 ^ _68950;
  wire _68952 = uncoded_block[1393] ^ uncoded_block[1405];
  wire _68953 = uncoded_block[1407] ^ uncoded_block[1435];
  wire _68954 = _68952 ^ _68953;
  wire _68955 = uncoded_block[1440] ^ uncoded_block[1473];
  wire _68956 = uncoded_block[1487] ^ uncoded_block[1503];
  wire _68957 = _68955 ^ _68956;
  wire _68958 = _68954 ^ _68957;
  wire _68959 = uncoded_block[1516] ^ uncoded_block[1543];
  wire _68960 = uncoded_block[1553] ^ uncoded_block[1567];
  wire _68961 = _68959 ^ _68960;
  wire _68962 = uncoded_block[1579] ^ uncoded_block[1610];
  wire _68963 = _68962 ^ _1633;
  wire _68964 = _68961 ^ _68963;
  wire _68965 = _68958 ^ _68964;
  wire _68966 = uncoded_block[1642] ^ uncoded_block[1655];
  wire _68967 = uncoded_block[1658] ^ uncoded_block[1675];
  wire _68968 = _68966 ^ _68967;
  wire _68969 = uncoded_block[1677] ^ uncoded_block[1713];
  wire _68970 = _68969 ^ uncoded_block[1715];
  wire _68971 = _68968 ^ _68970;
  wire _68972 = _68965 ^ _68971;
  wire _68973 = _68951 ^ _68972;
  wire _68974 = _68928 ^ _68973;
  wire _68975 = uncoded_block[90] ^ uncoded_block[104];
  wire _68976 = _9135 ^ _68975;
  wire _68977 = uncoded_block[138] ^ uncoded_block[155];
  wire _68978 = uncoded_block[177] ^ uncoded_block[221];
  wire _68979 = _68977 ^ _68978;
  wire _68980 = _68976 ^ _68979;
  wire _68981 = uncoded_block[252] ^ uncoded_block[271];
  wire _68982 = uncoded_block[287] ^ uncoded_block[310];
  wire _68983 = _68981 ^ _68982;
  wire _68984 = uncoded_block[357] ^ uncoded_block[390];
  wire _68985 = uncoded_block[405] ^ uncoded_block[410];
  wire _68986 = _68984 ^ _68985;
  wire _68987 = _68983 ^ _68986;
  wire _68988 = _68980 ^ _68987;
  wire _68989 = uncoded_block[451] ^ uncoded_block[475];
  wire _68990 = _68989 ^ _26081;
  wire _68991 = uncoded_block[567] ^ uncoded_block[608];
  wire _68992 = uncoded_block[653] ^ uncoded_block[665];
  wire _68993 = _68991 ^ _68992;
  wire _68994 = _68990 ^ _68993;
  wire _68995 = uncoded_block[687] ^ uncoded_block[698];
  wire _68996 = uncoded_block[742] ^ uncoded_block[747];
  wire _68997 = _68995 ^ _68996;
  wire _68998 = uncoded_block[810] ^ uncoded_block[818];
  wire _68999 = uncoded_block[851] ^ uncoded_block[868];
  wire _69000 = _68998 ^ _68999;
  wire _69001 = _68997 ^ _69000;
  wire _69002 = _68994 ^ _69001;
  wire _69003 = _68988 ^ _69002;
  wire _69004 = uncoded_block[911] ^ uncoded_block[927];
  wire _69005 = uncoded_block[984] ^ uncoded_block[994];
  wire _69006 = _69004 ^ _69005;
  wire _69007 = uncoded_block[1083] ^ uncoded_block[1092];
  wire _69008 = _56539 ^ _69007;
  wire _69009 = _69006 ^ _69008;
  wire _69010 = uncoded_block[1159] ^ uncoded_block[1203];
  wire _69011 = uncoded_block[1218] ^ uncoded_block[1244];
  wire _69012 = _69010 ^ _69011;
  wire _69013 = uncoded_block[1247] ^ uncoded_block[1278];
  wire _69014 = uncoded_block[1293] ^ uncoded_block[1314];
  wire _69015 = _69013 ^ _69014;
  wire _69016 = _69012 ^ _69015;
  wire _69017 = _69009 ^ _69016;
  wire _69018 = uncoded_block[1350] ^ uncoded_block[1390];
  wire _69019 = uncoded_block[1393] ^ uncoded_block[1429];
  wire _69020 = _69018 ^ _69019;
  wire _69021 = uncoded_block[1465] ^ uncoded_block[1514];
  wire _69022 = uncoded_block[1517] ^ uncoded_block[1536];
  wire _69023 = _69021 ^ _69022;
  wire _69024 = _69020 ^ _69023;
  wire _69025 = uncoded_block[1550] ^ uncoded_block[1592];
  wire _69026 = uncoded_block[1636] ^ uncoded_block[1668];
  wire _69027 = _69025 ^ _69026;
  wire _69028 = _69027 ^ uncoded_block[1669];
  wire _69029 = _69024 ^ _69028;
  wire _69030 = _69017 ^ _69029;
  wire _69031 = _69003 ^ _69030;
  wire _69032 = uncoded_block[18] ^ uncoded_block[26];
  wire _69033 = uncoded_block[83] ^ uncoded_block[94];
  wire _69034 = _69032 ^ _69033;
  wire _69035 = uncoded_block[120] ^ uncoded_block[166];
  wire _69036 = _69035 ^ _4766;
  wire _69037 = _69034 ^ _69036;
  wire _69038 = _46580 ^ _63796;
  wire _69039 = _38366 ^ _5580;
  wire _69040 = _69038 ^ _69039;
  wire _69041 = _69037 ^ _69040;
  wire _69042 = uncoded_block[457] ^ uncoded_block[492];
  wire _69043 = uncoded_block[525] ^ uncoded_block[541];
  wire _69044 = _69042 ^ _69043;
  wire _69045 = uncoded_block[568] ^ uncoded_block[578];
  wire _69046 = uncoded_block[659] ^ uncoded_block[675];
  wire _69047 = _69045 ^ _69046;
  wire _69048 = _69044 ^ _69047;
  wire _69049 = uncoded_block[692] ^ uncoded_block[754];
  wire _69050 = uncoded_block[770] ^ uncoded_block[781];
  wire _69051 = _69049 ^ _69050;
  wire _69052 = uncoded_block[782] ^ uncoded_block[840];
  wire _69053 = uncoded_block[855] ^ uncoded_block[902];
  wire _69054 = _69052 ^ _69053;
  wire _69055 = _69051 ^ _69054;
  wire _69056 = _69048 ^ _69055;
  wire _69057 = _69041 ^ _69056;
  wire _69058 = uncoded_block[941] ^ uncoded_block[950];
  wire _69059 = uncoded_block[983] ^ uncoded_block[1004];
  wire _69060 = _69058 ^ _69059;
  wire _69061 = uncoded_block[1050] ^ uncoded_block[1071];
  wire _69062 = uncoded_block[1082] ^ uncoded_block[1140];
  wire _69063 = _69061 ^ _69062;
  wire _69064 = _69060 ^ _69063;
  wire _69065 = uncoded_block[1163] ^ uncoded_block[1179];
  wire _69066 = uncoded_block[1220] ^ uncoded_block[1233];
  wire _69067 = _69065 ^ _69066;
  wire _69068 = uncoded_block[1241] ^ uncoded_block[1282];
  wire _69069 = _69068 ^ _61024;
  wire _69070 = _69067 ^ _69069;
  wire _69071 = _69064 ^ _69070;
  wire _69072 = uncoded_block[1335] ^ uncoded_block[1381];
  wire _69073 = _69072 ^ _3850;
  wire _69074 = uncoded_block[1441] ^ uncoded_block[1475];
  wire _69075 = uncoded_block[1519] ^ uncoded_block[1594];
  wire _69076 = _69074 ^ _69075;
  wire _69077 = _69073 ^ _69076;
  wire _69078 = uncoded_block[1602] ^ uncoded_block[1627];
  wire _69079 = uncoded_block[1629] ^ uncoded_block[1656];
  wire _69080 = _69078 ^ _69079;
  wire _69081 = _69080 ^ uncoded_block[1671];
  wire _69082 = _69077 ^ _69081;
  wire _69083 = _69071 ^ _69082;
  wire _69084 = _69057 ^ _69083;
  wire _69085 = uncoded_block[22] ^ uncoded_block[36];
  wire _69086 = uncoded_block[40] ^ uncoded_block[62];
  wire _69087 = _69085 ^ _69086;
  wire _69088 = uncoded_block[67] ^ uncoded_block[79];
  wire _69089 = uncoded_block[133] ^ uncoded_block[165];
  wire _69090 = _69088 ^ _69089;
  wire _69091 = _69087 ^ _69090;
  wire _69092 = uncoded_block[170] ^ uncoded_block[188];
  wire _69093 = _69092 ^ _4773;
  wire _69094 = uncoded_block[233] ^ uncoded_block[254];
  wire _69095 = uncoded_block[275] ^ uncoded_block[292];
  wire _69096 = _69094 ^ _69095;
  wire _69097 = _69093 ^ _69096;
  wire _69098 = _69091 ^ _69097;
  wire _69099 = _8051 ^ _62858;
  wire _69100 = uncoded_block[351] ^ uncoded_block[433];
  wire _69101 = uncoded_block[442] ^ uncoded_block[459];
  wire _69102 = _69100 ^ _69101;
  wire _69103 = _69099 ^ _69102;
  wire _69104 = uncoded_block[466] ^ uncoded_block[486];
  wire _69105 = uncoded_block[518] ^ uncoded_block[543];
  wire _69106 = _69104 ^ _69105;
  wire _69107 = uncoded_block[546] ^ uncoded_block[584];
  wire _69108 = _69107 ^ _6957;
  wire _69109 = _69106 ^ _69108;
  wire _69110 = _69103 ^ _69109;
  wire _69111 = _69098 ^ _69110;
  wire _69112 = uncoded_block[617] ^ uncoded_block[626];
  wire _69113 = uncoded_block[646] ^ uncoded_block[677];
  wire _69114 = _69112 ^ _69113;
  wire _69115 = _35635 ^ _58817;
  wire _69116 = _69114 ^ _69115;
  wire _69117 = uncoded_block[738] ^ uncoded_block[777];
  wire _69118 = uncoded_block[805] ^ uncoded_block[813];
  wire _69119 = _69117 ^ _69118;
  wire _69120 = uncoded_block[829] ^ uncoded_block[856];
  wire _69121 = uncoded_block[869] ^ uncoded_block[874];
  wire _69122 = _69120 ^ _69121;
  wire _69123 = _69119 ^ _69122;
  wire _69124 = _69116 ^ _69123;
  wire _69125 = uncoded_block[900] ^ uncoded_block[916];
  wire _69126 = uncoded_block[931] ^ uncoded_block[991];
  wire _69127 = _69125 ^ _69126;
  wire _69128 = _3664 ^ _36938;
  wire _69129 = _69127 ^ _69128;
  wire _69130 = uncoded_block[1057] ^ uncoded_block[1082];
  wire _69131 = _69130 ^ _53242;
  wire _69132 = uncoded_block[1119] ^ uncoded_block[1144];
  wire _69133 = uncoded_block[1153] ^ uncoded_block[1175];
  wire _69134 = _69132 ^ _69133;
  wire _69135 = _69131 ^ _69134;
  wire _69136 = _69129 ^ _69135;
  wire _69137 = _69124 ^ _69136;
  wire _69138 = _69111 ^ _69137;
  wire _69139 = uncoded_block[1180] ^ uncoded_block[1216];
  wire _69140 = uncoded_block[1249] ^ uncoded_block[1259];
  wire _69141 = _69139 ^ _69140;
  wire _69142 = uncoded_block[1269] ^ uncoded_block[1277];
  wire _69143 = uncoded_block[1374] ^ uncoded_block[1383];
  wire _69144 = _69142 ^ _69143;
  wire _69145 = _69141 ^ _69144;
  wire _69146 = uncoded_block[1396] ^ uncoded_block[1442];
  wire _69147 = uncoded_block[1443] ^ uncoded_block[1490];
  wire _69148 = _69146 ^ _69147;
  wire _69149 = uncoded_block[1542] ^ uncoded_block[1552];
  wire _69150 = _60098 ^ _69149;
  wire _69151 = _69148 ^ _69150;
  wire _69152 = _69145 ^ _69151;
  wire _69153 = _29986 ^ _47625;
  wire _69154 = uncoded_block[1601] ^ uncoded_block[1609];
  wire _69155 = uncoded_block[1622] ^ uncoded_block[1670];
  wire _69156 = _69154 ^ _69155;
  wire _69157 = _69153 ^ _69156;
  wire _69158 = _69157 ^ uncoded_block[1707];
  wire _69159 = _69152 ^ _69158;
  wire _69160 = _69138 ^ _69159;
  wire _69161 = _61399 ^ _18076;
  wire _69162 = uncoded_block[130] ^ uncoded_block[170];
  wire _69163 = uncoded_block[192] ^ uncoded_block[216];
  wire _69164 = _69162 ^ _69163;
  wire _69165 = _69161 ^ _69164;
  wire _69166 = uncoded_block[234] ^ uncoded_block[278];
  wire _69167 = uncoded_block[294] ^ uncoded_block[311];
  wire _69168 = _69166 ^ _69167;
  wire _69169 = uncoded_block[347] ^ uncoded_block[377];
  wire _69170 = uncoded_block[436] ^ uncoded_block[446];
  wire _69171 = _69169 ^ _69170;
  wire _69172 = _69168 ^ _69171;
  wire _69173 = _69165 ^ _69172;
  wire _69174 = uncoded_block[468] ^ uncoded_block[505];
  wire _69175 = uncoded_block[520] ^ uncoded_block[556];
  wire _69176 = _69174 ^ _69175;
  wire _69177 = uncoded_block[621] ^ uncoded_block[649];
  wire _69178 = _61454 ^ _69177;
  wire _69179 = _69176 ^ _69178;
  wire _69180 = uncoded_block[724] ^ uncoded_block[740];
  wire _69181 = _61459 ^ _69180;
  wire _69182 = uncoded_block[807] ^ uncoded_block[825];
  wire _69183 = uncoded_block[841] ^ uncoded_block[872];
  wire _69184 = _69182 ^ _69183;
  wire _69185 = _69181 ^ _69184;
  wire _69186 = _69179 ^ _69185;
  wire _69187 = _69173 ^ _69186;
  wire _69188 = uncoded_block[903] ^ uncoded_block[922];
  wire _69189 = _69188 ^ _12737;
  wire _69190 = uncoded_block[1004] ^ uncoded_block[1050];
  wire _69191 = uncoded_block[1085] ^ uncoded_block[1102];
  wire _69192 = _69190 ^ _69191;
  wire _69193 = _69189 ^ _69192;
  wire _69194 = uncoded_block[1137] ^ uncoded_block[1155];
  wire _69195 = uncoded_block[1183] ^ uncoded_block[1215];
  wire _69196 = _69194 ^ _69195;
  wire _69197 = uncoded_block[1262] ^ uncoded_block[1279];
  wire _69198 = _17907 ^ _69197;
  wire _69199 = _69196 ^ _69198;
  wire _69200 = _69193 ^ _69199;
  wire _69201 = uncoded_block[1288] ^ uncoded_block[1317];
  wire _69202 = uncoded_block[1361] ^ uncoded_block[1387];
  wire _69203 = _69201 ^ _69202;
  wire _69204 = uncoded_block[1425] ^ uncoded_block[1468];
  wire _69205 = uncoded_block[1534] ^ uncoded_block[1545];
  wire _69206 = _69204 ^ _69205;
  wire _69207 = _69203 ^ _69206;
  wire _69208 = uncoded_block[1581] ^ uncoded_block[1601];
  wire _69209 = uncoded_block[1608] ^ uncoded_block[1651];
  wire _69210 = _69208 ^ _69209;
  wire _69211 = _69210 ^ uncoded_block[1685];
  wire _69212 = _69207 ^ _69211;
  wire _69213 = _69200 ^ _69212;
  wire _69214 = _69187 ^ _69213;
  wire _69215 = uncoded_block[47] ^ uncoded_block[51];
  wire _69216 = _69215 ^ _64780;
  wire _69217 = uncoded_block[194] ^ uncoded_block[206];
  wire _69218 = _64781 ^ _69217;
  wire _69219 = _69216 ^ _69218;
  wire _69220 = _64787 ^ _64792;
  wire _69221 = uncoded_block[363] ^ uncoded_block[389];
  wire _69222 = uncoded_block[407] ^ uncoded_block[428];
  wire _69223 = _69221 ^ _69222;
  wire _69224 = _69220 ^ _69223;
  wire _69225 = _69219 ^ _69224;
  wire _69226 = _64799 ^ _65947;
  wire _69227 = uncoded_block[572] ^ uncoded_block[593];
  wire _69228 = _69227 ^ _9340;
  wire _69229 = _69226 ^ _69228;
  wire _69230 = _64810 ^ _60534;
  wire _69231 = uncoded_block[835] ^ uncoded_block[857];
  wire _69232 = _64814 ^ _69231;
  wire _69233 = _69230 ^ _69232;
  wire _69234 = _69229 ^ _69233;
  wire _69235 = _69225 ^ _69234;
  wire _69236 = uncoded_block[921] ^ uncoded_block[933];
  wire _69237 = uncoded_block[948] ^ uncoded_block[999];
  wire _69238 = _69236 ^ _69237;
  wire _69239 = uncoded_block[1063] ^ uncoded_block[1076];
  wire _69240 = _49571 ^ _69239;
  wire _69241 = _69238 ^ _69240;
  wire _69242 = uncoded_block[1162] ^ uncoded_block[1212];
  wire _69243 = _64829 ^ _69242;
  wire _69244 = uncoded_block[1242] ^ uncoded_block[1303];
  wire _69245 = _66623 ^ _69244;
  wire _69246 = _69243 ^ _69245;
  wire _69247 = _69241 ^ _69246;
  wire _69248 = uncoded_block[1431] ^ uncoded_block[1448];
  wire _69249 = _64841 ^ _69248;
  wire _69250 = uncoded_block[1464] ^ uncoded_block[1484];
  wire _69251 = uncoded_block[1495] ^ uncoded_block[1532];
  wire _69252 = _69250 ^ _69251;
  wire _69253 = _69249 ^ _69252;
  wire _69254 = uncoded_block[1577] ^ uncoded_block[1614];
  wire _69255 = uncoded_block[1652] ^ uncoded_block[1690];
  wire _69256 = _69254 ^ _69255;
  wire _69257 = _69256 ^ uncoded_block[1708];
  wire _69258 = _69253 ^ _69257;
  wire _69259 = _69247 ^ _69258;
  wire _69260 = _69235 ^ _69259;
  wire _69261 = uncoded_block[30] ^ uncoded_block[57];
  wire _69262 = uncoded_block[78] ^ uncoded_block[95];
  wire _69263 = _69261 ^ _69262;
  wire _69264 = uncoded_block[119] ^ uncoded_block[142];
  wire _69265 = uncoded_block[143] ^ uncoded_block[172];
  wire _69266 = _69264 ^ _69265;
  wire _69267 = _69263 ^ _69266;
  wire _69268 = uncoded_block[183] ^ uncoded_block[218];
  wire _69269 = _69268 ^ _44837;
  wire _69270 = uncoded_block[271] ^ uncoded_block[307];
  wire _69271 = _69270 ^ _63045;
  wire _69272 = _69269 ^ _69271;
  wire _69273 = _69267 ^ _69272;
  wire _69274 = uncoded_block[367] ^ uncoded_block[399];
  wire _69275 = _1029 ^ _69274;
  wire _69276 = uncoded_block[410] ^ uncoded_block[443];
  wire _69277 = uncoded_block[449] ^ uncoded_block[477];
  wire _69278 = _69276 ^ _69277;
  wire _69279 = _69275 ^ _69278;
  wire _69280 = uncoded_block[499] ^ uncoded_block[513];
  wire _69281 = _69280 ^ _32722;
  wire _69282 = uncoded_block[575] ^ uncoded_block[602];
  wire _69283 = _69282 ^ _63067;
  wire _69284 = _69281 ^ _69283;
  wire _69285 = _69279 ^ _69284;
  wire _69286 = _69273 ^ _69285;
  wire _69287 = _60981 ^ _318;
  wire _69288 = uncoded_block[691] ^ uncoded_block[743];
  wire _69289 = _69288 ^ _1217;
  wire _69290 = _69287 ^ _69289;
  wire _69291 = _22071 ^ _26164;
  wire _69292 = uncoded_block[856] ^ uncoded_block[924];
  wire _69293 = uncoded_block[930] ^ uncoded_block[938];
  wire _69294 = _69292 ^ _69293;
  wire _69295 = _69291 ^ _69294;
  wire _69296 = _69290 ^ _69295;
  wire _69297 = uncoded_block[992] ^ uncoded_block[1025];
  wire _69298 = _42022 ^ _69297;
  wire _69299 = uncoded_block[1079] ^ uncoded_block[1094];
  wire _69300 = _63104 ^ _69299;
  wire _69301 = _69298 ^ _69300;
  wire _69302 = uncoded_block[1129] ^ uncoded_block[1140];
  wire _69303 = _7132 ^ _69302;
  wire _69304 = uncoded_block[1172] ^ uncoded_block[1203];
  wire _69305 = uncoded_block[1207] ^ uncoded_block[1225];
  wire _69306 = _69304 ^ _69305;
  wire _69307 = _69303 ^ _69306;
  wire _69308 = _69301 ^ _69307;
  wire _69309 = _69296 ^ _69308;
  wire _69310 = _69286 ^ _69309;
  wire _69311 = uncoded_block[1249] ^ uncoded_block[1272];
  wire _69312 = _69311 ^ _10646;
  wire _69313 = _61031 ^ _49067;
  wire _69314 = _69312 ^ _69313;
  wire _69315 = uncoded_block[1392] ^ uncoded_block[1400];
  wire _69316 = _69315 ^ _63137;
  wire _69317 = _63138 ^ _63142;
  wire _69318 = _69316 ^ _69317;
  wire _69319 = _69314 ^ _69318;
  wire _69320 = uncoded_block[1470] ^ uncoded_block[1488];
  wire _69321 = uncoded_block[1491] ^ uncoded_block[1511];
  wire _69322 = _69320 ^ _69321;
  wire _69323 = uncoded_block[1621] ^ uncoded_block[1683];
  wire _69324 = _69323 ^ _33025;
  wire _69325 = _69322 ^ _69324;
  wire _69326 = _69325 ^ uncoded_block[1722];
  wire _69327 = _69319 ^ _69326;
  wire _69328 = _69310 ^ _69327;
  wire _69329 = _35101 ^ _21873;
  wire _69330 = _23 ^ _4726;
  wire _69331 = _1703 ^ _2472;
  wire _69332 = _69330 ^ _69331;
  wire _69333 = _69329 ^ _69332;
  wire _69334 = _68441 ^ _69333;
  wire _69335 = _14586 ^ _2487;
  wire _69336 = _51488 ^ _69335;
  wire _69337 = _68449 ^ _69336;
  wire _69338 = _14591 ^ _3249;
  wire _69339 = _15097 ^ _4031;
  wire _69340 = _69338 ^ _69339;
  wire _69341 = _68455 ^ _42599;
  wire _69342 = _69340 ^ _69341;
  wire _69343 = _69337 ^ _69342;
  wire _69344 = _69334 ^ _69343;
  wire _69345 = _4750 ^ _23269;
  wire _69346 = _69345 ^ _35514;
  wire _69347 = _1735 ^ _8581;
  wire _69348 = _9729 ^ _11924;
  wire _69349 = _69347 ^ _69348;
  wire _69350 = _69346 ^ _69349;
  wire _69351 = _55477 ^ _9186;
  wire _69352 = _69351 ^ _15119;
  wire _69353 = _14087 ^ _32646;
  wire _69354 = _69352 ^ _69353;
  wire _69355 = _69350 ^ _69354;
  wire _69356 = _14093 ^ _24646;
  wire _69357 = _18111 ^ _3283;
  wire _69358 = _3284 ^ _4068;
  wire _69359 = _69357 ^ _69358;
  wire _69360 = _69356 ^ _69359;
  wire _69361 = _11405 ^ _12483;
  wire _69362 = _39141 ^ _69361;
  wire _69363 = _22376 ^ _25100;
  wire _69364 = _69362 ^ _69363;
  wire _69365 = _69360 ^ _69364;
  wire _69366 = _69355 ^ _69365;
  wire _69367 = _69344 ^ _69366;
  wire _69368 = _1781 ^ _2556;
  wire _69369 = _21466 ^ _69368;
  wire _69370 = _60179 ^ _69369;
  wire _69371 = _5512 ^ _10303;
  wire _69372 = _68494 ^ _69371;
  wire _69373 = _68493 ^ _69372;
  wire _69374 = _69370 ^ _69373;
  wire _69375 = _5515 ^ _40716;
  wire _69376 = _69375 ^ _39547;
  wire _69377 = _32675 ^ _60193;
  wire _69378 = _69376 ^ _69377;
  wire _69379 = _145 ^ _6850;
  wire _69380 = _69379 ^ _39558;
  wire _69381 = _9242 ^ _6218;
  wire _69382 = _68505 ^ _69381;
  wire _69383 = _69380 ^ _69382;
  wire _69384 = _69378 ^ _69383;
  wire _69385 = _69374 ^ _69384;
  wire _69386 = _1023 ^ _2599;
  wire _69387 = _2601 ^ _20554;
  wire _69388 = _69386 ^ _69387;
  wire _69389 = _35170 ^ _5548;
  wire _69390 = _69389 ^ _37596;
  wire _69391 = _69388 ^ _69390;
  wire _69392 = _4149 ^ _12006;
  wire _69393 = _69392 ^ _30137;
  wire _69394 = _68516 ^ _69393;
  wire _69395 = _69391 ^ _69394;
  wire _69396 = _60214 ^ _47373;
  wire _69397 = _14160 ^ _2633;
  wire _69398 = _1062 ^ _34771;
  wire _69399 = _69397 ^ _69398;
  wire _69400 = _69396 ^ _69399;
  wire _69401 = _10352 ^ _23349;
  wire _69402 = _69401 ^ _68529;
  wire _69403 = uncoded_block[464] ^ uncoded_block[468];
  wire _69404 = _13662 ^ _69403;
  wire _69405 = _39982 ^ _69404;
  wire _69406 = _69402 ^ _69405;
  wire _69407 = _69400 ^ _69406;
  wire _69408 = _69395 ^ _69407;
  wire _69409 = _69385 ^ _69408;
  wire _69410 = _69367 ^ _69409;
  wire _69411 = _33987 ^ _4897;
  wire _69412 = _21527 ^ _69411;
  wire _69413 = _7516 ^ _21987;
  wire _69414 = _4905 ^ _1892;
  wire _69415 = _69413 ^ _69414;
  wire _69416 = _69412 ^ _69415;
  wire _69417 = _23370 ^ _1108;
  wire _69418 = _33579 ^ _69417;
  wire _69419 = _9301 ^ _6929;
  wire _69420 = _69419 ^ _23374;
  wire _69421 = _69418 ^ _69420;
  wire _69422 = _69416 ^ _69421;
  wire _69423 = _32324 ^ _2687;
  wire _69424 = _69423 ^ _60245;
  wire _69425 = _9320 ^ _3467;
  wire _69426 = _69425 ^ _68554;
  wire _69427 = _69424 ^ _69426;
  wire _69428 = _1931 ^ _1133;
  wire _69429 = _69428 ^ _58464;
  wire _69430 = _17721 ^ _2707;
  wire _69431 = _15753 ^ _69430;
  wire _69432 = _69429 ^ _69431;
  wire _69433 = _69427 ^ _69432;
  wire _69434 = _69422 ^ _69433;
  wire _69435 = _3489 ^ _14218;
  wire _69436 = _69435 ^ _68566;
  wire _69437 = _15261 ^ _5658;
  wire _69438 = _11538 ^ _69437;
  wire _69439 = _69436 ^ _69438;
  wire _69440 = _58804 ^ _36018;
  wire _69441 = _18705 ^ _15270;
  wire _69442 = _40796 ^ _69441;
  wire _69443 = _69440 ^ _69442;
  wire _69444 = _69439 ^ _69443;
  wire _69445 = _13726 ^ _311;
  wire _69446 = _69445 ^ _16254;
  wire _69447 = _69446 ^ _68577;
  wire _69448 = _329 ^ _17258;
  wire _69449 = _68578 ^ _69448;
  wire _69450 = _5685 ^ _33204;
  wire _69451 = _69450 ^ _55603;
  wire _69452 = _69449 ^ _69451;
  wire _69453 = _69447 ^ _69452;
  wire _69454 = _69444 ^ _69453;
  wire _69455 = _69434 ^ _69454;
  wire _69456 = _6367 ^ _4283;
  wire _69457 = _7002 ^ _1996;
  wire _69458 = _69456 ^ _69457;
  wire _69459 = _69458 ^ _68592;
  wire _69460 = uncoded_block[761] ^ uncoded_block[766];
  wire _69461 = _3556 ^ _69460;
  wire _69462 = _53732 ^ _69461;
  wire _69463 = _17776 ^ _14271;
  wire _69464 = _69463 ^ _41207;
  wire _69465 = _69462 ^ _69464;
  wire _69466 = _69459 ^ _69465;
  wire _69467 = _19705 ^ _2015;
  wire _69468 = _69467 ^ _58512;
  wire _69469 = _14282 ^ _7029;
  wire _69470 = _4317 ^ _12127;
  wire _69471 = _69469 ^ _69470;
  wire _69472 = _69468 ^ _69471;
  wire _69473 = uncoded_block[812] ^ uncoded_block[815];
  wire _69474 = _1238 ^ _69473;
  wire _69475 = _4325 ^ _2809;
  wire _69476 = _69474 ^ _69475;
  wire _69477 = _2813 ^ _57415;
  wire _69478 = _69476 ^ _69477;
  wire _69479 = _69472 ^ _69478;
  wire _69480 = _69466 ^ _69479;
  wire _69481 = _47836 ^ _1256;
  wire _69482 = _1257 ^ _2044;
  wire _69483 = _69481 ^ _69482;
  wire _69484 = _15330 ^ _23010;
  wire _69485 = _69484 ^ _14303;
  wire _69486 = _69483 ^ _69485;
  wire _69487 = _9953 ^ _41628;
  wire _69488 = _69487 ^ _48967;
  wire _69489 = _1277 ^ _20704;
  wire _69490 = _1280 ^ _19252;
  wire _69491 = _69489 ^ _69490;
  wire _69492 = _69488 ^ _69491;
  wire _69493 = _69486 ^ _69492;
  wire _69494 = _68624 ^ _2076;
  wire _69495 = _448 ^ _21649;
  wire _69496 = _69494 ^ _69495;
  wire _69497 = _58542 ^ _8842;
  wire _69498 = _454 ^ _69497;
  wire _69499 = _69496 ^ _69498;
  wire _69500 = _22566 ^ _22568;
  wire _69501 = _467 ^ _5112;
  wire _69502 = _17836 ^ _10537;
  wire _69503 = _69501 ^ _69502;
  wire _69504 = _69500 ^ _69503;
  wire _69505 = _69499 ^ _69504;
  wire _69506 = _69493 ^ _69505;
  wire _69507 = _69480 ^ _69506;
  wire _69508 = _69455 ^ _69507;
  wire _69509 = _69410 ^ _69508;
  wire _69510 = _12186 ^ _23938;
  wire _69511 = _3663 ^ _8293;
  wire _69512 = _69510 ^ _69511;
  wire _69513 = _7691 ^ _43085;
  wire _69514 = _13283 ^ _5131;
  wire _69515 = _69513 ^ _69514;
  wire _69516 = _69512 ^ _69515;
  wire _69517 = uncoded_block[1016] ^ uncoded_block[1021];
  wire _69518 = _69517 ^ _5137;
  wire _69519 = _69518 ^ _60338;
  wire _69520 = _7707 ^ _48641;
  wire _69521 = _59337 ^ _518;
  wire _69522 = _69520 ^ _69521;
  wire _69523 = _69519 ^ _69522;
  wire _69524 = _69516 ^ _69523;
  wire _69525 = _13295 ^ _38137;
  wire _69526 = _69525 ^ _68656;
  wire _69527 = _530 ^ _20753;
  wire _69528 = _68657 ^ _69527;
  wire _69529 = _69526 ^ _69528;
  wire _69530 = _48266 ^ _10580;
  wire _69531 = _15405 ^ _14372;
  wire _69532 = _69531 ^ _41682;
  wire _69533 = _69530 ^ _69532;
  wire _69534 = _69529 ^ _69533;
  wire _69535 = _69524 ^ _69534;
  wire _69536 = _68665 ^ _14886;
  wire _69537 = _62076 ^ _8929;
  wire _69538 = _4462 ^ _4465;
  wire _69539 = _69537 ^ _69538;
  wire _69540 = _69536 ^ _69539;
  wire _69541 = _65826 ^ _40539;
  wire _69542 = _19327 ^ _69541;
  wire _69543 = _584 ^ _17396;
  wire _69544 = _2195 ^ _35354;
  wire _69545 = _69543 ^ _69544;
  wire _69546 = _69542 ^ _69545;
  wire _69547 = _69540 ^ _69546;
  wire _69548 = _15431 ^ _2210;
  wire _69549 = _11171 ^ _1428;
  wire _69550 = _69548 ^ _69549;
  wire _69551 = _60375 ^ _69550;
  wire _69552 = _31228 ^ _13360;
  wire _69553 = _30775 ^ _69552;
  wire _69554 = _60381 ^ _69553;
  wire _69555 = _69551 ^ _69554;
  wire _69556 = _69547 ^ _69555;
  wire _69557 = _69535 ^ _69556;
  wire _69558 = _2230 ^ _59168;
  wire _69559 = uncoded_block[1254] ^ uncoded_block[1259];
  wire _69560 = _69559 ^ _30361;
  wire _69561 = _69558 ^ _69560;
  wire _69562 = _26718 ^ _1463;
  wire _69563 = _9534 ^ _69562;
  wire _69564 = _69561 ^ _69563;
  wire _69565 = _27136 ^ _17427;
  wire _69566 = _4531 ^ _13915;
  wire _69567 = _4530 ^ _69566;
  wire _69568 = _69565 ^ _69567;
  wire _69569 = _69564 ^ _69568;
  wire _69570 = _8407 ^ _7805;
  wire _69571 = _68706 ^ _69570;
  wire _69572 = _3032 ^ _8413;
  wire _69573 = _3822 ^ _9564;
  wire _69574 = _69572 ^ _69573;
  wire _69575 = _69571 ^ _69574;
  wire _69576 = _60403 ^ _16443;
  wire _69577 = _12861 ^ _54880;
  wire _69578 = _69577 ^ _5286;
  wire _69579 = _69576 ^ _69578;
  wire _69580 = _69575 ^ _69579;
  wire _69581 = _69569 ^ _69580;
  wire _69582 = _68720 ^ _68725;
  wire _69583 = _21316 ^ _60413;
  wire _69584 = _69582 ^ _69583;
  wire _69585 = _68728 ^ _17961;
  wire _69586 = _1534 ^ _13432;
  wire _69587 = _68731 ^ _69586;
  wire _69588 = _69585 ^ _69587;
  wire _69589 = _69584 ^ _69588;
  wire _69590 = _6613 ^ _11246;
  wire _69591 = _20852 ^ _23176;
  wire _69592 = _69590 ^ _69591;
  wire _69593 = _35423 ^ _41757;
  wire _69594 = _3101 ^ _17980;
  wire _69595 = _69593 ^ _69594;
  wire _69596 = _69592 ^ _69595;
  wire _69597 = _1565 ^ _43955;
  wire _69598 = _3109 ^ _3894;
  wire _69599 = _69597 ^ _69598;
  wire _69600 = _23628 ^ _60435;
  wire _69601 = _69599 ^ _69600;
  wire _69602 = _69596 ^ _69601;
  wire _69603 = _69589 ^ _69602;
  wire _69604 = _69581 ^ _69603;
  wire _69605 = _69557 ^ _69604;
  wire _69606 = _36235 ^ _68755;
  wire _69607 = _60440 ^ _11832;
  wire _69608 = _69606 ^ _69607;
  wire _69609 = _25451 ^ _6664;
  wire _69610 = _40243 ^ _6673;
  wire _69611 = uncoded_block[1600] ^ uncoded_block[1604];
  wire _69612 = _11295 ^ _69611;
  wire _69613 = _69610 ^ _69612;
  wire _69614 = _69609 ^ _69613;
  wire _69615 = _69608 ^ _69614;
  wire _69616 = _68768 ^ _29557;
  wire _69617 = _33421 ^ _69616;
  wire _69618 = _1636 ^ _5388;
  wire _69619 = uncoded_block[1637] ^ uncoded_block[1641];
  wire _69620 = _69619 ^ _34255;
  wire _69621 = _69618 ^ _69620;
  wire _69622 = _69617 ^ _69621;
  wire _69623 = _42182 ^ _19465;
  wire _69624 = _9667 ^ _25030;
  wire _69625 = _69623 ^ _69624;
  wire _69626 = _69622 ^ _69625;
  wire _69627 = _69615 ^ _69626;
  wire _69628 = _3183 ^ _11321;
  wire _69629 = _69628 ^ _38681;
  wire _69630 = _14544 ^ _48779;
  wire _69631 = _69629 ^ _69630;
  wire _69632 = uncoded_block[1699] ^ uncoded_block[1705];
  wire _69633 = _69632 ^ _2437;
  wire _69634 = _55813 ^ _1677;
  wire _69635 = _69633 ^ _69634;
  wire _69636 = _69635 ^ uncoded_block[1722];
  wire _69637 = _69631 ^ _69636;
  wire _69638 = _69627 ^ _69637;
  wire _69639 = _69605 ^ _69638;
  wire _69640 = _69509 ^ _69639;
  wire _69641 = uncoded_block[0] ^ uncoded_block[25];
  wire _69642 = uncoded_block[38] ^ uncoded_block[78];
  wire _69643 = _69641 ^ _69642;
  wire _69644 = uncoded_block[116] ^ uncoded_block[147];
  wire _69645 = _58721 ^ _69644;
  wire _69646 = _69643 ^ _69645;
  wire _69647 = uncoded_block[184] ^ uncoded_block[224];
  wire _69648 = _59935 ^ _69647;
  wire _69649 = uncoded_block[231] ^ uncoded_block[247];
  wire _69650 = _69649 ^ _65353;
  wire _69651 = _69648 ^ _69650;
  wire _69652 = _69646 ^ _69651;
  wire _69653 = uncoded_block[340] ^ uncoded_block[364];
  wire _69654 = _16648 ^ _69653;
  wire _69655 = uncoded_block[380] ^ uncoded_block[413];
  wire _69656 = _69655 ^ _25150;
  wire _69657 = _69654 ^ _69656;
  wire _69658 = uncoded_block[482] ^ uncoded_block[520];
  wire _69659 = _29280 ^ _69658;
  wire _69660 = uncoded_block[521] ^ uncoded_block[545];
  wire _69661 = uncoded_block[565] ^ uncoded_block[581];
  wire _69662 = _69660 ^ _69661;
  wire _69663 = _69659 ^ _69662;
  wire _69664 = _69657 ^ _69663;
  wire _69665 = _69652 ^ _69664;
  wire _69666 = uncoded_block[606] ^ uncoded_block[621];
  wire _69667 = uncoded_block[623] ^ uncoded_block[647];
  wire _69668 = _69666 ^ _69667;
  wire _69669 = _18719 ^ _65372;
  wire _69670 = _69668 ^ _69669;
  wire _69671 = uncoded_block[765] ^ uncoded_block[790];
  wire _69672 = uncoded_block[795] ^ uncoded_block[803];
  wire _69673 = _69671 ^ _69672;
  wire _69674 = uncoded_block[848] ^ uncoded_block[860];
  wire _69675 = uncoded_block[863] ^ uncoded_block[905];
  wire _69676 = _69674 ^ _69675;
  wire _69677 = _69673 ^ _69676;
  wire _69678 = _69670 ^ _69677;
  wire _69679 = uncoded_block[919] ^ uncoded_block[933];
  wire _69680 = uncoded_block[967] ^ uncoded_block[984];
  wire _69681 = _69679 ^ _69680;
  wire _69682 = uncoded_block[1029] ^ uncoded_block[1052];
  wire _69683 = _62406 ^ _69682;
  wire _69684 = _69681 ^ _69683;
  wire _69685 = uncoded_block[1086] ^ uncoded_block[1127];
  wire _69686 = _49575 ^ _69685;
  wire _69687 = uncoded_block[1166] ^ uncoded_block[1175];
  wire _69688 = _50600 ^ _69687;
  wire _69689 = _69686 ^ _69688;
  wire _69690 = _69684 ^ _69689;
  wire _69691 = _69678 ^ _69690;
  wire _69692 = _69665 ^ _69691;
  wire _69693 = uncoded_block[1219] ^ uncoded_block[1230];
  wire _69694 = _5209 ^ _69693;
  wire _69695 = uncoded_block[1260] ^ uncoded_block[1266];
  wire _69696 = uncoded_block[1298] ^ uncoded_block[1313];
  wire _69697 = _69695 ^ _69696;
  wire _69698 = _69694 ^ _69697;
  wire _69699 = uncoded_block[1327] ^ uncoded_block[1346];
  wire _69700 = uncoded_block[1394] ^ uncoded_block[1406];
  wire _69701 = _69699 ^ _69700;
  wire _69702 = _60087 ^ _5309;
  wire _69703 = _69701 ^ _69702;
  wire _69704 = _69698 ^ _69703;
  wire _69705 = uncoded_block[1473] ^ uncoded_block[1493];
  wire _69706 = uncoded_block[1495] ^ uncoded_block[1579];
  wire _69707 = _69705 ^ _69706;
  wire _69708 = _7912 ^ _36687;
  wire _69709 = _69707 ^ _69708;
  wire _69710 = _3979 ^ uncoded_block[1715];
  wire _69711 = _69709 ^ _69710;
  wire _69712 = _69704 ^ _69711;
  wire _69713 = _69692 ^ _69712;
  wire _69714 = uncoded_block[5] ^ uncoded_block[28];
  wire _69715 = uncoded_block[77] ^ uncoded_block[104];
  wire _69716 = _69714 ^ _69715;
  wire _69717 = uncoded_block[183] ^ uncoded_block[202];
  wire _69718 = _71 ^ _69717;
  wire _69719 = _69716 ^ _69718;
  wire _69720 = uncoded_block[251] ^ uncoded_block[261];
  wire _69721 = uncoded_block[295] ^ uncoded_block[320];
  wire _69722 = _69720 ^ _69721;
  wire _69723 = uncoded_block[421] ^ uncoded_block[432];
  wire _69724 = _16664 ^ _69723;
  wire _69725 = _69722 ^ _69724;
  wire _69726 = _69719 ^ _69725;
  wire _69727 = uncoded_block[508] ^ uncoded_block[526];
  wire _69728 = _8111 ^ _69727;
  wire _69729 = uncoded_block[627] ^ uncoded_block[651];
  wire _69730 = _2715 ^ _69729;
  wire _69731 = _69728 ^ _69730;
  wire _69732 = uncoded_block[757] ^ uncoded_block[773];
  wire _69733 = _51599 ^ _69732;
  wire _69734 = uncoded_block[865] ^ uncoded_block[871];
  wire _69735 = _4322 ^ _69734;
  wire _69736 = _69733 ^ _69735;
  wire _69737 = _69731 ^ _69736;
  wire _69738 = _69726 ^ _69737;
  wire _69739 = uncoded_block[915] ^ uncoded_block[939];
  wire _69740 = uncoded_block[956] ^ uncoded_block[1002];
  wire _69741 = _69739 ^ _69740;
  wire _69742 = uncoded_block[1013] ^ uncoded_block[1034];
  wire _69743 = uncoded_block[1076] ^ uncoded_block[1148];
  wire _69744 = _69742 ^ _69743;
  wire _69745 = _69741 ^ _69744;
  wire _69746 = uncoded_block[1151] ^ uncoded_block[1177];
  wire _69747 = _69746 ^ _54471;
  wire _69748 = uncoded_block[1277] ^ uncoded_block[1302];
  wire _69749 = _59835 ^ _69748;
  wire _69750 = _69747 ^ _69749;
  wire _69751 = _69745 ^ _69750;
  wire _69752 = uncoded_block[1313] ^ uncoded_block[1343];
  wire _69753 = uncoded_block[1352] ^ uncoded_block[1397];
  wire _69754 = _69752 ^ _69753;
  wire _69755 = uncoded_block[1399] ^ uncoded_block[1436];
  wire _69756 = uncoded_block[1492] ^ uncoded_block[1560];
  wire _69757 = _69755 ^ _69756;
  wire _69758 = _69754 ^ _69757;
  wire _69759 = uncoded_block[1586] ^ uncoded_block[1593];
  wire _69760 = uncoded_block[1610] ^ uncoded_block[1698];
  wire _69761 = _69759 ^ _69760;
  wire _69762 = _69761 ^ uncoded_block[1712];
  wire _69763 = _69758 ^ _69762;
  wire _69764 = _69751 ^ _69763;
  wire _69765 = _69738 ^ _69764;
  wire _69766 = uncoded_block[10] ^ uncoded_block[51];
  wire _69767 = uncoded_block[56] ^ uncoded_block[107];
  wire _69768 = _69766 ^ _69767;
  wire _69769 = uncoded_block[116] ^ uncoded_block[157];
  wire _69770 = uncoded_block[172] ^ uncoded_block[186];
  wire _69771 = _69769 ^ _69770;
  wire _69772 = _69768 ^ _69771;
  wire _69773 = uncoded_block[255] ^ uncoded_block[276];
  wire _69774 = uncoded_block[305] ^ uncoded_block[324];
  wire _69775 = _69773 ^ _69774;
  wire _69776 = uncoded_block[402] ^ uncoded_block[425];
  wire _69777 = _29257 ^ _69776;
  wire _69778 = _69775 ^ _69777;
  wire _69779 = _69772 ^ _69778;
  wire _69780 = uncoded_block[531] ^ uncoded_block[547];
  wire _69781 = _4902 ^ _69780;
  wire _69782 = uncoded_block[561] ^ uncoded_block[596];
  wire _69783 = uncoded_block[630] ^ uncoded_block[643];
  wire _69784 = _69782 ^ _69783;
  wire _69785 = _69781 ^ _69784;
  wire _69786 = uncoded_block[723] ^ uncoded_block[813];
  wire _69787 = _62696 ^ _69786;
  wire _69788 = uncoded_block[824] ^ uncoded_block[857];
  wire _69789 = uncoded_block[868] ^ uncoded_block[939];
  wire _69790 = _69788 ^ _69789;
  wire _69791 = _69787 ^ _69790;
  wire _69792 = _69785 ^ _69791;
  wire _69793 = _69779 ^ _69792;
  wire _69794 = uncoded_block[954] ^ uncoded_block[1039];
  wire _69795 = _8841 ^ _69794;
  wire _69796 = uncoded_block[1053] ^ uncoded_block[1090];
  wire _69797 = uncoded_block[1107] ^ uncoded_block[1119];
  wire _69798 = _69796 ^ _69797;
  wire _69799 = _69795 ^ _69798;
  wire _69800 = uncoded_block[1155] ^ uncoded_block[1209];
  wire _69801 = _69800 ^ _23105;
  wire _69802 = uncoded_block[1224] ^ uncoded_block[1291];
  wire _69803 = uncoded_block[1305] ^ uncoded_block[1348];
  wire _69804 = _69802 ^ _69803;
  wire _69805 = _69801 ^ _69804;
  wire _69806 = _69799 ^ _69805;
  wire _69807 = uncoded_block[1371] ^ uncoded_block[1404];
  wire _69808 = uncoded_block[1413] ^ uncoded_block[1429];
  wire _69809 = _69807 ^ _69808;
  wire _69810 = uncoded_block[1499] ^ uncoded_block[1564];
  wire _69811 = uncoded_block[1586] ^ uncoded_block[1597];
  wire _69812 = _69810 ^ _69811;
  wire _69813 = _69809 ^ _69812;
  wire _69814 = uncoded_block[1655] ^ uncoded_block[1705];
  wire _69815 = _67850 ^ _69814;
  wire _69816 = _69815 ^ uncoded_block[1713];
  wire _69817 = _69813 ^ _69816;
  wire _69818 = _69806 ^ _69817;
  wire _69819 = _69793 ^ _69818;
  wire _69820 = uncoded_block[13] ^ uncoded_block[19];
  wire _69821 = _69820 ^ _34682;
  wire _69822 = uncoded_block[57] ^ uncoded_block[76];
  wire _69823 = uncoded_block[117] ^ uncoded_block[126];
  wire _69824 = _69822 ^ _69823;
  wire _69825 = _69821 ^ _69824;
  wire _69826 = uncoded_block[161] ^ uncoded_block[173];
  wire _69827 = _69826 ^ _58738;
  wire _69828 = _4095 ^ _61792;
  wire _69829 = _69827 ^ _69828;
  wire _69830 = _69825 ^ _69829;
  wire _69831 = uncoded_block[306] ^ uncoded_block[328];
  wire _69832 = _69831 ^ _173;
  wire _69833 = uncoded_block[379] ^ uncoded_block[402];
  wire _69834 = uncoded_block[403] ^ uncoded_block[429];
  wire _69835 = _69833 ^ _69834;
  wire _69836 = _69832 ^ _69835;
  wire _69837 = uncoded_block[467] ^ uncoded_block[494];
  wire _69838 = uncoded_block[495] ^ uncoded_block[535];
  wire _69839 = _69837 ^ _69838;
  wire _69840 = uncoded_block[540] ^ uncoded_block[548];
  wire _69841 = uncoded_block[565] ^ uncoded_block[597];
  wire _69842 = _69840 ^ _69841;
  wire _69843 = _69839 ^ _69842;
  wire _69844 = _69836 ^ _69843;
  wire _69845 = _69830 ^ _69844;
  wire _69846 = uncoded_block[612] ^ uncoded_block[634];
  wire _69847 = uncoded_block[635] ^ uncoded_block[644];
  wire _69848 = _69846 ^ _69847;
  wire _69849 = uncoded_block[697] ^ uncoded_block[710];
  wire _69850 = _69849 ^ _66715;
  wire _69851 = _69848 ^ _69850;
  wire _69852 = uncoded_block[750] ^ uncoded_block[793];
  wire _69853 = _69852 ^ _61860;
  wire _69854 = uncoded_block[872] ^ uncoded_block[891];
  wire _69855 = _66170 ^ _69854;
  wire _69856 = _69853 ^ _69855;
  wire _69857 = _69851 ^ _69856;
  wire _69858 = uncoded_block[925] ^ uncoded_block[940];
  wire _69859 = _69858 ^ _14329;
  wire _69860 = uncoded_block[968] ^ uncoded_block[1026];
  wire _69861 = uncoded_block[1043] ^ uncoded_block[1054];
  wire _69862 = _69860 ^ _69861;
  wire _69863 = _69859 ^ _69862;
  wire _69864 = uncoded_block[1120] ^ uncoded_block[1140];
  wire _69865 = _1378 ^ _69864;
  wire _69866 = uncoded_block[1159] ^ uncoded_block[1210];
  wire _69867 = uncoded_block[1221] ^ uncoded_block[1238];
  wire _69868 = _69866 ^ _69867;
  wire _69869 = _69865 ^ _69868;
  wire _69870 = _69863 ^ _69869;
  wire _69871 = _69857 ^ _69870;
  wire _69872 = _69845 ^ _69871;
  wire _69873 = uncoded_block[1240] ^ uncoded_block[1278];
  wire _69874 = _69873 ^ _9545;
  wire _69875 = uncoded_block[1309] ^ uncoded_block[1352];
  wire _69876 = uncoded_block[1355] ^ uncoded_block[1372];
  wire _69877 = _69875 ^ _69876;
  wire _69878 = _69874 ^ _69877;
  wire _69879 = uncoded_block[1395] ^ uncoded_block[1408];
  wire _69880 = _69879 ^ _66520;
  wire _69881 = _66523 ^ _38247;
  wire _69882 = _69880 ^ _69881;
  wire _69883 = _69878 ^ _69882;
  wire _69884 = uncoded_block[1568] ^ uncoded_block[1587];
  wire _69885 = uncoded_block[1592] ^ uncoded_block[1600];
  wire _69886 = _69884 ^ _69885;
  wire _69887 = _804 ^ _67554;
  wire _69888 = _69886 ^ _69887;
  wire _69889 = uncoded_block[1691] ^ uncoded_block[1706];
  wire _69890 = _69889 ^ uncoded_block[1716];
  wire _69891 = _69888 ^ _69890;
  wire _69892 = _69883 ^ _69891;
  wire _69893 = _69872 ^ _69892;
  wire _69894 = uncoded_block[47] ^ uncoded_block[66];
  wire _69895 = _14565 ^ _69894;
  wire _69896 = uncoded_block[73] ^ uncoded_block[105];
  wire _69897 = _69896 ^ _4034;
  wire _69898 = _69895 ^ _69897;
  wire _69899 = uncoded_block[124] ^ uncoded_block[198];
  wire _69900 = _69899 ^ _64342;
  wire _69901 = uncoded_block[225] ^ uncoded_block[254];
  wire _69902 = uncoded_block[269] ^ uncoded_block[284];
  wire _69903 = _69901 ^ _69902;
  wire _69904 = _69900 ^ _69903;
  wire _69905 = _69898 ^ _69904;
  wire _69906 = uncoded_block[337] ^ uncoded_block[379];
  wire _69907 = _64350 ^ _69906;
  wire _69908 = uncoded_block[390] ^ uncoded_block[412];
  wire _69909 = uncoded_block[415] ^ uncoded_block[439];
  wire _69910 = _69908 ^ _69909;
  wire _69911 = _69907 ^ _69910;
  wire _69912 = uncoded_block[449] ^ uncoded_block[484];
  wire _69913 = uncoded_block[499] ^ uncoded_block[523];
  wire _69914 = _69912 ^ _69913;
  wire _69915 = uncoded_block[526] ^ uncoded_block[546];
  wire _69916 = _69915 ^ _1130;
  wire _69917 = _69914 ^ _69916;
  wire _69918 = _69911 ^ _69917;
  wire _69919 = _69905 ^ _69918;
  wire _69920 = uncoded_block[599] ^ uncoded_block[645];
  wire _69921 = uncoded_block[680] ^ uncoded_block[692];
  wire _69922 = _69920 ^ _69921;
  wire _69923 = uncoded_block[718] ^ uncoded_block[736];
  wire _69924 = _69923 ^ _64383;
  wire _69925 = _69922 ^ _69924;
  wire _69926 = _61155 ^ _5066;
  wire _69927 = uncoded_block[882] ^ uncoded_block[895];
  wire _69928 = uncoded_block[902] ^ uncoded_block[939];
  wire _69929 = _69927 ^ _69928;
  wire _69930 = _69926 ^ _69929;
  wire _69931 = _69925 ^ _69930;
  wire _69932 = uncoded_block[977] ^ uncoded_block[1042];
  wire _69933 = _11643 ^ _69932;
  wire _69934 = _23966 ^ _64406;
  wire _69935 = _69933 ^ _69934;
  wire _69936 = uncoded_block[1121] ^ uncoded_block[1146];
  wire _69937 = uncoded_block[1176] ^ uncoded_block[1193];
  wire _69938 = _69936 ^ _69937;
  wire _69939 = uncoded_block[1202] ^ uncoded_block[1252];
  wire _69940 = uncoded_block[1258] ^ uncoded_block[1264];
  wire _69941 = _69939 ^ _69940;
  wire _69942 = _69938 ^ _69941;
  wire _69943 = _69935 ^ _69942;
  wire _69944 = _69931 ^ _69943;
  wire _69945 = _69919 ^ _69944;
  wire _69946 = uncoded_block[1297] ^ uncoded_block[1318];
  wire _69947 = _69946 ^ _11207;
  wire _69948 = _64425 ^ _69202;
  wire _69949 = _69947 ^ _69948;
  wire _69950 = uncoded_block[1440] ^ uncoded_block[1461];
  wire _69951 = _32942 ^ _69950;
  wire _69952 = _27184 ^ _11266;
  wire _69953 = _69951 ^ _69952;
  wire _69954 = _69949 ^ _69953;
  wire _69955 = uncoded_block[1527] ^ uncoded_block[1540];
  wire _69956 = uncoded_block[1604] ^ uncoded_block[1663];
  wire _69957 = _69955 ^ _69956;
  wire _69958 = _64450 ^ _3190;
  wire _69959 = _69957 ^ _69958;
  wire _69960 = _69959 ^ uncoded_block[1710];
  wire _69961 = _69954 ^ _69960;
  wire _69962 = _69945 ^ _69961;
  wire _69963 = uncoded_block[2] ^ uncoded_block[27];
  wire _69964 = uncoded_block[30] ^ uncoded_block[69];
  wire _69965 = _69963 ^ _69964;
  wire _69966 = uncoded_block[72] ^ uncoded_block[84];
  wire _69967 = uncoded_block[118] ^ uncoded_block[161];
  wire _69968 = _69966 ^ _69967;
  wire _69969 = _69965 ^ _69968;
  wire _69970 = uncoded_block[185] ^ uncoded_block[203];
  wire _69971 = _61262 ^ _69970;
  wire _69972 = uncoded_block[226] ^ uncoded_block[257];
  wire _69973 = uncoded_block[273] ^ uncoded_block[288];
  wire _69974 = _69972 ^ _69973;
  wire _69975 = _69971 ^ _69974;
  wire _69976 = _69969 ^ _69975;
  wire _69977 = uncoded_block[335] ^ uncoded_block[357];
  wire _69978 = _37581 ^ _69977;
  wire _69979 = uncoded_block[388] ^ uncoded_block[435];
  wire _69980 = _69979 ^ _5580;
  wire _69981 = _69978 ^ _69980;
  wire _69982 = uncoded_block[481] ^ uncoded_block[512];
  wire _69983 = _1076 ^ _69982;
  wire _69984 = _67684 ^ _22936;
  wire _69985 = _69983 ^ _69984;
  wire _69986 = _69981 ^ _69985;
  wire _69987 = _69976 ^ _69986;
  wire _69988 = uncoded_block[597] ^ uncoded_block[618];
  wire _69989 = _69988 ^ _58805;
  wire _69990 = uncoded_block[670] ^ uncoded_block[676];
  wire _69991 = uncoded_block[707] ^ uncoded_block[741];
  wire _69992 = _69990 ^ _69991;
  wire _69993 = _69989 ^ _69992;
  wire _69994 = _59511 ^ _38464;
  wire _69995 = uncoded_block[815] ^ uncoded_block[832];
  wire _69996 = _69995 ^ _60675;
  wire _69997 = _69994 ^ _69996;
  wire _69998 = _69993 ^ _69997;
  wire _69999 = uncoded_block[908] ^ uncoded_block[951];
  wire _70000 = _69999 ^ _26197;
  wire _70001 = uncoded_block[1035] ^ uncoded_block[1065];
  wire _70002 = _484 ^ _70001;
  wire _70003 = _70000 ^ _70002;
  wire _70004 = uncoded_block[1083] ^ uncoded_block[1117];
  wire _70005 = uncoded_block[1141] ^ uncoded_block[1158];
  wire _70006 = _70004 ^ _70005;
  wire _70007 = uncoded_block[1194] ^ uncoded_block[1222];
  wire _70008 = _590 ^ _70007;
  wire _70009 = _70006 ^ _70008;
  wire _70010 = _70003 ^ _70009;
  wire _70011 = _69998 ^ _70010;
  wire _70012 = _69987 ^ _70011;
  wire _70013 = uncoded_block[1234] ^ uncoded_block[1290];
  wire _70014 = uncoded_block[1311] ^ uncoded_block[1324];
  wire _70015 = _70013 ^ _70014;
  wire _70016 = uncoded_block[1329] ^ uncoded_block[1345];
  wire _70017 = uncoded_block[1366] ^ uncoded_block[1382];
  wire _70018 = _70016 ^ _70017;
  wire _70019 = _70015 ^ _70018;
  wire _70020 = _27590 ^ _7842;
  wire _70021 = uncoded_block[1443] ^ uncoded_block[1456];
  wire _70022 = uncoded_block[1506] ^ uncoded_block[1524];
  wire _70023 = _70021 ^ _70022;
  wire _70024 = _70020 ^ _70023;
  wire _70025 = _70019 ^ _70024;
  wire _70026 = uncoded_block[1540] ^ uncoded_block[1595];
  wire _70027 = uncoded_block[1630] ^ uncoded_block[1657];
  wire _70028 = _70026 ^ _70027;
  wire _70029 = uncoded_block[1661] ^ uncoded_block[1667];
  wire _70030 = uncoded_block[1695] ^ uncoded_block[1702];
  wire _70031 = _70029 ^ _70030;
  wire _70032 = _70028 ^ _70031;
  wire _70033 = _70032 ^ uncoded_block[1709];
  wire _70034 = _70025 ^ _70033;
  wire _70035 = _70012 ^ _70034;
  wire _70036 = uncoded_block[4] ^ uncoded_block[31];
  wire _70037 = uncoded_block[48] ^ uncoded_block[68];
  wire _70038 = _70036 ^ _70037;
  wire _70039 = uncoded_block[119] ^ uncoded_block[185];
  wire _70040 = _26393 ^ _70039;
  wire _70041 = _70038 ^ _70040;
  wire _70042 = uncoded_block[242] ^ uncoded_block[264];
  wire _70043 = _60626 ^ _70042;
  wire _70044 = uncoded_block[274] ^ uncoded_block[284];
  wire _70045 = uncoded_block[289] ^ uncoded_block[315];
  wire _70046 = _70044 ^ _70045;
  wire _70047 = _70043 ^ _70046;
  wire _70048 = _70041 ^ _70047;
  wire _70049 = uncoded_block[336] ^ uncoded_block[372];
  wire _70050 = _70049 ^ _67795;
  wire _70051 = uncoded_block[433] ^ uncoded_block[445];
  wire _70052 = uncoded_block[456] ^ uncoded_block[473];
  wire _70053 = _70051 ^ _70052;
  wire _70054 = _70050 ^ _70053;
  wire _70055 = uncoded_block[476] ^ uncoded_block[518];
  wire _70056 = uncoded_block[537] ^ uncoded_block[553];
  wire _70057 = _70055 ^ _70056;
  wire _70058 = uncoded_block[564] ^ uncoded_block[581];
  wire _70059 = uncoded_block[583] ^ uncoded_block[652];
  wire _70060 = _70058 ^ _70059;
  wire _70061 = _70057 ^ _70060;
  wire _70062 = _70054 ^ _70061;
  wire _70063 = _70048 ^ _70062;
  wire _70064 = uncoded_block[688] ^ uncoded_block[704];
  wire _70065 = _4975 ^ _70064;
  wire _70066 = _62223 ^ _56505;
  wire _70067 = _70065 ^ _70066;
  wire _70068 = _49309 ^ _4331;
  wire _70069 = uncoded_block[864] ^ uncoded_block[909];
  wire _70070 = uncoded_block[920] ^ uncoded_block[940];
  wire _70071 = _70069 ^ _70070;
  wire _70072 = _70068 ^ _70071;
  wire _70073 = _70067 ^ _70072;
  wire _70074 = uncoded_block[969] ^ uncoded_block[979];
  wire _70075 = uncoded_block[992] ^ uncoded_block[1005];
  wire _70076 = _70074 ^ _70075;
  wire _70077 = uncoded_block[1012] ^ uncoded_block[1039];
  wire _70078 = uncoded_block[1097] ^ uncoded_block[1109];
  wire _70079 = _70077 ^ _70078;
  wire _70080 = _70076 ^ _70079;
  wire _70081 = uncoded_block[1118] ^ uncoded_block[1182];
  wire _70082 = _56844 ^ _70081;
  wire _70083 = uncoded_block[1186] ^ uncoded_block[1205];
  wire _70084 = _70083 ^ _56863;
  wire _70085 = _70082 ^ _70084;
  wire _70086 = _70080 ^ _70085;
  wire _70087 = _70073 ^ _70086;
  wire _70088 = _70063 ^ _70087;
  wire _70089 = uncoded_block[1289] ^ uncoded_block[1325];
  wire _70090 = _32082 ^ _70089;
  wire _70091 = uncoded_block[1357] ^ uncoded_block[1367];
  wire _70092 = uncoded_block[1380] ^ uncoded_block[1389];
  wire _70093 = _70091 ^ _70092;
  wire _70094 = _70090 ^ _70093;
  wire _70095 = uncoded_block[1398] ^ uncoded_block[1420];
  wire _70096 = uncoded_block[1423] ^ uncoded_block[1436];
  wire _70097 = _70095 ^ _70096;
  wire _70098 = uncoded_block[1444] ^ uncoded_block[1462];
  wire _70099 = uncoded_block[1469] ^ uncoded_block[1476];
  wire _70100 = _70098 ^ _70099;
  wire _70101 = _70097 ^ _70100;
  wire _70102 = _70094 ^ _70101;
  wire _70103 = uncoded_block[1512] ^ uncoded_block[1530];
  wire _70104 = uncoded_block[1554] ^ uncoded_block[1605];
  wire _70105 = _70103 ^ _70104;
  wire _70106 = uncoded_block[1617] ^ uncoded_block[1630];
  wire _70107 = uncoded_block[1639] ^ uncoded_block[1654];
  wire _70108 = _70106 ^ _70107;
  wire _70109 = _70105 ^ _70108;
  wire _70110 = _70109 ^ uncoded_block[1718];
  wire _70111 = _70102 ^ _70110;
  wire _70112 = _70088 ^ _70111;
  wire _70113 = uncoded_block[14] ^ uncoded_block[37];
  wire _70114 = uncoded_block[51] ^ uncoded_block[79];
  wire _70115 = _70113 ^ _70114;
  wire _70116 = _50014 ^ _59257;
  wire _70117 = _70115 ^ _70116;
  wire _70118 = uncoded_block[166] ^ uncoded_block[174];
  wire _70119 = uncoded_block[194] ^ uncoded_block[208];
  wire _70120 = _70118 ^ _70119;
  wire _70121 = _50418 ^ _66227;
  wire _70122 = _70120 ^ _70121;
  wire _70123 = _70117 ^ _70122;
  wire _70124 = uncoded_block[294] ^ uncoded_block[317];
  wire _70125 = _70124 ^ _6859;
  wire _70126 = uncoded_block[363] ^ uncoded_block[394];
  wire _70127 = uncoded_block[428] ^ uncoded_block[440];
  wire _70128 = _70126 ^ _70127;
  wire _70129 = _70125 ^ _70128;
  wire _70130 = uncoded_block[488] ^ uncoded_block[536];
  wire _70131 = _13662 ^ _70130;
  wire _70132 = uncoded_block[575] ^ uncoded_block[586];
  wire _70133 = _63063 ^ _70132;
  wire _70134 = _70131 ^ _70133;
  wire _70135 = _70129 ^ _70134;
  wire _70136 = _70123 ^ _70135;
  wire _70137 = uncoded_block[627] ^ uncoded_block[655];
  wire _70138 = _64807 ^ _70137;
  wire _70139 = uncoded_block[689] ^ uncoded_block[747];
  wire _70140 = _43772 ^ _70139;
  wire _70141 = _70138 ^ _70140;
  wire _70142 = _63462 ^ _63465;
  wire _70143 = uncoded_block[798] ^ uncoded_block[835];
  wire _70144 = _70143 ^ _2814;
  wire _70145 = _70142 ^ _70144;
  wire _70146 = _70141 ^ _70145;
  wire _70147 = uncoded_block[914] ^ uncoded_block[933];
  wire _70148 = uncoded_block[937] ^ uncoded_block[975];
  wire _70149 = _70147 ^ _70148;
  wire _70150 = uncoded_block[980] ^ uncoded_block[999];
  wire _70151 = _70150 ^ _42728;
  wire _70152 = _70149 ^ _70151;
  wire _70153 = uncoded_block[1046] ^ uncoded_block[1062];
  wire _70154 = uncoded_block[1068] ^ uncoded_block[1076];
  wire _70155 = _70153 ^ _70154;
  wire _70156 = uncoded_block[1108] ^ uncoded_block[1123];
  wire _70157 = _70156 ^ _2188;
  wire _70158 = _70155 ^ _70157;
  wire _70159 = _70152 ^ _70158;
  wire _70160 = _70146 ^ _70159;
  wire _70161 = _70136 ^ _70160;
  wire _70162 = uncoded_block[1168] ^ uncoded_block[1187];
  wire _70163 = uncoded_block[1213] ^ uncoded_block[1239];
  wire _70164 = _70162 ^ _70163;
  wire _70165 = uncoded_block[1240] ^ uncoded_block[1263];
  wire _70166 = _70165 ^ _17431;
  wire _70167 = _70164 ^ _70166;
  wire _70168 = uncoded_block[1354] ^ uncoded_block[1372];
  wire _70169 = _70168 ^ _63519;
  wire _70170 = uncoded_block[1449] ^ uncoded_block[1464];
  wire _70171 = _13951 ^ _70170;
  wire _70172 = _70169 ^ _70171;
  wire _70173 = _70167 ^ _70172;
  wire _70174 = _9042 ^ _36230;
  wire _70175 = uncoded_block[1534] ^ uncoded_block[1599];
  wire _70176 = uncoded_block[1625] ^ uncoded_block[1652];
  wire _70177 = _70175 ^ _70176;
  wire _70178 = _70174 ^ _70177;
  wire _70179 = uncoded_block[1690] ^ uncoded_block[1698];
  wire _70180 = _70179 ^ uncoded_block[1699];
  wire _70181 = _70178 ^ _70180;
  wire _70182 = _70173 ^ _70181;
  wire _70183 = _70161 ^ _70182;
  wire _70184 = uncoded_block[26] ^ uncoded_block[40];
  wire _70185 = _70184 ^ _28438;
  wire _70186 = uncoded_block[127] ^ uncoded_block[166];
  wire _70187 = uncoded_block[173] ^ uncoded_block[211];
  wire _70188 = _70186 ^ _70187;
  wire _70189 = _70185 ^ _70188;
  wire _70190 = uncoded_block[229] ^ uncoded_block[256];
  wire _70191 = uncoded_block[297] ^ uncoded_block[305];
  wire _70192 = _70190 ^ _70191;
  wire _70193 = uncoded_block[345] ^ uncoded_block[356];
  wire _70194 = uncoded_block[397] ^ uncoded_block[447];
  wire _70195 = _70193 ^ _70194;
  wire _70196 = _70192 ^ _70195;
  wire _70197 = _70189 ^ _70196;
  wire _70198 = uncoded_block[457] ^ uncoded_block[464];
  wire _70199 = uncoded_block[525] ^ uncoded_block[560];
  wire _70200 = _70198 ^ _70199;
  wire _70201 = uncoded_block[568] ^ uncoded_block[588];
  wire _70202 = _70201 ^ _3513;
  wire _70203 = _70200 ^ _70202;
  wire _70204 = _1180 ^ _49300;
  wire _70205 = uncoded_block[841] ^ uncoded_block[855];
  wire _70206 = _41210 ^ _70205;
  wire _70207 = _70204 ^ _70206;
  wire _70208 = _70203 ^ _70207;
  wire _70209 = _70197 ^ _70208;
  wire _70210 = uncoded_block[902] ^ uncoded_block[916];
  wire _70211 = uncoded_block[950] ^ uncoded_block[978];
  wire _70212 = _70210 ^ _70211;
  wire _70213 = uncoded_block[1004] ^ uncoded_block[1012];
  wire _70214 = uncoded_block[1065] ^ uncoded_block[1082];
  wire _70215 = _70213 ^ _70214;
  wire _70216 = _70212 ^ _70215;
  wire _70217 = uncoded_block[1126] ^ uncoded_block[1140];
  wire _70218 = uncoded_block[1179] ^ uncoded_block[1190];
  wire _70219 = _70217 ^ _70218;
  wire _70220 = uncoded_block[1233] ^ uncoded_block[1266];
  wire _70221 = uncoded_block[1282] ^ uncoded_block[1289];
  wire _70222 = _70220 ^ _70221;
  wire _70223 = _70219 ^ _70222;
  wire _70224 = _70216 ^ _70223;
  wire _70225 = uncoded_block[1420] ^ uncoded_block[1431];
  wire _70226 = _62771 ^ _70225;
  wire _70227 = uncoded_block[1451] ^ uncoded_block[1475];
  wire _70228 = uncoded_block[1486] ^ uncoded_block[1531];
  wire _70229 = _70227 ^ _70228;
  wire _70230 = _70226 ^ _70229;
  wire _70231 = uncoded_block[1539] ^ uncoded_block[1594];
  wire _70232 = _70231 ^ _61057;
  wire _70233 = _70232 ^ uncoded_block[1656];
  wire _70234 = _70230 ^ _70233;
  wire _70235 = _70224 ^ _70234;
  wire _70236 = _70209 ^ _70235;
  wire _70237 = uncoded_block[14] ^ uncoded_block[82];
  wire _70238 = uncoded_block[86] ^ uncoded_block[128];
  wire _70239 = _70237 ^ _70238;
  wire _70240 = uncoded_block[133] ^ uncoded_block[179];
  wire _70241 = uncoded_block[212] ^ uncoded_block[230];
  wire _70242 = _70240 ^ _70241;
  wire _70243 = _70239 ^ _70242;
  wire _70244 = uncoded_block[267] ^ uncoded_block[298];
  wire _70245 = uncoded_block[317] ^ uncoded_block[346];
  wire _70246 = _70244 ^ _70245;
  wire _70247 = uncoded_block[398] ^ uncoded_block[464];
  wire _70248 = _56452 ^ _70247;
  wire _70249 = _70246 ^ _70248;
  wire _70250 = _70243 ^ _70249;
  wire _70251 = uncoded_block[465] ^ uncoded_block[506];
  wire _70252 = uncoded_block[530] ^ uncoded_block[589];
  wire _70253 = _70251 ^ _70252;
  wire _70254 = uncoded_block[605] ^ uncoded_block[640];
  wire _70255 = uncoded_block[659] ^ uncoded_block[678];
  wire _70256 = _70254 ^ _70255;
  wire _70257 = _70253 ^ _70256;
  wire _70258 = uncoded_block[787] ^ uncoded_block[811];
  wire _70259 = _67506 ^ _70258;
  wire _70260 = uncoded_block[832] ^ uncoded_block[842];
  wire _70261 = uncoded_block[917] ^ uncoded_block[939];
  wire _70262 = _70260 ^ _70261;
  wire _70263 = _70259 ^ _70262;
  wire _70264 = _70257 ^ _70263;
  wire _70265 = _70250 ^ _70264;
  wire _70266 = uncoded_block[1013] ^ uncoded_block[1043];
  wire _70267 = _62404 ^ _70266;
  wire _70268 = uncoded_block[1066] ^ uncoded_block[1080];
  wire _70269 = uncoded_block[1127] ^ uncoded_block[1149];
  wire _70270 = _70268 ^ _70269;
  wire _70271 = _70267 ^ _70270;
  wire _70272 = uncoded_block[1191] ^ uncoded_block[1204];
  wire _70273 = _70272 ^ _24018;
  wire _70274 = uncoded_block[1283] ^ uncoded_block[1312];
  wire _70275 = uncoded_block[1376] ^ uncoded_block[1432];
  wire _70276 = _70274 ^ _70275;
  wire _70277 = _70273 ^ _70276;
  wire _70278 = _70271 ^ _70277;
  wire _70279 = _1544 ^ _57765;
  wire _70280 = uncoded_block[1533] ^ uncoded_block[1576];
  wire _70281 = _21338 ^ _70280;
  wire _70282 = _70279 ^ _70281;
  wire _70283 = uncoded_block[1638] ^ uncoded_block[1663];
  wire _70284 = _70283 ^ _62447;
  wire _70285 = _70284 ^ uncoded_block[1714];
  wire _70286 = _70282 ^ _70285;
  wire _70287 = _70278 ^ _70286;
  wire _70288 = _70265 ^ _70287;
  wire _70289 = uncoded_block[87] ^ uncoded_block[111];
  wire _70290 = uncoded_block[198] ^ uncoded_block[237];
  wire _70291 = _70289 ^ _70290;
  wire _70292 = uncoded_block[323] ^ uncoded_block[371];
  wire _70293 = uncoded_block[437] ^ uncoded_block[471];
  wire _70294 = _70292 ^ _70293;
  wire _70295 = _70291 ^ _70294;
  wire _70296 = uncoded_block[547] ^ uncoded_block[603];
  wire _70297 = _70296 ^ _65565;
  wire _70298 = uncoded_block[851] ^ uncoded_block[894];
  wire _70299 = _65569 ^ _70298;
  wire _70300 = _70297 ^ _70299;
  wire _70301 = _70295 ^ _70300;
  wire _70302 = uncoded_block[958] ^ uncoded_block[1033];
  wire _70303 = uncoded_block[1091] ^ uncoded_block[1124];
  wire _70304 = _70302 ^ _70303;
  wire _70305 = uncoded_block[1178] ^ uncoded_block[1260];
  wire _70306 = uncoded_block[1324] ^ uncoded_block[1331];
  wire _70307 = _70305 ^ _70306;
  wire _70308 = _70304 ^ _70307;
  wire _70309 = uncoded_block[1376] ^ uncoded_block[1396];
  wire _70310 = uncoded_block[1562] ^ uncoded_block[1588];
  wire _70311 = _70309 ^ _70310;
  wire _70312 = uncoded_block[1628] ^ uncoded_block[1708];
  wire _70313 = _70312 ^ uncoded_block[1720];
  wire _70314 = _70311 ^ _70313;
  wire _70315 = _70308 ^ _70314;
  wire _70316 = _70301 ^ _70315;
  wire _70317 = uncoded_block[77] ^ uncoded_block[118];
  wire _70318 = uncoded_block[182] ^ uncoded_block[270];
  wire _70319 = _70317 ^ _70318;
  wire _70320 = uncoded_block[317] ^ uncoded_block[356];
  wire _70321 = uncoded_block[398] ^ uncoded_block[498];
  wire _70322 = _70320 ^ _70321;
  wire _70323 = _70319 ^ _70322;
  wire _70324 = uncoded_block[512] ^ uncoded_block[574];
  wire _70325 = uncoded_block[650] ^ uncoded_block[677];
  wire _70326 = _70324 ^ _70325;
  wire _70327 = uncoded_block[742] ^ uncoded_block[801];
  wire _70328 = uncoded_block[852] ^ uncoded_block[923];
  wire _70329 = _70327 ^ _70328;
  wire _70330 = _70326 ^ _70329;
  wire _70331 = _70323 ^ _70330;
  wire _70332 = uncoded_block[976] ^ uncoded_block[1036];
  wire _70333 = uncoded_block[1171] ^ uncoded_block[1248];
  wire _70334 = _70332 ^ _70333;
  wire _70335 = uncoded_block[1316] ^ uncoded_block[1358];
  wire _70336 = uncoded_block[1403] ^ uncoded_block[1446];
  wire _70337 = _70335 ^ _70336;
  wire _70338 = _70334 ^ _70337;
  wire _70339 = uncoded_block[1559] ^ uncoded_block[1587];
  wire _70340 = _23624 ^ _70339;
  wire _70341 = uncoded_block[1674] ^ uncoded_block[1713];
  wire _70342 = _70341 ^ uncoded_block[1721];
  wire _70343 = _70340 ^ _70342;
  wire _70344 = _70338 ^ _70343;
  wire _70345 = _70331 ^ _70344;
  wire _70346 = uncoded_block[14] ^ uncoded_block[91];
  wire _70347 = uncoded_block[116] ^ uncoded_block[174];
  wire _70348 = _70346 ^ _70347;
  wire _70349 = uncoded_block[345] ^ uncoded_block[440];
  wire _70350 = _66227 ^ _70349;
  wire _70351 = _70348 ^ _70350;
  wire _70352 = uncoded_block[488] ^ uncoded_block[537];
  wire _70353 = uncoded_block[575] ^ uncoded_block[627];
  wire _70354 = _70352 ^ _70353;
  wire _70355 = uncoded_block[689] ^ uncoded_block[767];
  wire _70356 = uncoded_block[779] ^ uncoded_block[836];
  wire _70357 = _70355 ^ _70356;
  wire _70358 = _70354 ^ _70357;
  wire _70359 = _70351 ^ _70358;
  wire _70360 = uncoded_block[937] ^ uncoded_block[980];
  wire _70361 = _70360 ^ _68017;
  wire _70362 = uncoded_block[1239] ^ uncoded_block[1298];
  wire _70363 = _66256 ^ _70362;
  wire _70364 = _70361 ^ _70363;
  wire _70365 = uncoded_block[1414] ^ uncoded_block[1438];
  wire _70366 = _70365 ^ _64607;
  wire _70367 = _66271 ^ uncoded_block[1698];
  wire _70368 = _70366 ^ _70367;
  wire _70369 = _70364 ^ _70368;
  wire _70370 = _70359 ^ _70369;
  wire _70371 = uncoded_block[27] ^ uncoded_block[73];
  wire _70372 = uncoded_block[124] ^ uncoded_block[199];
  wire _70373 = _70371 ^ _70372;
  wire _70374 = uncoded_block[225] ^ uncoded_block[328];
  wire _70375 = uncoded_block[337] ^ uncoded_block[412];
  wire _70376 = _70374 ^ _70375;
  wire _70377 = _70373 ^ _70376;
  wire _70378 = uncoded_block[572] ^ uncoded_block[625];
  wire _70379 = _69913 ^ _70378;
  wire _70380 = uncoded_block[680] ^ uncoded_block[745];
  wire _70381 = uncoded_block[796] ^ uncoded_block[858];
  wire _70382 = _70380 ^ _70381;
  wire _70383 = _70379 ^ _70382;
  wire _70384 = _70377 ^ _70383;
  wire _70385 = uncoded_block[939] ^ uncoded_block[959];
  wire _70386 = _70385 ^ _66671;
  wire _70387 = uncoded_block[1121] ^ uncoded_block[1202];
  wire _70388 = uncoded_block[1264] ^ uncoded_block[1297];
  wire _70389 = _70387 ^ _70388;
  wire _70390 = _70386 ^ _70389;
  wire _70391 = uncoded_block[1330] ^ uncoded_block[1360];
  wire _70392 = uncoded_block[1387] ^ uncoded_block[1540];
  wire _70393 = _70391 ^ _70392;
  wire _70394 = uncoded_block[1604] ^ uncoded_block[1666];
  wire _70395 = _70394 ^ uncoded_block[1710];
  wire _70396 = _70393 ^ _70395;
  wire _70397 = _70390 ^ _70396;
  wire _70398 = _70384 ^ _70397;
  wire _70399 = uncoded_block[143] ^ uncoded_block[218];
  wire _70400 = _69261 ^ _70399;
  wire _70401 = uncoded_block[238] ^ uncoded_block[307];
  wire _70402 = uncoded_block[367] ^ uncoded_block[443];
  wire _70403 = _70401 ^ _70402;
  wire _70404 = _70400 ^ _70403;
  wire _70405 = uncoded_block[449] ^ uncoded_block[514];
  wire _70406 = uncoded_block[613] ^ uncoded_block[659];
  wire _70407 = _70405 ^ _70406;
  wire _70408 = uncoded_block[673] ^ uncoded_block[763];
  wire _70409 = uncoded_block[805] ^ uncoded_block[850];
  wire _70410 = _70408 ^ _70409;
  wire _70411 = _70407 ^ _70410;
  wire _70412 = _70404 ^ _70411;
  wire _70413 = uncoded_block[938] ^ uncoded_block[971];
  wire _70414 = uncoded_block[1053] ^ uncoded_block[1094];
  wire _70415 = _70413 ^ _70414;
  wire _70416 = uncoded_block[1129] ^ uncoded_block[1207];
  wire _70417 = uncoded_block[1272] ^ uncoded_block[1293];
  wire _70418 = _70416 ^ _70417;
  wire _70419 = _70415 ^ _70418;
  wire _70420 = uncoded_block[1351] ^ uncoded_block[1400];
  wire _70421 = _70420 ^ _66402;
  wire _70422 = uncoded_block[1470] ^ uncoded_block[1621];
  wire _70423 = _70422 ^ uncoded_block[1675];
  wire _70424 = _70421 ^ _70423;
  wire _70425 = _70419 ^ _70424;
  wire _70426 = _70412 ^ _70425;
  wire _70427 = uncoded_block[35] ^ uncoded_block[96];
  wire _70428 = uncoded_block[163] ^ uncoded_block[216];
  wire _70429 = _70427 ^ _70428;
  wire _70430 = uncoded_block[247] ^ uncoded_block[322];
  wire _70431 = uncoded_block[389] ^ uncoded_block[426];
  wire _70432 = _70430 ^ _70431;
  wire _70433 = _70429 ^ _70432;
  wire _70434 = uncoded_block[459] ^ uncoded_block[550];
  wire _70435 = uncoded_block[600] ^ uncoded_block[660];
  wire _70436 = _70434 ^ _70435;
  wire _70437 = uncoded_block[718] ^ uncoded_block[738];
  wire _70438 = uncoded_block[791] ^ uncoded_block[873];
  wire _70439 = _70437 ^ _70438;
  wire _70440 = _70436 ^ _70439;
  wire _70441 = _70433 ^ _70440;
  wire _70442 = uncoded_block[898] ^ uncoded_block[1002];
  wire _70443 = uncoded_block[1032] ^ uncoded_block[1100];
  wire _70444 = _70442 ^ _70443;
  wire _70445 = _66882 ^ _65227;
  wire _70446 = _70444 ^ _70445;
  wire _70447 = uncoded_block[1299] ^ uncoded_block[1368];
  wire _70448 = uncoded_block[1397] ^ uncoded_block[1563];
  wire _70449 = _70447 ^ _70448;
  wire _70450 = _66897 ^ uncoded_block[1649];
  wire _70451 = _70449 ^ _70450;
  wire _70452 = _70446 ^ _70451;
  wire _70453 = _70441 ^ _70452;
  wire _70454 = uncoded_block[44] ^ uncoded_block[97];
  wire _70455 = uncoded_block[131] ^ uncoded_block[212];
  wire _70456 = _70454 ^ _70455;
  wire _70457 = uncoded_block[255] ^ uncoded_block[280];
  wire _70458 = uncoded_block[348] ^ uncoded_block[420];
  wire _70459 = _70457 ^ _70458;
  wire _70460 = _70456 ^ _70459;
  wire _70461 = uncoded_block[494] ^ uncoded_block[516];
  wire _70462 = uncoded_block[599] ^ uncoded_block[665];
  wire _70463 = _70461 ^ _70462;
  wire _70464 = uncoded_block[671] ^ uncoded_block[760];
  wire _70465 = uncoded_block[782] ^ uncoded_block[833];
  wire _70466 = _70464 ^ _70465;
  wire _70467 = _70463 ^ _70466;
  wire _70468 = _70460 ^ _70467;
  wire _70469 = uncoded_block[907] ^ uncoded_block[947];
  wire _70470 = uncoded_block[1047] ^ uncoded_block[1065];
  wire _70471 = _70469 ^ _70470;
  wire _70472 = uncoded_block[1148] ^ uncoded_block[1268];
  wire _70473 = uncoded_block[1278] ^ uncoded_block[1361];
  wire _70474 = _70472 ^ _70473;
  wire _70475 = _70471 ^ _70474;
  wire _70476 = uncoded_block[1607] ^ uncoded_block[1626];
  wire _70477 = _70476 ^ uncoded_block[1667];
  wire _70478 = _67959 ^ _70477;
  wire _70479 = _70475 ^ _70478;
  wire _70480 = _70468 ^ _70479;
  wire _70481 = uncoded_block[137] ^ uncoded_block[185];
  wire _70482 = _67781 ^ _70481;
  wire _70483 = uncoded_block[242] ^ uncoded_block[284];
  wire _70484 = _70483 ^ _67795;
  wire _70485 = _70482 ^ _70484;
  wire _70486 = uncoded_block[583] ^ uncoded_block[653];
  wire _70487 = _70055 ^ _70486;
  wire _70488 = uncoded_block[704] ^ uncoded_block[753];
  wire _70489 = uncoded_block[784] ^ uncoded_block[832];
  wire _70490 = _70488 ^ _70489;
  wire _70491 = _70487 ^ _70490;
  wire _70492 = _70485 ^ _70491;
  wire _70493 = uncoded_block[940] ^ uncoded_block[979];
  wire _70494 = uncoded_block[1012] ^ uncoded_block[1097];
  wire _70495 = _70493 ^ _70494;
  wire _70496 = uncoded_block[1186] ^ uncoded_block[1227];
  wire _70497 = uncoded_block[1289] ^ uncoded_block[1357];
  wire _70498 = _70496 ^ _70497;
  wire _70499 = _70495 ^ _70498;
  wire _70500 = uncoded_block[1462] ^ uncoded_block[1512];
  wire _70501 = _66202 ^ _70500;
  wire _70502 = uncoded_block[1554] ^ uncoded_block[1617];
  wire _70503 = _70502 ^ uncoded_block[1718];
  wire _70504 = _70501 ^ _70503;
  wire _70505 = _70499 ^ _70504;
  wire _70506 = _70492 ^ _70505;
  wire _70507 = uncoded_block[49] ^ uncoded_block[109];
  wire _70508 = uncoded_block[113] ^ uncoded_block[223];
  wire _70509 = _70507 ^ _70508;
  wire _70510 = uncoded_block[273] ^ uncoded_block[302];
  wire _70511 = uncoded_block[369] ^ uncoded_block[400];
  wire _70512 = _70510 ^ _70511;
  wire _70513 = _70509 ^ _70512;
  wire _70514 = uncoded_block[490] ^ uncoded_block[544];
  wire _70515 = uncoded_block[593] ^ uncoded_block[640];
  wire _70516 = _70514 ^ _70515;
  wire _70517 = uncoded_block[693] ^ uncoded_block[821];
  wire _70518 = uncoded_block[855] ^ uncoded_block[936];
  wire _70519 = _70517 ^ _70518;
  wire _70520 = _70516 ^ _70519;
  wire _70521 = _70513 ^ _70520;
  wire _70522 = uncoded_block[951] ^ uncoded_block[1050];
  wire _70523 = _70522 ^ _66948;
  wire _70524 = uncoded_block[1169] ^ uncoded_block[1206];
  wire _70525 = uncoded_block[1237] ^ uncoded_block[1288];
  wire _70526 = _70524 ^ _70525;
  wire _70527 = _70523 ^ _70526;
  wire _70528 = uncoded_block[1369] ^ uncoded_block[1411];
  wire _70529 = uncoded_block[1427] ^ uncoded_block[1499];
  wire _70530 = _70528 ^ _70529;
  wire _70531 = uncoded_block[1614] ^ uncoded_block[1653];
  wire _70532 = _70531 ^ uncoded_block[1704];
  wire _70533 = _70530 ^ _70532;
  wire _70534 = _70527 ^ _70533;
  wire _70535 = _70521 ^ _70534;
  wire _70536 = uncoded_block[52] ^ uncoded_block[66];
  wire _70537 = uncoded_block[151] ^ uncoded_block[221];
  wire _70538 = _70536 ^ _70537;
  wire _70539 = uncoded_block[237] ^ uncoded_block[289];
  wire _70540 = uncoded_block[361] ^ uncoded_block[411];
  wire _70541 = _70539 ^ _70540;
  wire _70542 = _70538 ^ _70541;
  wire _70543 = uncoded_block[473] ^ uncoded_block[539];
  wire _70544 = uncoded_block[585] ^ uncoded_block[631];
  wire _70545 = _70543 ^ _70544;
  wire _70546 = uncoded_block[711] ^ uncoded_block[734];
  wire _70547 = uncoded_block[797] ^ uncoded_block[883];
  wire _70548 = _70546 ^ _70547;
  wire _70549 = _70545 ^ _70548;
  wire _70550 = _70542 ^ _70549;
  wire _70551 = uncoded_block[904] ^ uncoded_block[978];
  wire _70552 = uncoded_block[1046] ^ uncoded_block[1106];
  wire _70553 = _70551 ^ _70552;
  wire _70554 = uncoded_block[1130] ^ uncoded_block[1231];
  wire _70555 = uncoded_block[1305] ^ uncoded_block[1368];
  wire _70556 = _70554 ^ _70555;
  wire _70557 = _70553 ^ _70556;
  wire _70558 = uncoded_block[1416] ^ uncoded_block[1475];
  wire _70559 = uncoded_block[1485] ^ uncoded_block[1515];
  wire _70560 = _70558 ^ _70559;
  wire _70561 = uncoded_block[1595] ^ uncoded_block[1661];
  wire _70562 = _70561 ^ uncoded_block[1695];
  wire _70563 = _70560 ^ _70562;
  wire _70564 = _70557 ^ _70563;
  wire _70565 = _70550 ^ _70564;
  wire _70566 = uncoded_block[78] ^ uncoded_block[119];
  wire _70567 = uncoded_block[183] ^ uncoded_block[271];
  wire _70568 = _70566 ^ _70567;
  wire _70569 = uncoded_block[318] ^ uncoded_block[357];
  wire _70570 = uncoded_block[399] ^ uncoded_block[499];
  wire _70571 = _70569 ^ _70570;
  wire _70572 = _70568 ^ _70571;
  wire _70573 = uncoded_block[513] ^ uncoded_block[575];
  wire _70574 = uncoded_block[651] ^ uncoded_block[678];
  wire _70575 = _70573 ^ _70574;
  wire _70576 = uncoded_block[743] ^ uncoded_block[802];
  wire _70577 = uncoded_block[853] ^ uncoded_block[924];
  wire _70578 = _70576 ^ _70577;
  wire _70579 = _70575 ^ _70578;
  wire _70580 = _70572 ^ _70579;
  wire _70581 = uncoded_block[977] ^ uncoded_block[1037];
  wire _70582 = uncoded_block[1111] ^ uncoded_block[1172];
  wire _70583 = _70581 ^ _70582;
  wire _70584 = uncoded_block[1249] ^ uncoded_block[1317];
  wire _70585 = uncoded_block[1359] ^ uncoded_block[1404];
  wire _70586 = _70584 ^ _70585;
  wire _70587 = _70583 ^ _70586;
  wire _70588 = uncoded_block[1488] ^ uncoded_block[1511];
  wire _70589 = _61042 ^ _70588;
  wire _70590 = uncoded_block[1675] ^ uncoded_block[1714];
  wire _70591 = _70590 ^ uncoded_block[1722];
  wire _70592 = _70589 ^ _70591;
  wire _70593 = _70587 ^ _70592;
  wire _70594 = _70580 ^ _70593;
  wire _70595 = uncoded_block[6] ^ uncoded_block[80];
  wire _70596 = uncoded_block[115] ^ uncoded_block[209];
  wire _70597 = _70595 ^ _70596;
  wire _70598 = uncoded_block[276] ^ uncoded_block[323];
  wire _70599 = uncoded_block[342] ^ uncoded_block[443];
  wire _70600 = _70598 ^ _70599;
  wire _70601 = _70597 ^ _70600;
  wire _70602 = uncoded_block[501] ^ uncoded_block[533];
  wire _70603 = uncoded_block[588] ^ uncoded_block[636];
  wire _70604 = _70602 ^ _70603;
  wire _70605 = uncoded_block[707] ^ uncoded_block[733];
  wire _70606 = uncoded_block[813] ^ uncoded_block[844];
  wire _70607 = _70605 ^ _70606;
  wire _70608 = _70604 ^ _70607;
  wire _70609 = _70601 ^ _70608;
  wire _70610 = uncoded_block[906] ^ uncoded_block[974];
  wire _70611 = uncoded_block[1104] ^ uncoded_block[1112];
  wire _70612 = _70610 ^ _70611;
  wire _70613 = uncoded_block[1133] ^ uncoded_block[1170];
  wire _70614 = uncoded_block[1258] ^ uncoded_block[1292];
  wire _70615 = _70613 ^ _70614;
  wire _70616 = _70612 ^ _70615;
  wire _70617 = uncoded_block[1338] ^ uncoded_block[1436];
  wire _70618 = uncoded_block[1505] ^ uncoded_block[1604];
  wire _70619 = _70617 ^ _70618;
  wire _70620 = uncoded_block[1626] ^ uncoded_block[1685];
  wire _70621 = _70620 ^ uncoded_block[1702];
  wire _70622 = _70619 ^ _70621;
  wire _70623 = _70616 ^ _70622;
  wire _70624 = _70609 ^ _70623;
  wire _70625 = uncoded_block[16] ^ uncoded_block[73];
  wire _70626 = uncoded_block[123] ^ uncoded_block[196];
  wire _70627 = _70625 ^ _70626;
  wire _70628 = uncoded_block[258] ^ uncoded_block[284];
  wire _70629 = uncoded_block[373] ^ uncoded_block[400];
  wire _70630 = _70628 ^ _70629;
  wire _70631 = _70627 ^ _70630;
  wire _70632 = uncoded_block[465] ^ uncoded_block[537];
  wire _70633 = uncoded_block[609] ^ uncoded_block[632];
  wire _70634 = _70632 ^ _70633;
  wire _70635 = uncoded_block[713] ^ uncoded_block[748];
  wire _70636 = uncoded_block[791] ^ uncoded_block[831];
  wire _70637 = _70635 ^ _70636;
  wire _70638 = _70634 ^ _70637;
  wire _70639 = _70631 ^ _70638;
  wire _70640 = uncoded_block[922] ^ uncoded_block[965];
  wire _70641 = uncoded_block[1024] ^ uncoded_block[1094];
  wire _70642 = _70640 ^ _70641;
  wire _70643 = uncoded_block[1138] ^ uncoded_block[1217];
  wire _70644 = uncoded_block[1235] ^ uncoded_block[1287];
  wire _70645 = _70643 ^ _70644;
  wire _70646 = _70642 ^ _70645;
  wire _70647 = uncoded_block[1353] ^ uncoded_block[1393];
  wire _70648 = _70647 ^ _63966;
  wire _70649 = uncoded_block[1624] ^ uncoded_block[1686];
  wire _70650 = _70649 ^ uncoded_block[1689];
  wire _70651 = _70648 ^ _70650;
  wire _70652 = _70646 ^ _70651;
  wire _70653 = _70639 ^ _70652;
  wire _70654 = uncoded_block[17] ^ uncoded_block[77];
  wire _70655 = uncoded_block[113] ^ uncoded_block[197];
  wire _70656 = _70654 ^ _70655;
  wire _70657 = uncoded_block[306] ^ uncoded_block[354];
  wire _70658 = uncoded_block[397] ^ uncoded_block[479];
  wire _70659 = _70657 ^ _70658;
  wire _70660 = _70656 ^ _70659;
  wire _70661 = uncoded_block[516] ^ uncoded_block[579];
  wire _70662 = uncoded_block[668] ^ uncoded_block[712];
  wire _70663 = _70661 ^ _70662;
  wire _70664 = uncoded_block[732] ^ uncoded_block[818];
  wire _70665 = uncoded_block[864] ^ uncoded_block[930];
  wire _70666 = _70664 ^ _70665;
  wire _70667 = _70663 ^ _70666;
  wire _70668 = _70660 ^ _70667;
  wire _70669 = uncoded_block[993] ^ uncoded_block[1045];
  wire _70670 = uncoded_block[1085] ^ uncoded_block[1119];
  wire _70671 = _70669 ^ _70670;
  wire _70672 = uncoded_block[1214] ^ uncoded_block[1274];
  wire _70673 = uncoded_block[1302] ^ uncoded_block[1379];
  wire _70674 = _70672 ^ _70673;
  wire _70675 = _70671 ^ _70674;
  wire _70676 = uncoded_block[1448] ^ uncoded_block[1548];
  wire _70677 = uncoded_block[1567] ^ uncoded_block[1582];
  wire _70678 = _70676 ^ _70677;
  wire _70679 = uncoded_block[1636] ^ uncoded_block[1662];
  wire _70680 = _70679 ^ uncoded_block[1696];
  wire _70681 = _70678 ^ _70680;
  wire _70682 = _70675 ^ _70681;
  wire _70683 = _70668 ^ _70682;
  wire _70684 = uncoded_block[18] ^ uncoded_block[62];
  wire _70685 = uncoded_block[139] ^ uncoded_block[177];
  wire _70686 = _70684 ^ _70685;
  wire _70687 = uncoded_block[257] ^ uncoded_block[313];
  wire _70688 = uncoded_block[367] ^ uncoded_block[416];
  wire _70689 = _70687 ^ _70688;
  wire _70690 = _70686 ^ _70689;
  wire _70691 = uncoded_block[453] ^ uncoded_block[554];
  wire _70692 = uncoded_block[592] ^ uncoded_block[633];
  wire _70693 = _70691 ^ _70692;
  wire _70694 = uncoded_block[690] ^ uncoded_block[745];
  wire _70695 = uncoded_block[806] ^ uncoded_block[873];
  wire _70696 = _70694 ^ _70695;
  wire _70697 = _70693 ^ _70696;
  wire _70698 = _70690 ^ _70697;
  wire _70699 = uncoded_block[897] ^ uncoded_block[985];
  wire _70700 = uncoded_block[1017] ^ uncoded_block[1074];
  wire _70701 = _70699 ^ _70700;
  wire _70702 = uncoded_block[1122] ^ uncoded_block[1197];
  wire _70703 = uncoded_block[1226] ^ uncoded_block[1321];
  wire _70704 = _70702 ^ _70703;
  wire _70705 = _70701 ^ _70704;
  wire _70706 = uncoded_block[1365] ^ uncoded_block[1403];
  wire _70707 = uncoded_block[1575] ^ uncoded_block[1594];
  wire _70708 = _70706 ^ _70707;
  wire _70709 = uncoded_block[1630] ^ uncoded_block[1663];
  wire _70710 = _70709 ^ uncoded_block[1705];
  wire _70711 = _70708 ^ _70710;
  wire _70712 = _70705 ^ _70711;
  wire _70713 = _70698 ^ _70712;
  wire _70714 = uncoded_block[22] ^ uncoded_block[75];
  wire _70715 = uncoded_block[161] ^ uncoded_block[224];
  wire _70716 = _70714 ^ _70715;
  wire _70717 = uncoded_block[228] ^ uncoded_block[308];
  wire _70718 = uncoded_block[337] ^ uncoded_block[410];
  wire _70719 = _70717 ^ _70718;
  wire _70720 = _70716 ^ _70719;
  wire _70721 = uncoded_block[468] ^ uncoded_block[542];
  wire _70722 = uncoded_block[578] ^ uncoded_block[644];
  wire _70723 = _70721 ^ _70722;
  wire _70724 = uncoded_block[695] ^ uncoded_block[763];
  wire _70725 = uncoded_block[787] ^ uncoded_block[845];
  wire _70726 = _70724 ^ _70725;
  wire _70727 = _70723 ^ _70726;
  wire _70728 = _70720 ^ _70727;
  wire _70729 = uncoded_block[916] ^ uncoded_block[964];
  wire _70730 = uncoded_block[1010] ^ uncoded_block[1061];
  wire _70731 = _70729 ^ _70730;
  wire _70732 = uncoded_block[1135] ^ uncoded_block[1168];
  wire _70733 = uncoded_block[1206] ^ uncoded_block[1263];
  wire _70734 = _70732 ^ _70733;
  wire _70735 = _70731 ^ _70734;
  wire _70736 = uncoded_block[1324] ^ uncoded_block[1405];
  wire _70737 = uncoded_block[1473] ^ uncoded_block[1487];
  wire _70738 = _70736 ^ _70737;
  wire _70739 = _68178 ^ uncoded_block[1713];
  wire _70740 = _70738 ^ _70739;
  wire _70741 = _70735 ^ _70740;
  wire _70742 = _70728 ^ _70741;
  wire _70743 = uncoded_block[23] ^ uncoded_block[101];
  wire _70744 = uncoded_block[142] ^ uncoded_block[193];
  wire _70745 = _70743 ^ _70744;
  wire _70746 = uncoded_block[240] ^ uncoded_block[322];
  wire _70747 = uncoded_block[375] ^ uncoded_block[429];
  wire _70748 = _70746 ^ _70747;
  wire _70749 = _70745 ^ _70748;
  wire _70750 = uncoded_block[610] ^ uncoded_block[643];
  wire _70751 = _67493 ^ _70750;
  wire _70752 = uncoded_block[724] ^ uncoded_block[784];
  wire _70753 = _67503 ^ _70752;
  wire _70754 = _70751 ^ _70753;
  wire _70755 = _70749 ^ _70754;
  wire _70756 = uncoded_block[884] ^ uncoded_block[903];
  wire _70757 = uncoded_block[981] ^ uncoded_block[1028];
  wire _70758 = _70756 ^ _70757;
  wire _70759 = uncoded_block[1068] ^ uncoded_block[1121];
  wire _70760 = uncoded_block[1188] ^ uncoded_block[1267];
  wire _70761 = _70759 ^ _70760;
  wire _70762 = _70758 ^ _70761;
  wire _70763 = uncoded_block[1366] ^ uncoded_block[1476];
  wire _70764 = _66457 ^ _70763;
  wire _70765 = uncoded_block[1551] ^ uncoded_block[1611];
  wire _70766 = _70765 ^ uncoded_block[1687];
  wire _70767 = _70764 ^ _70766;
  wire _70768 = _70762 ^ _70767;
  wire _70769 = _70755 ^ _70768;
  wire _70770 = uncoded_block[26] ^ uncoded_block[100];
  wire _70771 = uncoded_block[137] ^ uncoded_block[181];
  wire _70772 = _70770 ^ _70771;
  wire _70773 = uncoded_block[245] ^ uncoded_block[320];
  wire _70774 = uncoded_block[353] ^ uncoded_block[436];
  wire _70775 = _70773 ^ _70774;
  wire _70776 = _70772 ^ _70775;
  wire _70777 = uncoded_block[572] ^ uncoded_block[662];
  wire _70778 = _68201 ^ _70777;
  wire _70779 = uncoded_block[803] ^ uncoded_block[881];
  wire _70780 = _68208 ^ _70779;
  wire _70781 = _70778 ^ _70780;
  wire _70782 = _70776 ^ _70781;
  wire _70783 = uncoded_block[928] ^ uncoded_block[961];
  wire _70784 = uncoded_block[1018] ^ uncoded_block[1088];
  wire _70785 = _70783 ^ _70784;
  wire _70786 = uncoded_block[1128] ^ uncoded_block[1164];
  wire _70787 = _70786 ^ _68227;
  wire _70788 = _70785 ^ _70787;
  wire _70789 = uncoded_block[1291] ^ uncoded_block[1374];
  wire _70790 = uncoded_block[1418] ^ uncoded_block[1432];
  wire _70791 = _70789 ^ _70790;
  wire _70792 = uncoded_block[1583] ^ uncoded_block[1640];
  wire _70793 = _70792 ^ uncoded_block[1684];
  wire _70794 = _70791 ^ _70793;
  wire _70795 = _70788 ^ _70794;
  wire _70796 = _70782 ^ _70795;
  wire _70797 = uncoded_block[29] ^ uncoded_block[90];
  wire _70798 = uncoded_block[163] ^ uncoded_block[182];
  wire _70799 = _70797 ^ _70798;
  wire _70800 = uncoded_block[236] ^ uncoded_block[298];
  wire _70801 = uncoded_block[340] ^ uncoded_block[422];
  wire _70802 = _70800 ^ _70801;
  wire _70803 = _70799 ^ _70802;
  wire _70804 = uncoded_block[449] ^ uncoded_block[557];
  wire _70805 = uncoded_block[569] ^ uncoded_block[648];
  wire _70806 = _70804 ^ _70805;
  wire _70807 = uncoded_block[700] ^ uncoded_block[771];
  wire _70808 = uncoded_block[799] ^ uncoded_block[875];
  wire _70809 = _70807 ^ _70808;
  wire _70810 = _70806 ^ _70809;
  wire _70811 = _70803 ^ _70810;
  wire _70812 = uncoded_block[931] ^ uncoded_block[950];
  wire _70813 = _70812 ^ _30731;
  wire _70814 = uncoded_block[1099] ^ uncoded_block[1120];
  wire _70815 = uncoded_block[1190] ^ uncoded_block[1237];
  wire _70816 = _70814 ^ _70815;
  wire _70817 = _70813 ^ _70816;
  wire _70818 = uncoded_block[1308] ^ uncoded_block[1356];
  wire _70819 = uncoded_block[1545] ^ uncoded_block[1560];
  wire _70820 = _70818 ^ _70819;
  wire _70821 = uncoded_block[1591] ^ uncoded_block[1617];
  wire _70822 = _70821 ^ uncoded_block[1666];
  wire _70823 = _70820 ^ _70822;
  wire _70824 = _70817 ^ _70823;
  wire _70825 = _70811 ^ _70824;
  wire _70826 = uncoded_block[34] ^ uncoded_block[69];
  wire _70827 = uncoded_block[126] ^ uncoded_block[205];
  wire _70828 = _70826 ^ _70827;
  wire _70829 = uncoded_block[259] ^ uncoded_block[297];
  wire _70830 = uncoded_block[407] ^ uncoded_block[492];
  wire _70831 = _70829 ^ _70830;
  wire _70832 = _70828 ^ _70831;
  wire _70833 = uncoded_block[552] ^ uncoded_block[615];
  wire _70834 = uncoded_block[667] ^ uncoded_block[714];
  wire _70835 = _70833 ^ _70834;
  wire _70836 = uncoded_block[773] ^ uncoded_block[801];
  wire _70837 = uncoded_block[843] ^ uncoded_block[929];
  wire _70838 = _70836 ^ _70837;
  wire _70839 = _70835 ^ _70838;
  wire _70840 = _70832 ^ _70839;
  wire _70841 = uncoded_block[969] ^ uncoded_block[1009];
  wire _70842 = uncoded_block[1093] ^ uncoded_block[1166];
  wire _70843 = _70841 ^ _70842;
  wire _70844 = uncoded_block[1191] ^ uncoded_block[1264];
  wire _70845 = uncoded_block[1314] ^ uncoded_block[1456];
  wire _70846 = _70844 ^ _70845;
  wire _70847 = _70843 ^ _70846;
  wire _70848 = uncoded_block[1496] ^ uncoded_block[1533];
  wire _70849 = uncoded_block[1543] ^ uncoded_block[1578];
  wire _70850 = _70848 ^ _70849;
  wire _70851 = uncoded_block[1644] ^ uncoded_block[1653];
  wire _70852 = _70851 ^ uncoded_block[1688];
  wire _70853 = _70850 ^ _70852;
  wire _70854 = _70847 ^ _70853;
  wire _70855 = _70840 ^ _70854;
  wire _70856 = uncoded_block[38] ^ uncoded_block[94];
  wire _70857 = uncoded_block[116] ^ uncoded_block[184];
  wire _70858 = _70856 ^ _70857;
  wire _70859 = _65353 ^ _65359;
  wire _70860 = _70858 ^ _70859;
  wire _70861 = uncoded_block[565] ^ uncoded_block[621];
  wire _70862 = _65363 ^ _70861;
  wire _70863 = uncoded_block[795] ^ uncoded_block[863];
  wire _70864 = _65372 ^ _70863;
  wire _70865 = _70862 ^ _70864;
  wire _70866 = _70860 ^ _70865;
  wire _70867 = uncoded_block[905] ^ uncoded_block[984];
  wire _70868 = _70867 ^ _66726;
  wire _70869 = uncoded_block[1127] ^ uncoded_block[1175];
  wire _70870 = uncoded_block[1260] ^ uncoded_block[1313];
  wire _70871 = _70869 ^ _70870;
  wire _70872 = _70868 ^ _70871;
  wire _70873 = uncoded_block[1346] ^ uncoded_block[1406];
  wire _70874 = uncoded_block[1433] ^ uncoded_block[1455];
  wire _70875 = _70873 ^ _70874;
  wire _70876 = uncoded_block[1621] ^ uncoded_block[1657];
  wire _70877 = _70876 ^ uncoded_block[1706];
  wire _70878 = _70875 ^ _70877;
  wire _70879 = _70872 ^ _70878;
  wire _70880 = _70866 ^ _70879;
  wire _70881 = uncoded_block[40] ^ uncoded_block[79];
  wire _70882 = _70881 ^ _67400;
  wire _70883 = uncoded_block[344] ^ uncoded_block[433];
  wire _70884 = _69095 ^ _70883;
  wire _70885 = _70882 ^ _70884;
  wire _70886 = uncoded_block[466] ^ uncoded_block[518];
  wire _70887 = uncoded_block[612] ^ uncoded_block[646];
  wire _70888 = _70886 ^ _70887;
  wire _70889 = uncoded_block[680] ^ uncoded_block[737];
  wire _70890 = uncoded_block[805] ^ uncoded_block[869];
  wire _70891 = _70889 ^ _70890;
  wire _70892 = _70888 ^ _70891;
  wire _70893 = _70885 ^ _70892;
  wire _70894 = uncoded_block[900] ^ uncoded_block[991];
  wire _70895 = uncoded_block[1057] ^ uncoded_block[1100];
  wire _70896 = _70894 ^ _70895;
  wire _70897 = uncoded_block[1153] ^ uncoded_block[1180];
  wire _70898 = _70897 ^ _67444;
  wire _70899 = _70896 ^ _70898;
  wire _70900 = uncoded_block[1383] ^ uncoded_block[1442];
  wire _70901 = _70900 ^ _67455;
  wire _70902 = uncoded_block[1609] ^ uncoded_block[1683];
  wire _70903 = _70902 ^ uncoded_block[1707];
  wire _70904 = _70901 ^ _70903;
  wire _70905 = _70899 ^ _70904;
  wire _70906 = _70893 ^ _70905;
  wire _70907 = uncoded_block[41] ^ uncoded_block[109];
  wire _70908 = uncoded_block[118] ^ uncoded_block[216];
  wire _70909 = _70907 ^ _70908;
  wire _70910 = uncoded_block[266] ^ uncoded_block[325];
  wire _70911 = uncoded_block[360] ^ uncoded_block[412];
  wire _70912 = _70910 ^ _70911;
  wire _70913 = _70909 ^ _70912;
  wire _70914 = uncoded_block[464] ^ uncoded_block[559];
  wire _70915 = uncoded_block[570] ^ uncoded_block[652];
  wire _70916 = _70914 ^ _70915;
  wire _70917 = uncoded_block[705] ^ uncoded_block[775];
  wire _70918 = uncoded_block[792] ^ uncoded_block[921];
  wire _70919 = _70917 ^ _70918;
  wire _70920 = _70916 ^ _70919;
  wire _70921 = _70913 ^ _70920;
  wire _70922 = uncoded_block[987] ^ uncoded_block[1029];
  wire _70923 = uncoded_block[1072] ^ uncoded_block[1114];
  wire _70924 = _70922 ^ _70923;
  wire _70925 = uncoded_block[1176] ^ uncoded_block[1233];
  wire _70926 = uncoded_block[1309] ^ uncoded_block[1335];
  wire _70927 = _70925 ^ _70926;
  wire _70928 = _70924 ^ _70927;
  wire _70929 = uncoded_block[1391] ^ uncoded_block[1430];
  wire _70930 = uncoded_block[1449] ^ uncoded_block[1459];
  wire _70931 = _70929 ^ _70930;
  wire _70932 = uncoded_block[1616] ^ uncoded_block[1678];
  wire _70933 = _70932 ^ uncoded_block[1711];
  wire _70934 = _70931 ^ _70933;
  wire _70935 = _70928 ^ _70934;
  wire _70936 = _70921 ^ _70935;
  wire _70937 = uncoded_block[51] ^ uncoded_block[85];
  wire _70938 = uncoded_block[166] ^ uncoded_block[194];
  wire _70939 = _70937 ^ _70938;
  wire _70940 = uncoded_block[232] ^ uncoded_block[317];
  wire _70941 = uncoded_block[363] ^ uncoded_block[428];
  wire _70942 = _70940 ^ _70941;
  wire _70943 = _70939 ^ _70942;
  wire _70944 = uncoded_block[463] ^ uncoded_block[536];
  wire _70945 = _70944 ^ _64807;
  wire _70946 = uncoded_block[671] ^ uncoded_block[750];
  wire _70947 = _70946 ^ _70143;
  wire _70948 = _70945 ^ _70947;
  wire _70949 = _70943 ^ _70948;
  wire _70950 = uncoded_block[933] ^ uncoded_block[999];
  wire _70951 = uncoded_block[1016] ^ uncoded_block[1076];
  wire _70952 = _70950 ^ _70951;
  wire _70953 = uncoded_block[1108] ^ uncoded_block[1162];
  wire _70954 = _70953 ^ _66623;
  wire _70955 = _70952 ^ _70954;
  wire _70956 = uncoded_block[1303] ^ uncoded_block[1354];
  wire _70957 = _70956 ^ _66629;
  wire _70958 = uncoded_block[1484] ^ uncoded_block[1652];
  wire _70959 = _70958 ^ uncoded_block[1690];
  wire _70960 = _70957 ^ _70959;
  wire _70961 = _70955 ^ _70960;
  wire _70962 = _70949 ^ _70961;
  wire _70963 = uncoded_block[0] ^ uncoded_block[87];
  wire _70964 = uncoded_block[151] ^ uncoded_block[189];
  wire _70965 = _70963 ^ _70964;
  wire _70966 = uncoded_block[248] ^ uncoded_block[280];
  wire _70967 = uncoded_block[357] ^ uncoded_block[404];
  wire _70968 = _70966 ^ _70967;
  wire _70969 = _70965 ^ _70968;
  wire _70970 = uncoded_block[497] ^ uncoded_block[559];
  wire _70971 = uncoded_block[592] ^ uncoded_block[643];
  wire _70972 = _70970 ^ _70971;
  wire _70973 = uncoded_block[717] ^ uncoded_block[729];
  wire _70974 = uncoded_block[801] ^ uncoded_block[831];
  wire _70975 = _70973 ^ _70974;
  wire _70976 = _70972 ^ _70975;
  wire _70977 = _70969 ^ _70976;
  wire _70978 = uncoded_block[920] ^ uncoded_block[1002];
  wire _70979 = uncoded_block[1051] ^ uncoded_block[1104];
  wire _70980 = _70978 ^ _70979;
  wire _70981 = uncoded_block[1257] ^ uncoded_block[1279];
  wire _70982 = _68085 ^ _70981;
  wire _70983 = _70980 ^ _70982;
  wire _70984 = uncoded_block[1377] ^ uncoded_block[1401];
  wire _70985 = uncoded_block[1431] ^ uncoded_block[1490];
  wire _70986 = _70984 ^ _70985;
  wire _70987 = uncoded_block[1529] ^ uncoded_block[1597];
  wire _70988 = _70987 ^ uncoded_block[1658];
  wire _70989 = _70986 ^ _70988;
  wire _70990 = _70983 ^ _70989;
  wire _70991 = _70977 ^ _70990;
  wire _70992 = uncoded_block[2] ^ uncoded_block[69];
  wire _70993 = uncoded_block[161] ^ uncoded_block[185];
  wire _70994 = _70992 ^ _70993;
  wire _70995 = uncoded_block[226] ^ uncoded_block[302];
  wire _70996 = _70995 ^ _69979;
  wire _70997 = _70994 ^ _70996;
  wire _70998 = _69982 ^ _69988;
  wire _70999 = uncoded_block[707] ^ uncoded_block[748];
  wire _71000 = uncoded_block[815] ^ uncoded_block[863];
  wire _71001 = _70999 ^ _71000;
  wire _71002 = _70998 ^ _71001;
  wire _71003 = _70997 ^ _71002;
  wire _71004 = uncoded_block[903] ^ uncoded_block[972];
  wire _71005 = _71004 ^ _70001;
  wire _71006 = uncoded_block[1158] ^ uncoded_block[1194];
  wire _71007 = uncoded_block[1222] ^ uncoded_block[1311];
  wire _71008 = _71006 ^ _71007;
  wire _71009 = _71005 ^ _71008;
  wire _71010 = uncoded_block[1345] ^ uncoded_block[1384];
  wire _71011 = uncoded_block[1524] ^ uncoded_block[1540];
  wire _71012 = _71010 ^ _71011;
  wire _71013 = uncoded_block[1630] ^ uncoded_block[1661];
  wire _71014 = _71013 ^ uncoded_block[1709];
  wire _71015 = _71012 ^ _71014;
  wire _71016 = _71009 ^ _71015;
  wire _71017 = _71003 ^ _71016;
  wire _71018 = uncoded_block[9] ^ uncoded_block[103];
  wire _71019 = uncoded_block[113] ^ uncoded_block[179];
  wire _71020 = _71018 ^ _71019;
  wire _71021 = uncoded_block[236] ^ uncoded_block[294];
  wire _71022 = uncoded_block[383] ^ uncoded_block[416];
  wire _71023 = _71021 ^ _71022;
  wire _71024 = _71020 ^ _71023;
  wire _71025 = uncoded_block[582] ^ uncoded_block[641];
  wire _71026 = _61621 ^ _71025;
  wire _71027 = uncoded_block[687] ^ uncoded_block[728];
  wire _71028 = uncoded_block[824] ^ uncoded_block[837];
  wire _71029 = _71027 ^ _71028;
  wire _71030 = _71026 ^ _71029;
  wire _71031 = _71024 ^ _71030;
  wire _71032 = uncoded_block[891] ^ uncoded_block[948];
  wire _71033 = uncoded_block[1028] ^ uncoded_block[1059];
  wire _71034 = _71032 ^ _71033;
  wire _71035 = uncoded_block[1079] ^ uncoded_block[1145];
  wire _71036 = uncoded_block[1182] ^ uncoded_block[1297];
  wire _71037 = _71035 ^ _71036;
  wire _71038 = _71034 ^ _71037;
  wire _71039 = uncoded_block[1374] ^ uncoded_block[1469];
  wire _71040 = uncoded_block[1521] ^ uncoded_block[1547];
  wire _71041 = _71039 ^ _71040;
  wire _71042 = uncoded_block[1593] ^ uncoded_block[1643];
  wire _71043 = _71042 ^ uncoded_block[1715];
  wire _71044 = _71041 ^ _71043;
  wire _71045 = _71038 ^ _71044;
  wire _71046 = _71031 ^ _71045;
  wire _71047 = uncoded_block[11] ^ uncoded_block[104];
  wire _71048 = uncoded_block[155] ^ uncoded_block[221];
  wire _71049 = _71047 ^ _71048;
  wire _71050 = uncoded_block[271] ^ uncoded_block[310];
  wire _71051 = uncoded_block[390] ^ uncoded_block[410];
  wire _71052 = _71050 ^ _71051;
  wire _71053 = _71049 ^ _71052;
  wire _71054 = uncoded_block[475] ^ uncoded_block[527];
  wire _71055 = uncoded_block[608] ^ uncoded_block[653];
  wire _71056 = _71054 ^ _71055;
  wire _71057 = uncoded_block[698] ^ uncoded_block[742];
  wire _71058 = uncoded_block[810] ^ uncoded_block[851];
  wire _71059 = _71057 ^ _71058;
  wire _71060 = _71056 ^ _71059;
  wire _71061 = _71053 ^ _71060;
  wire _71062 = uncoded_block[927] ^ uncoded_block[984];
  wire _71063 = uncoded_block[1020] ^ uncoded_block[1083];
  wire _71064 = _71062 ^ _71063;
  wire _71065 = uncoded_block[1244] ^ uncoded_block[1278];
  wire _71066 = uncoded_block[1293] ^ uncoded_block[1350];
  wire _71067 = _71065 ^ _71066;
  wire _71068 = _71064 ^ _71067;
  wire _71069 = _69019 ^ _751;
  wire _71070 = uncoded_block[1592] ^ uncoded_block[1636];
  wire _71071 = _71070 ^ uncoded_block[1669];
  wire _71072 = _71069 ^ _71071;
  wire _71073 = _71068 ^ _71072;
  wire _71074 = _71061 ^ _71073;
  wire _71075 = uncoded_block[19] ^ uncoded_block[63];
  wire _71076 = uncoded_block[140] ^ uncoded_block[178];
  wire _71077 = _71075 ^ _71076;
  wire _71078 = uncoded_block[258] ^ uncoded_block[314];
  wire _71079 = uncoded_block[368] ^ uncoded_block[417];
  wire _71080 = _71078 ^ _71079;
  wire _71081 = _71077 ^ _71080;
  wire _71082 = uncoded_block[454] ^ uncoded_block[555];
  wire _71083 = _71082 ^ _68315;
  wire _71084 = uncoded_block[691] ^ uncoded_block[746];
  wire _71085 = uncoded_block[807] ^ uncoded_block[874];
  wire _71086 = _71084 ^ _71085;
  wire _71087 = _71083 ^ _71086;
  wire _71088 = _71081 ^ _71087;
  wire _71089 = uncoded_block[1018] ^ uncoded_block[1075];
  wire _71090 = _68328 ^ _71089;
  wire _71091 = uncoded_block[1123] ^ uncoded_block[1198];
  wire _71092 = uncoded_block[1227] ^ uncoded_block[1322];
  wire _71093 = _71091 ^ _71092;
  wire _71094 = _71090 ^ _71093;
  wire _71095 = uncoded_block[1445] ^ uncoded_block[1575];
  wire _71096 = _68343 ^ _71095;
  wire _71097 = uncoded_block[1595] ^ uncoded_block[1631];
  wire _71098 = _71097 ^ uncoded_block[1706];
  wire _71099 = _71096 ^ _71098;
  wire _71100 = _71094 ^ _71099;
  wire _71101 = _71088 ^ _71100;
  wire _71102 = uncoded_block[22] ^ uncoded_block[90];
  wire _71103 = uncoded_block[135] ^ uncoded_block[193];
  wire _71104 = _71102 ^ _71103;
  wire _71105 = uncoded_block[270] ^ uncoded_block[328];
  wire _71106 = uncoded_block[366] ^ uncoded_block[419];
  wire _71107 = _71105 ^ _71106;
  wire _71108 = _71104 ^ _71107;
  wire _71109 = uncoded_block[472] ^ uncoded_block[520];
  wire _71110 = uncoded_block[623] ^ uncoded_block[718];
  wire _71111 = _71109 ^ _71110;
  wire _71112 = uncoded_block[865] ^ uncoded_block[914];
  wire _71113 = _11022 ^ _71112;
  wire _71114 = _71111 ^ _71113;
  wire _71115 = _71108 ^ _71114;
  wire _71116 = uncoded_block[967] ^ uncoded_block[1022];
  wire _71117 = uncoded_block[1066] ^ uncoded_block[1112];
  wire _71118 = _71116 ^ _71117;
  wire _71119 = uncoded_block[1174] ^ uncoded_block[1228];
  wire _71120 = uncoded_block[1284] ^ uncoded_block[1373];
  wire _71121 = _71119 ^ _71120;
  wire _71122 = _71118 ^ _71121;
  wire _71123 = uncoded_block[1411] ^ uncoded_block[1442];
  wire _71124 = uncoded_block[1480] ^ uncoded_block[1511];
  wire _71125 = _71123 ^ _71124;
  wire _71126 = uncoded_block[1615] ^ uncoded_block[1655];
  wire _71127 = _71126 ^ uncoded_block[1708];
  wire _71128 = _71125 ^ _71127;
  wire _71129 = _71122 ^ _71128;
  wire _71130 = _71115 ^ _71129;
  wire _71131 = uncoded_block[23] ^ uncoded_block[76];
  wire _71132 = uncoded_block[162] ^ uncoded_block[224];
  wire _71133 = _71131 ^ _71132;
  wire _71134 = uncoded_block[229] ^ uncoded_block[309];
  wire _71135 = uncoded_block[338] ^ uncoded_block[411];
  wire _71136 = _71134 ^ _71135;
  wire _71137 = _71133 ^ _71136;
  wire _71138 = uncoded_block[469] ^ uncoded_block[543];
  wire _71139 = uncoded_block[579] ^ uncoded_block[645];
  wire _71140 = _71138 ^ _71139;
  wire _71141 = uncoded_block[696] ^ uncoded_block[788];
  wire _71142 = uncoded_block[846] ^ uncoded_block[917];
  wire _71143 = _71141 ^ _71142;
  wire _71144 = _71140 ^ _71143;
  wire _71145 = _71137 ^ _71144;
  wire _71146 = uncoded_block[965] ^ uncoded_block[1011];
  wire _71147 = uncoded_block[1062] ^ uncoded_block[1136];
  wire _71148 = _71146 ^ _71147;
  wire _71149 = uncoded_block[1169] ^ uncoded_block[1207];
  wire _71150 = uncoded_block[1264] ^ uncoded_block[1325];
  wire _71151 = _71149 ^ _71150;
  wire _71152 = _71148 ^ _71151;
  wire _71153 = uncoded_block[1336] ^ uncoded_block[1406];
  wire _71154 = uncoded_block[1474] ^ uncoded_block[1577];
  wire _71155 = _71153 ^ _71154;
  wire _71156 = uncoded_block[1620] ^ uncoded_block[1659];
  wire _71157 = _71156 ^ uncoded_block[1714];
  wire _71158 = _71155 ^ _71157;
  wire _71159 = _71152 ^ _71158;
  wire _71160 = _71145 ^ _71159;
  wire _71161 = uncoded_block[26] ^ uncoded_block[83];
  wire _71162 = _71161 ^ _60941;
  wire _71163 = uncoded_block[256] ^ uncoded_block[305];
  wire _71164 = uncoded_block[356] ^ uncoded_block[447];
  wire _71165 = _71163 ^ _71164;
  wire _71166 = _71162 ^ _71165;
  wire _71167 = uncoded_block[457] ^ uncoded_block[525];
  wire _71168 = uncoded_block[568] ^ uncoded_block[659];
  wire _71169 = _71167 ^ _71168;
  wire _71170 = uncoded_block[675] ^ uncoded_block[754];
  wire _71171 = uncoded_block[781] ^ uncoded_block[855];
  wire _71172 = _71170 ^ _71171;
  wire _71173 = _71169 ^ _71172;
  wire _71174 = _71166 ^ _71173;
  wire _71175 = uncoded_block[902] ^ uncoded_block[950];
  wire _71176 = uncoded_block[1004] ^ uncoded_block[1082];
  wire _71177 = _71175 ^ _71176;
  wire _71178 = uncoded_block[1140] ^ uncoded_block[1179];
  wire _71179 = uncoded_block[1233] ^ uncoded_block[1282];
  wire _71180 = _71178 ^ _71179;
  wire _71181 = _71177 ^ _71180;
  wire _71182 = uncoded_block[1289] ^ uncoded_block[1381];
  wire _71183 = uncoded_block[1420] ^ uncoded_block[1475];
  wire _71184 = _71182 ^ _71183;
  wire _71185 = uncoded_block[1594] ^ uncoded_block[1629];
  wire _71186 = _71185 ^ uncoded_block[1656];
  wire _71187 = _71184 ^ _71186;
  wire _71188 = _71181 ^ _71187;
  wire _71189 = _71174 ^ _71188;
  wire _71190 = uncoded_block[28] ^ uncoded_block[77];
  wire _71191 = uncoded_block[154] ^ uncoded_block[202];
  wire _71192 = _71190 ^ _71191;
  wire _71193 = uncoded_block[261] ^ uncoded_block[295];
  wire _71194 = uncoded_block[375] ^ uncoded_block[432];
  wire _71195 = _71193 ^ _71194;
  wire _71196 = _71192 ^ _71195;
  wire _71197 = uncoded_block[483] ^ uncoded_block[508];
  wire _71198 = uncoded_block[616] ^ uncoded_block[651];
  wire _71199 = _71197 ^ _71198;
  wire _71200 = uncoded_block[693] ^ uncoded_block[757];
  wire _71201 = uncoded_block[811] ^ uncoded_block[871];
  wire _71202 = _71200 ^ _71201;
  wire _71203 = _71199 ^ _71202;
  wire _71204 = _71196 ^ _71203;
  wire _71205 = uncoded_block[915] ^ uncoded_block[956];
  wire _71206 = uncoded_block[1013] ^ uncoded_block[1076];
  wire _71207 = _71205 ^ _71206;
  wire _71208 = uncoded_block[1148] ^ uncoded_block[1177];
  wire _71209 = uncoded_block[1225] ^ uncoded_block[1277];
  wire _71210 = _71208 ^ _71209;
  wire _71211 = _71207 ^ _71210;
  wire _71212 = uncoded_block[1313] ^ uncoded_block[1352];
  wire _71213 = uncoded_block[1397] ^ uncoded_block[1436];
  wire _71214 = _71212 ^ _71213;
  wire _71215 = uncoded_block[1492] ^ uncoded_block[1586];
  wire _71216 = _71215 ^ uncoded_block[1698];
  wire _71217 = _71214 ^ _71216;
  wire _71218 = _71211 ^ _71217;
  wire _71219 = _71204 ^ _71218;
  wire _71220 = uncoded_block[29] ^ uncoded_block[75];
  wire _71221 = uncoded_block[126] ^ uncoded_block[201];
  wire _71222 = _71220 ^ _71221;
  wire _71223 = uncoded_block[227] ^ uncoded_block[329];
  wire _71224 = uncoded_block[339] ^ uncoded_block[414];
  wire _71225 = _71223 ^ _71224;
  wire _71226 = _71222 ^ _71225;
  wire _71227 = uncoded_block[501] ^ uncoded_block[524];
  wire _71228 = uncoded_block[574] ^ uncoded_block[627];
  wire _71229 = _71227 ^ _71228;
  wire _71230 = uncoded_block[681] ^ uncoded_block[747];
  wire _71231 = uncoded_block[797] ^ uncoded_block[860];
  wire _71232 = _71230 ^ _71231;
  wire _71233 = _71229 ^ _71232;
  wire _71234 = _71226 ^ _71233;
  wire _71235 = uncoded_block[941] ^ uncoded_block[961];
  wire _71236 = uncoded_block[1044] ^ uncoded_block[1078];
  wire _71237 = _71235 ^ _71236;
  wire _71238 = uncoded_block[1122] ^ uncoded_block[1204];
  wire _71239 = _71238 ^ _65720;
  wire _71240 = _71237 ^ _71239;
  wire _71241 = uncoded_block[1332] ^ uncoded_block[1362];
  wire _71242 = uncoded_block[1389] ^ uncoded_block[1542];
  wire _71243 = _71241 ^ _71242;
  wire _71244 = uncoded_block[1606] ^ uncoded_block[1628];
  wire _71245 = _71244 ^ uncoded_block[1667];
  wire _71246 = _71243 ^ _71245;
  wire _71247 = _71240 ^ _71246;
  wire _71248 = _71234 ^ _71247;
  wire _71249 = uncoded_block[31] ^ uncoded_block[85];
  wire _71250 = uncoded_block[130] ^ uncoded_block[216];
  wire _71251 = _71249 ^ _71250;
  wire _71252 = uncoded_block[234] ^ uncoded_block[311];
  wire _71253 = uncoded_block[377] ^ uncoded_block[446];
  wire _71254 = _71252 ^ _71253;
  wire _71255 = _71251 ^ _71254;
  wire _71256 = uncoded_block[505] ^ uncoded_block[556];
  wire _71257 = uncoded_block[607] ^ uncoded_block[621];
  wire _71258 = _71256 ^ _71257;
  wire _71259 = uncoded_block[676] ^ uncoded_block[724];
  wire _71260 = uncoded_block[825] ^ uncoded_block[841];
  wire _71261 = _71259 ^ _71260;
  wire _71262 = _71258 ^ _71261;
  wire _71263 = _71255 ^ _71262;
  wire _71264 = uncoded_block[922] ^ uncoded_block[990];
  wire _71265 = uncoded_block[1050] ^ uncoded_block[1085];
  wire _71266 = _71264 ^ _71265;
  wire _71267 = uncoded_block[1137] ^ uncoded_block[1215];
  wire _71268 = _71267 ^ _17907;
  wire _71269 = _71266 ^ _71268;
  wire _71270 = uncoded_block[1317] ^ uncoded_block[1361];
  wire _71271 = uncoded_block[1387] ^ uncoded_block[1425];
  wire _71272 = _71270 ^ _71271;
  wire _71273 = _19921 ^ uncoded_block[1651];
  wire _71274 = _71272 ^ _71273;
  wire _71275 = _71269 ^ _71274;
  wire _71276 = _71263 ^ _71275;
  wire _71277 = uncoded_block[32] ^ uncoded_block[59];
  wire _71278 = uncoded_block[145] ^ uncoded_block[220];
  wire _71279 = _71277 ^ _71278;
  wire _71280 = uncoded_block[240] ^ uncoded_block[308];
  wire _71281 = uncoded_block[369] ^ uncoded_block[445];
  wire _71282 = _71280 ^ _71281;
  wire _71283 = _71279 ^ _71282;
  wire _71284 = uncoded_block[451] ^ uncoded_block[515];
  wire _71285 = uncoded_block[615] ^ uncoded_block[661];
  wire _71286 = _71284 ^ _71285;
  wire _71287 = uncoded_block[674] ^ uncoded_block[764];
  wire _71288 = uncoded_block[806] ^ uncoded_block[852];
  wire _71289 = _71287 ^ _71288;
  wire _71290 = _71286 ^ _71289;
  wire _71291 = _71283 ^ _71290;
  wire _71292 = uncoded_block[940] ^ uncoded_block[973];
  wire _71293 = uncoded_block[1055] ^ uncoded_block[1095];
  wire _71294 = _71292 ^ _71293;
  wire _71295 = uncoded_block[1130] ^ uncoded_block[1209];
  wire _71296 = uncoded_block[1274] ^ uncoded_block[1295];
  wire _71297 = _71295 ^ _71296;
  wire _71298 = _71294 ^ _71297;
  wire _71299 = uncoded_block[1353] ^ uncoded_block[1402];
  wire _71300 = _71299 ^ _63953;
  wire _71301 = uncoded_block[1472] ^ uncoded_block[1623];
  wire _71302 = _71301 ^ uncoded_block[1677];
  wire _71303 = _71300 ^ _71302;
  wire _71304 = _71298 ^ _71303;
  wire _71305 = _71291 ^ _71304;
  wire _71306 = uncoded_block[36] ^ uncoded_block[60];
  wire _71307 = uncoded_block[129] ^ uncoded_block[180];
  wire _71308 = _71306 ^ _71307;
  wire _71309 = uncoded_block[246] ^ uncoded_block[330];
  wire _71310 = uncoded_block[335] ^ uncoded_block[395];
  wire _71311 = _71309 ^ _71310;
  wire _71312 = _71308 ^ _71311;
  wire _71313 = uncoded_block[462] ^ uncoded_block[547];
  wire _71314 = uncoded_block[598] ^ uncoded_block[630];
  wire _71315 = _71313 ^ _71314;
  wire _71316 = uncoded_block[671] ^ uncoded_block[731];
  wire _71317 = uncoded_block[818] ^ uncoded_block[867];
  wire _71318 = _71316 ^ _71317;
  wire _71319 = _71315 ^ _71318;
  wire _71320 = _71312 ^ _71319;
  wire _71321 = _68268 ^ _68271;
  wire _71322 = uncoded_block[1116] ^ uncoded_block[1164];
  wire _71323 = _71322 ^ _68276;
  wire _71324 = _71321 ^ _71323;
  wire _71325 = uncoded_block[1287] ^ uncoded_block[1341];
  wire _71326 = uncoded_block[1408] ^ uncoded_block[1441];
  wire _71327 = _71325 ^ _71326;
  wire _71328 = uncoded_block[1459] ^ uncoded_block[1491];
  wire _71329 = _71328 ^ uncoded_block[1694];
  wire _71330 = _71327 ^ _71329;
  wire _71331 = _71324 ^ _71330;
  wire _71332 = _71320 ^ _71331;
  wire _71333 = uncoded_block[45] ^ uncoded_block[102];
  wire _71334 = uncoded_block[134] ^ uncoded_block[204];
  wire _71335 = _71333 ^ _71334;
  wire _71336 = uncoded_block[245] ^ uncoded_block[300];
  wire _71337 = _71336 ^ _65677;
  wire _71338 = _71335 ^ _71337;
  wire _71339 = uncoded_block[448] ^ uncoded_block[554];
  wire _71340 = uncoded_block[570] ^ uncoded_block[628];
  wire _71341 = _71339 ^ _71340;
  wire _71342 = uncoded_block[711] ^ uncoded_block[760];
  wire _71343 = uncoded_block[820] ^ uncoded_block[856];
  wire _71344 = _71342 ^ _71343;
  wire _71345 = _71341 ^ _71344;
  wire _71346 = _71338 ^ _71345;
  wire _71347 = uncoded_block[919] ^ uncoded_block[946];
  wire _71348 = _71347 ^ _67595;
  wire _71349 = uncoded_block[1139] ^ uncoded_block[1210];
  wire _71350 = uncoded_block[1241] ^ uncoded_block[1356];
  wire _71351 = _71349 ^ _71350;
  wire _71352 = _71348 ^ _71351;
  wire _71353 = uncoded_block[1386] ^ uncoded_block[1446];
  wire _71354 = uncoded_block[1532] ^ uncoded_block[1576];
  wire _71355 = _71353 ^ _71354;
  wire _71356 = uncoded_block[1613] ^ uncoded_block[1685];
  wire _71357 = _71356 ^ uncoded_block[1707];
  wire _71358 = _71355 ^ _71357;
  wire _71359 = _71352 ^ _71358;
  wire _71360 = _71346 ^ _71359;
  wire _71361 = uncoded_block[47] ^ uncoded_block[105];
  wire _71362 = uncoded_block[111] ^ uncoded_block[208];
  wire _71363 = _71361 ^ _71362;
  wire _71364 = uncoded_block[254] ^ uncoded_block[316];
  wire _71365 = uncoded_block[379] ^ uncoded_block[415];
  wire _71366 = _71364 ^ _71365;
  wire _71367 = _71363 ^ _71366;
  wire _71368 = uncoded_block[484] ^ uncoded_block[526];
  wire _71369 = _71368 ^ _60980;
  wire _71370 = uncoded_block[692] ^ uncoded_block[739];
  wire _71371 = uncoded_block[789] ^ uncoded_block[859];
  wire _71372 = _71370 ^ _71371;
  wire _71373 = _71369 ^ _71372;
  wire _71374 = _71367 ^ _71373;
  wire _71375 = uncoded_block[895] ^ uncoded_block[977];
  wire _71376 = uncoded_block[1057] ^ uncoded_block[1146];
  wire _71377 = _71375 ^ _71376;
  wire _71378 = uncoded_block[1348] ^ uncoded_block[1422];
  wire _71379 = _67705 ^ _71378;
  wire _71380 = _71377 ^ _71379;
  wire _71381 = uncoded_block[1440] ^ uncoded_block[1484];
  wire _71382 = uncoded_block[1487] ^ uncoded_block[1509];
  wire _71383 = _71381 ^ _71382;
  wire _71384 = uncoded_block[1527] ^ uncoded_block[1674];
  wire _71385 = _71384 ^ uncoded_block[1689];
  wire _71386 = _71383 ^ _71385;
  wire _71387 = _71380 ^ _71386;
  wire _71388 = _71374 ^ _71387;
  wire _71389 = uncoded_block[48] ^ uncoded_block[96];
  wire _71390 = uncoded_block[150] ^ uncoded_block[213];
  wire _71391 = _71389 ^ _71390;
  wire _71392 = uncoded_block[273] ^ uncoded_block[320];
  wire _71393 = uncoded_block[363] ^ uncoded_block[504];
  wire _71394 = _71392 ^ _71393;
  wire _71395 = _71391 ^ _71394;
  wire _71396 = uncoded_block[523] ^ uncoded_block[614];
  wire _71397 = uncoded_block[636] ^ uncoded_block[703];
  wire _71398 = _71396 ^ _71397;
  wire _71399 = uncoded_block[732] ^ uncoded_block[872];
  wire _71400 = uncoded_block[887] ^ uncoded_block[913];
  wire _71401 = _71399 ^ _71400;
  wire _71402 = _71398 ^ _71401;
  wire _71403 = _71395 ^ _71402;
  wire _71404 = uncoded_block[958] ^ uncoded_block[1040];
  wire _71405 = uncoded_block[1068] ^ uncoded_block[1153];
  wire _71406 = _71404 ^ _71405;
  wire _71407 = uncoded_block[1184] ^ uncoded_block[1246];
  wire _71408 = uncoded_block[1312] ^ uncoded_block[1351];
  wire _71409 = _71407 ^ _71408;
  wire _71410 = _71406 ^ _71409;
  wire _71411 = uncoded_block[1403] ^ uncoded_block[1457];
  wire _71412 = uncoded_block[1481] ^ uncoded_block[1500];
  wire _71413 = _71411 ^ _71412;
  wire _71414 = uncoded_block[1634] ^ uncoded_block[1670];
  wire _71415 = _71414 ^ uncoded_block[1701];
  wire _71416 = _71413 ^ _71415;
  wire _71417 = _71410 ^ _71416;
  wire _71418 = _71403 ^ _71417;
  wire _71419 = uncoded_block[52] ^ uncoded_block[59];
  wire _71420 = uncoded_block[138] ^ uncoded_block[185];
  wire _71421 = _71419 ^ _71420;
  wire _71422 = uncoded_block[270] ^ uncoded_block[280];
  wire _71423 = uncoded_block[393] ^ uncoded_block[486];
  wire _71424 = _71422 ^ _71423;
  wire _71425 = _71421 ^ _71424;
  wire _71426 = uncoded_block[659] ^ uncoded_block[719];
  wire _71427 = _67265 ^ _71426;
  wire _71428 = uncoded_block[757] ^ uncoded_block[778];
  wire _71429 = uncoded_block[859] ^ uncoded_block[889];
  wire _71430 = _71428 ^ _71429;
  wire _71431 = _71427 ^ _71430;
  wire _71432 = _71425 ^ _71431;
  wire _71433 = uncoded_block[1078] ^ uncoded_block[1161];
  wire _71434 = _67022 ^ _71433;
  wire _71435 = uncoded_block[1236] ^ uncoded_block[1322];
  wire _71436 = _27912 ^ _71435;
  wire _71437 = _71434 ^ _71436;
  wire _71438 = uncoded_block[1333] ^ uncoded_block[1380];
  wire _71439 = uncoded_block[1548] ^ uncoded_block[1585];
  wire _71440 = _71438 ^ _71439;
  wire _71441 = uncoded_block[1634] ^ uncoded_block[1684];
  wire _71442 = _71441 ^ uncoded_block[1703];
  wire _71443 = _71440 ^ _71442;
  wire _71444 = _71437 ^ _71443;
  wire _71445 = _71432 ^ _71444;
  wire _71446 = uncoded_block[90] ^ uncoded_block[113];
  wire _71447 = uncoded_block[200] ^ uncoded_block[240];
  wire _71448 = _71446 ^ _71447;
  wire _71449 = uncoded_block[439] ^ uncoded_block[474];
  wire _71450 = _65299 ^ _71449;
  wire _71451 = _71448 ^ _71450;
  wire _71452 = uncoded_block[550] ^ uncoded_block[606];
  wire _71453 = _71452 ^ _65309;
  wire _71454 = uncoded_block[767] ^ uncoded_block[814];
  wire _71455 = _71454 ^ _65316;
  wire _71456 = _71453 ^ _71455;
  wire _71457 = _71451 ^ _71456;
  wire _71458 = uncoded_block[961] ^ uncoded_block[1035];
  wire _71459 = _71458 ^ _65325;
  wire _71460 = uncoded_block[1181] ^ uncoded_block[1263];
  wire _71461 = uncoded_block[1327] ^ uncoded_block[1378];
  wire _71462 = _71460 ^ _71461;
  wire _71463 = _71459 ^ _71462;
  wire _71464 = uncoded_block[1399] ^ uncoded_block[1554];
  wire _71465 = uncoded_block[1564] ^ uncoded_block[1590];
  wire _71466 = _71464 ^ _71465;
  wire _71467 = uncoded_block[1629] ^ uncoded_block[1672];
  wire _71468 = _71467 ^ uncoded_block[1722];
  wire _71469 = _71466 ^ _71468;
  wire _71470 = _71463 ^ _71469;
  wire _71471 = _71457 ^ _71470;
  wire _71472 = uncoded_block[0] ^ uncoded_block[106];
  wire _71473 = uncoded_block[153] ^ uncoded_block[193];
  wire _71474 = _71472 ^ _71473;
  wire _71475 = uncoded_block[226] ^ uncoded_block[318];
  wire _71476 = uncoded_block[354] ^ uncoded_block[444];
  wire _71477 = _71475 ^ _71476;
  wire _71478 = _71474 ^ _71477;
  wire _71479 = uncoded_block[484] ^ uncoded_block[545];
  wire _71480 = uncoded_block[603] ^ uncoded_block[658];
  wire _71481 = _71479 ^ _71480;
  wire _71482 = uncoded_block[783] ^ uncoded_block[850];
  wire _71483 = _65896 ^ _71482;
  wire _71484 = _71481 ^ _71483;
  wire _71485 = _71478 ^ _71484;
  wire _71486 = uncoded_block[909] ^ uncoded_block[1001];
  wire _71487 = _71486 ^ _65907;
  wire _71488 = uncoded_block[1125] ^ uncoded_block[1176];
  wire _71489 = uncoded_block[1305] ^ uncoded_block[1358];
  wire _71490 = _71488 ^ _71489;
  wire _71491 = _71487 ^ _71490;
  wire _71492 = uncoded_block[1412] ^ uncoded_block[1426];
  wire _71493 = uncoded_block[1463] ^ uncoded_block[1521];
  wire _71494 = _71492 ^ _71493;
  wire _71495 = uncoded_block[1558] ^ uncoded_block[1648];
  wire _71496 = _71495 ^ uncoded_block[1652];
  wire _71497 = _71494 ^ _71496;
  wire _71498 = _71491 ^ _71497;
  wire _71499 = _71485 ^ _71498;
  wire _71500 = uncoded_block[6] ^ uncoded_block[109];
  wire _71501 = uncoded_block[147] ^ uncoded_block[204];
  wire _71502 = _71500 ^ _71501;
  wire _71503 = uncoded_block[232] ^ uncoded_block[304];
  wire _71504 = uncoded_block[368] ^ uncoded_block[397];
  wire _71505 = _71503 ^ _71504;
  wire _71506 = _71502 ^ _71505;
  wire _71507 = uncoded_block[496] ^ uncoded_block[512];
  wire _71508 = uncoded_block[576] ^ uncoded_block[651];
  wire _71509 = _71507 ^ _71508;
  wire _71510 = uncoded_block[721] ^ uncoded_block[754];
  wire _71511 = uncoded_block[787] ^ uncoded_block[881];
  wire _71512 = _71510 ^ _71511;
  wire _71513 = _71509 ^ _71512;
  wire _71514 = _71506 ^ _71513;
  wire _71515 = uncoded_block[895] ^ uncoded_block[998];
  wire _71516 = uncoded_block[1027] ^ uncoded_block[1059];
  wire _71517 = _71515 ^ _71516;
  wire _71518 = uncoded_block[1093] ^ uncoded_block[1156];
  wire _71519 = uncoded_block[1320] ^ uncoded_block[1339];
  wire _71520 = _71518 ^ _71519;
  wire _71521 = _71517 ^ _71520;
  wire _71522 = uncoded_block[1472] ^ uncoded_block[1517];
  wire _71523 = _71522 ^ _63146;
  wire _71524 = uncoded_block[1597] ^ uncoded_block[1639];
  wire _71525 = _71524 ^ uncoded_block[1697];
  wire _71526 = _71523 ^ _71525;
  wire _71527 = _71521 ^ _71526;
  wire _71528 = _71514 ^ _71527;
  wire _71529 = uncoded_block[7] ^ uncoded_block[89];
  wire _71530 = _71529 ^ _67175;
  wire _71531 = uncoded_block[251] ^ uncoded_block[286];
  wire _71532 = uncoded_block[356] ^ uncoded_block[404];
  wire _71533 = _71531 ^ _71532;
  wire _71534 = _71530 ^ _71533;
  wire _71535 = uncoded_block[450] ^ uncoded_block[533];
  wire _71536 = uncoded_block[566] ^ uncoded_block[664];
  wire _71537 = _71535 ^ _71536;
  wire _71538 = uncoded_block[686] ^ uncoded_block[746];
  wire _71539 = uncoded_block[817] ^ uncoded_block[867];
  wire _71540 = _71538 ^ _71539;
  wire _71541 = _71537 ^ _71540;
  wire _71542 = _71534 ^ _71541;
  wire _71543 = uncoded_block[910] ^ uncoded_block[993];
  wire _71544 = uncoded_block[1032] ^ uncoded_block[1091];
  wire _71545 = _71543 ^ _71544;
  wire _71546 = uncoded_block[1202] ^ uncoded_block[1246];
  wire _71547 = _60567 ^ _71546;
  wire _71548 = _71545 ^ _71547;
  wire _71549 = uncoded_block[1313] ^ uncoded_block[1389];
  wire _71550 = _71549 ^ _67228;
  wire _71551 = uncoded_block[1549] ^ uncoded_block[1625];
  wire _71552 = _71551 ^ uncoded_block[1691];
  wire _71553 = _71550 ^ _71552;
  wire _71554 = _71548 ^ _71553;
  wire _71555 = _71542 ^ _71554;
  wire _71556 = uncoded_block[8] ^ uncoded_block[82];
  wire _71557 = uncoded_block[117] ^ uncoded_block[211];
  wire _71558 = _71556 ^ _71557;
  wire _71559 = uncoded_block[344] ^ uncoded_block[445];
  wire _71560 = _65936 ^ _71559;
  wire _71561 = _71558 ^ _71560;
  wire _71562 = uncoded_block[503] ^ uncoded_block[535];
  wire _71563 = uncoded_block[590] ^ uncoded_block[638];
  wire _71564 = _71562 ^ _71563;
  wire _71565 = uncoded_block[709] ^ uncoded_block[735];
  wire _71566 = _71565 ^ _68390;
  wire _71567 = _71564 ^ _71566;
  wire _71568 = _71561 ^ _71567;
  wire _71569 = uncoded_block[908] ^ uncoded_block[976];
  wire _71570 = uncoded_block[1106] ^ uncoded_block[1135];
  wire _71571 = _71569 ^ _71570;
  wire _71572 = uncoded_block[1164] ^ uncoded_block[1172];
  wire _71573 = uncoded_block[1260] ^ uncoded_block[1293];
  wire _71574 = _71572 ^ _71573;
  wire _71575 = _71571 ^ _71574;
  wire _71576 = uncoded_block[1340] ^ uncoded_block[1395];
  wire _71577 = uncoded_block[1438] ^ uncoded_block[1495];
  wire _71578 = _71576 ^ _71577;
  wire _71579 = uncoded_block[1505] ^ uncoded_block[1606];
  wire _71580 = _71579 ^ uncoded_block[1627];
  wire _71581 = _71578 ^ _71580;
  wire _71582 = _71575 ^ _71581;
  wire _71583 = _71568 ^ _71582;
  wire _71584 = uncoded_block[22] ^ uncoded_block[62];
  wire _71585 = uncoded_block[133] ^ uncoded_block[189];
  wire _71586 = _71584 ^ _71585;
  wire _71587 = uncoded_block[233] ^ uncoded_block[302];
  wire _71588 = uncoded_block[351] ^ uncoded_block[442];
  wire _71589 = _71587 ^ _71588;
  wire _71590 = _71586 ^ _71589;
  wire _71591 = uncoded_block[459] ^ uncoded_block[546];
  wire _71592 = _71591 ^ _59988;
  wire _71593 = uncoded_block[677] ^ uncoded_block[731];
  wire _71594 = uncoded_block[813] ^ uncoded_block[874];
  wire _71595 = _71593 ^ _71594;
  wire _71596 = _71592 ^ _71595;
  wire _71597 = _71590 ^ _71596;
  wire _71598 = uncoded_block[931] ^ uncoded_block[994];
  wire _71599 = uncoded_block[1030] ^ uncoded_block[1109];
  wire _71600 = _71598 ^ _71599;
  wire _71601 = uncoded_block[1144] ^ uncoded_block[1175];
  wire _71602 = uncoded_block[1249] ^ uncoded_block[1443];
  wire _71603 = _71601 ^ _71602;
  wire _71604 = _71600 ^ _71603;
  wire _71605 = uncoded_block[1576] ^ uncoded_block[1622];
  wire _71606 = _71605 ^ uncoded_block[1683];
  wire _71607 = _67158 ^ _71606;
  wire _71608 = _71604 ^ _71607;
  wire _71609 = _71597 ^ _71608;
  wire _71610 = uncoded_block[24] ^ uncoded_block[77];
  wire _71611 = uncoded_block[163] ^ uncoded_block[224];
  wire _71612 = _71610 ^ _71611;
  wire _71613 = uncoded_block[230] ^ uncoded_block[310];
  wire _71614 = uncoded_block[339] ^ uncoded_block[412];
  wire _71615 = _71613 ^ _71614;
  wire _71616 = _71612 ^ _71615;
  wire _71617 = uncoded_block[470] ^ uncoded_block[544];
  wire _71618 = uncoded_block[580] ^ uncoded_block[646];
  wire _71619 = _71617 ^ _71618;
  wire _71620 = uncoded_block[697] ^ uncoded_block[764];
  wire _71621 = uncoded_block[789] ^ uncoded_block[847];
  wire _71622 = _71620 ^ _71621;
  wire _71623 = _71619 ^ _71622;
  wire _71624 = _71616 ^ _71623;
  wire _71625 = uncoded_block[918] ^ uncoded_block[966];
  wire _71626 = uncoded_block[1012] ^ uncoded_block[1063];
  wire _71627 = _71625 ^ _71626;
  wire _71628 = uncoded_block[1137] ^ uncoded_block[1208];
  wire _71629 = uncoded_block[1218] ^ uncoded_block[1265];
  wire _71630 = _71628 ^ _71629;
  wire _71631 = _71627 ^ _71630;
  wire _71632 = uncoded_block[1326] ^ uncoded_block[1337];
  wire _71633 = uncoded_block[1407] ^ uncoded_block[1475];
  wire _71634 = _71632 ^ _71633;
  wire _71635 = uncoded_block[1578] ^ uncoded_block[1621];
  wire _71636 = _71635 ^ uncoded_block[1660];
  wire _71637 = _71634 ^ _71636;
  wire _71638 = _71631 ^ _71637;
  wire _71639 = _71624 ^ _71638;
  wire _71640 = uncoded_block[25] ^ uncoded_block[102];
  wire _71641 = uncoded_block[144] ^ uncoded_block[194];
  wire _71642 = _71640 ^ _71641;
  wire _71643 = uncoded_block[323] ^ uncoded_block[377];
  wire _71644 = uncoded_block[431] ^ uncoded_block[488];
  wire _71645 = _71643 ^ _71644;
  wire _71646 = _71642 ^ _71645;
  wire _71647 = uncoded_block[515] ^ uncoded_block[612];
  wire _71648 = uncoded_block[645] ^ uncoded_block[717];
  wire _71649 = _71647 ^ _71648;
  wire _71650 = uncoded_block[725] ^ uncoded_block[785];
  wire _71651 = uncoded_block[830] ^ uncoded_block[886];
  wire _71652 = _71650 ^ _71651;
  wire _71653 = _71649 ^ _71652;
  wire _71654 = _71646 ^ _71653;
  wire _71655 = uncoded_block[905] ^ uncoded_block[983];
  wire _71656 = uncoded_block[1029] ^ uncoded_block[1069];
  wire _71657 = _71655 ^ _71656;
  wire _71658 = uncoded_block[1122] ^ uncoded_block[1190];
  wire _71659 = uncoded_block[1269] ^ uncoded_block[1297];
  wire _71660 = _71658 ^ _71659;
  wire _71661 = _71657 ^ _71660;
  wire _71662 = uncoded_block[1368] ^ uncoded_block[1384];
  wire _71663 = uncoded_block[1392] ^ uncoded_block[1477];
  wire _71664 = _71662 ^ _71663;
  wire _71665 = uncoded_block[1612] ^ uncoded_block[1687];
  wire _71666 = _71665 ^ uncoded_block[1696];
  wire _71667 = _71664 ^ _71666;
  wire _71668 = _71661 ^ _71667;
  wire _71669 = _71654 ^ _71668;
  wire _71670 = uncoded_block[27] ^ uncoded_block[84];
  wire _71671 = _71670 ^ _61262;
  wire _71672 = uncoded_block[257] ^ uncoded_block[306];
  wire _71673 = uncoded_block[357] ^ uncoded_block[447];
  wire _71674 = _71672 ^ _71673;
  wire _71675 = _71671 ^ _71674;
  wire _71676 = uncoded_block[458] ^ uncoded_block[526];
  wire _71677 = uncoded_block[569] ^ uncoded_block[660];
  wire _71678 = _71676 ^ _71677;
  wire _71679 = uncoded_block[676] ^ uncoded_block[755];
  wire _71680 = uncoded_block[782] ^ uncoded_block[856];
  wire _71681 = _71679 ^ _71680;
  wire _71682 = _71678 ^ _71681;
  wire _71683 = _71675 ^ _71682;
  wire _71684 = uncoded_block[903] ^ uncoded_block[951];
  wire _71685 = uncoded_block[1005] ^ uncoded_block[1083];
  wire _71686 = _71684 ^ _71685;
  wire _71687 = uncoded_block[1141] ^ uncoded_block[1180];
  wire _71688 = _71687 ^ _70013;
  wire _71689 = _71686 ^ _71688;
  wire _71690 = uncoded_block[1329] ^ uncoded_block[1382];
  wire _71691 = uncoded_block[1421] ^ uncoded_block[1456];
  wire _71692 = _71690 ^ _71691;
  wire _71693 = uncoded_block[1595] ^ uncoded_block[1657];
  wire _71694 = _71693 ^ uncoded_block[1702];
  wire _71695 = _71692 ^ _71694;
  wire _71696 = _71689 ^ _71695;
  wire _71697 = _71683 ^ _71696;
  wire _71698 = uncoded_block[37] ^ uncoded_block[61];
  wire _71699 = uncoded_block[130] ^ uncoded_block[181];
  wire _71700 = _71698 ^ _71699;
  wire _71701 = uncoded_block[247] ^ uncoded_block[331];
  wire _71702 = uncoded_block[336] ^ uncoded_block[396];
  wire _71703 = _71701 ^ _71702;
  wire _71704 = _71700 ^ _71703;
  wire _71705 = uncoded_block[463] ^ uncoded_block[548];
  wire _71706 = uncoded_block[599] ^ uncoded_block[631];
  wire _71707 = _71705 ^ _71706;
  wire _71708 = uncoded_block[672] ^ uncoded_block[732];
  wire _71709 = uncoded_block[819] ^ uncoded_block[868];
  wire _71710 = _71708 ^ _71709;
  wire _71711 = _71707 ^ _71710;
  wire _71712 = _71704 ^ _71711;
  wire _71713 = uncoded_block[1024] ^ uncoded_block[1071];
  wire _71714 = _66562 ^ _71713;
  wire _71715 = uncoded_block[1191] ^ uncoded_block[1227];
  wire _71716 = _66568 ^ _71715;
  wire _71717 = _71714 ^ _71716;
  wire _71718 = uncoded_block[1288] ^ uncoded_block[1342];
  wire _71719 = uncoded_block[1409] ^ uncoded_block[1442];
  wire _71720 = _71718 ^ _71719;
  wire _71721 = uncoded_block[1460] ^ uncoded_block[1492];
  wire _71722 = _71721 ^ uncoded_block[1669];
  wire _71723 = _71720 ^ _71722;
  wire _71724 = _71717 ^ _71723;
  wire _71725 = _71712 ^ _71724;
  wire _71726 = uncoded_block[39] ^ uncoded_block[83];
  wire _71727 = uncoded_block[158] ^ uncoded_block[192];
  wire _71728 = _71726 ^ _71727;
  wire _71729 = uncoded_block[273] ^ uncoded_block[287];
  wire _71730 = uncoded_block[373] ^ uncoded_block[394];
  wire _71731 = _71729 ^ _71730;
  wire _71732 = _71728 ^ _71731;
  wire _71733 = uncoded_block[495] ^ uncoded_block[543];
  wire _71734 = uncoded_block[589] ^ uncoded_block[661];
  wire _71735 = _71733 ^ _71734;
  wire _71736 = uncoded_block[671] ^ uncoded_block[771];
  wire _71737 = uncoded_block[862] ^ uncoded_block[912];
  wire _71738 = _71736 ^ _71737;
  wire _71739 = _71735 ^ _71738;
  wire _71740 = _71732 ^ _71739;
  wire _71741 = uncoded_block[964] ^ uncoded_block[1008];
  wire _71742 = uncoded_block[1075] ^ uncoded_block[1145];
  wire _71743 = _71741 ^ _71742;
  wire _71744 = uncoded_block[1199] ^ uncoded_block[1252];
  wire _71745 = uncoded_block[1299] ^ uncoded_block[1360];
  wire _71746 = _71744 ^ _71745;
  wire _71747 = _71743 ^ _71746;
  wire _71748 = uncoded_block[1391] ^ uncoded_block[1436];
  wire _71749 = uncoded_block[1455] ^ uncoded_block[1592];
  wire _71750 = _71748 ^ _71749;
  wire _71751 = uncoded_block[1615] ^ uncoded_block[1679];
  wire _71752 = _71751 ^ uncoded_block[1688];
  wire _71753 = _71750 ^ _71752;
  wire _71754 = _71747 ^ _71753;
  wire _71755 = _71740 ^ _71754;
  wire _71756 = uncoded_block[41] ^ uncoded_block[80];
  wire _71757 = uncoded_block[170] ^ uncoded_block[191];
  wire _71758 = _71756 ^ _71757;
  wire _71759 = uncoded_block[277] ^ uncoded_block[293];
  wire _71760 = uncoded_block[346] ^ uncoded_block[435];
  wire _71761 = _71759 ^ _71760;
  wire _71762 = _71758 ^ _71761;
  wire _71763 = uncoded_block[467] ^ uncoded_block[519];
  wire _71764 = uncoded_block[614] ^ uncoded_block[648];
  wire _71765 = _71763 ^ _71764;
  wire _71766 = uncoded_block[681] ^ uncoded_block[739];
  wire _71767 = uncoded_block[806] ^ uncoded_block[871];
  wire _71768 = _71766 ^ _71767;
  wire _71769 = _71765 ^ _71768;
  wire _71770 = _71762 ^ _71769;
  wire _71771 = uncoded_block[902] ^ uncoded_block[992];
  wire _71772 = uncoded_block[1101] ^ uncoded_block[1154];
  wire _71773 = _71771 ^ _71772;
  wire _71774 = uncoded_block[1182] ^ uncoded_block[1261];
  wire _71775 = _71774 ^ _66960;
  wire _71776 = _71773 ^ _71775;
  wire _71777 = uncoded_block[1467] ^ uncoded_block[1504];
  wire _71778 = _71777 ^ _68424;
  wire _71779 = uncoded_block[1580] ^ uncoded_block[1611];
  wire _71780 = _71779 ^ uncoded_block[1708];
  wire _71781 = _71778 ^ _71780;
  wire _71782 = _71776 ^ _71781;
  wire _71783 = _71770 ^ _71782;
  wire _71784 = uncoded_block[116] ^ uncoded_block[172];
  wire _71785 = _33041 ^ _71784;
  wire _71786 = uncoded_block[276] ^ uncoded_block[305];
  wire _71787 = uncoded_block[372] ^ uncoded_block[402];
  wire _71788 = _71786 ^ _71787;
  wire _71789 = _71785 ^ _71788;
  wire _71790 = uncoded_block[493] ^ uncoded_block[547];
  wire _71791 = uncoded_block[596] ^ uncoded_block[643];
  wire _71792 = _71790 ^ _71791;
  wire _71793 = uncoded_block[696] ^ uncoded_block[824];
  wire _71794 = uncoded_block[857] ^ uncoded_block[939];
  wire _71795 = _71793 ^ _71794;
  wire _71796 = _71792 ^ _71795;
  wire _71797 = _71789 ^ _71796;
  wire _71798 = uncoded_block[954] ^ uncoded_block[1053];
  wire _71799 = _71798 ^ _69797;
  wire _71800 = uncoded_block[1209] ^ uncoded_block[1220];
  wire _71801 = uncoded_block[1291] ^ uncoded_block[1371];
  wire _71802 = _71800 ^ _71801;
  wire _71803 = _71799 ^ _71802;
  wire _71804 = uncoded_block[1499] ^ uncoded_block[1586];
  wire _71805 = _69808 ^ _71804;
  wire _71806 = uncoded_block[1617] ^ uncoded_block[1655];
  wire _71807 = _71806 ^ uncoded_block[1705];
  wire _71808 = _71805 ^ _71807;
  wire _71809 = _71803 ^ _71808;
  wire _71810 = _71797 ^ _71809;
  wire _71811 = uncoded_block[117] ^ uncoded_block[173];
  wire _71812 = _43266 ^ _71811;
  wire _71813 = uncoded_block[277] ^ uncoded_block[306];
  wire _71814 = _71813 ^ _66014;
  wire _71815 = _71812 ^ _71814;
  wire _71816 = uncoded_block[494] ^ uncoded_block[548];
  wire _71817 = _71816 ^ _66024;
  wire _71818 = uncoded_block[697] ^ uncoded_block[825];
  wire _71819 = uncoded_block[858] ^ uncoded_block[940];
  wire _71820 = _71818 ^ _71819;
  wire _71821 = _71817 ^ _71820;
  wire _71822 = _71815 ^ _71821;
  wire _71823 = uncoded_block[955] ^ uncoded_block[1054];
  wire _71824 = uncoded_block[1120] ^ uncoded_block[1210];
  wire _71825 = _71823 ^ _71824;
  wire _71826 = uncoded_block[1292] ^ uncoded_block[1372];
  wire _71827 = _66512 ^ _71826;
  wire _71828 = _71825 ^ _71827;
  wire _71829 = _66520 ^ _66523;
  wire _71830 = _66526 ^ uncoded_block[1706];
  wire _71831 = _71829 ^ _71830;
  wire _71832 = _71828 ^ _71831;
  wire _71833 = _71822 ^ _71832;
  wire _71834 = uncoded_block[4] ^ uncoded_block[68];
  wire _71835 = uncoded_block[137] ^ uncoded_block[209];
  wire _71836 = _71834 ^ _71835;
  wire _71837 = uncoded_block[264] ^ uncoded_block[315];
  wire _71838 = uncoded_block[372] ^ uncoded_block[433];
  wire _71839 = _71837 ^ _71838;
  wire _71840 = _71836 ^ _71839;
  wire _71841 = uncoded_block[473] ^ uncoded_block[537];
  wire _71842 = uncoded_block[564] ^ uncoded_block[654];
  wire _71843 = _71841 ^ _71842;
  wire _71844 = uncoded_block[688] ^ uncoded_block[771];
  wire _71845 = uncoded_block[789] ^ uncoded_block[864];
  wire _71846 = _71844 ^ _71845;
  wire _71847 = _71843 ^ _71846;
  wire _71848 = _71840 ^ _71847;
  wire _71849 = uncoded_block[920] ^ uncoded_block[992];
  wire _71850 = uncoded_block[1039] ^ uncoded_block[1111];
  wire _71851 = _71849 ^ _71850;
  wire _71852 = uncoded_block[1117] ^ uncoded_block[1205];
  wire _71853 = uncoded_block[1222] ^ uncoded_block[1255];
  wire _71854 = _71852 ^ _71853;
  wire _71855 = _71851 ^ _71854;
  wire _71856 = uncoded_block[1380] ^ uncoded_block[1420];
  wire _71857 = uncoded_block[1469] ^ uncoded_block[1530];
  wire _71858 = _71856 ^ _71857;
  wire _71859 = uncoded_block[1605] ^ uncoded_block[1639];
  wire _71860 = _71859 ^ uncoded_block[1654];
  wire _71861 = _71858 ^ _71860;
  wire _71862 = _71855 ^ _71861;
  wire _71863 = _71848 ^ _71862;
  wire _71864 = uncoded_block[7] ^ uncoded_block[54];
  wire _71865 = uncoded_block[148] ^ uncoded_block[205];
  wire _71866 = _71864 ^ _71865;
  wire _71867 = uncoded_block[233] ^ uncoded_block[305];
  wire _71868 = uncoded_block[369] ^ uncoded_block[398];
  wire _71869 = _71867 ^ _71868;
  wire _71870 = _71866 ^ _71869;
  wire _71871 = uncoded_block[497] ^ uncoded_block[513];
  wire _71872 = uncoded_block[577] ^ uncoded_block[652];
  wire _71873 = _71871 ^ _71872;
  wire _71874 = uncoded_block[669] ^ uncoded_block[755];
  wire _71875 = uncoded_block[788] ^ uncoded_block[882];
  wire _71876 = _71874 ^ _71875;
  wire _71877 = _71873 ^ _71876;
  wire _71878 = _71870 ^ _71877;
  wire _71879 = uncoded_block[896] ^ uncoded_block[999];
  wire _71880 = uncoded_block[1028] ^ uncoded_block[1060];
  wire _71881 = _71879 ^ _71880;
  wire _71882 = uncoded_block[1094] ^ uncoded_block[1157];
  wire _71883 = _71882 ^ _66819;
  wire _71884 = _71881 ^ _71883;
  wire _71885 = uncoded_block[1473] ^ uncoded_block[1518];
  wire _71886 = uncoded_block[1524] ^ uncoded_block[1598];
  wire _71887 = _71885 ^ _71886;
  wire _71888 = uncoded_block[1640] ^ uncoded_block[1667];
  wire _71889 = _71888 ^ uncoded_block[1698];
  wire _71890 = _71887 ^ _71889;
  wire _71891 = _71884 ^ _71890;
  wire _71892 = _71878 ^ _71891;
  wire _71893 = uncoded_block[9] ^ uncoded_block[83];
  wire _71894 = uncoded_block[118] ^ uncoded_block[212];
  wire _71895 = _71893 ^ _71894;
  wire _71896 = uncoded_block[225] ^ uncoded_block[326];
  wire _71897 = uncoded_block[345] ^ uncoded_block[446];
  wire _71898 = _71896 ^ _71897;
  wire _71899 = _71895 ^ _71898;
  wire _71900 = uncoded_block[504] ^ uncoded_block[536];
  wire _71901 = uncoded_block[591] ^ uncoded_block[639];
  wire _71902 = _71900 ^ _71901;
  wire _71903 = uncoded_block[710] ^ uncoded_block[736];
  wire _71904 = uncoded_block[816] ^ uncoded_block[847];
  wire _71905 = _71903 ^ _71904;
  wire _71906 = _71902 ^ _71905;
  wire _71907 = _71899 ^ _71906;
  wire _71908 = uncoded_block[909] ^ uncoded_block[977];
  wire _71909 = uncoded_block[1107] ^ uncoded_block[1136];
  wire _71910 = _71908 ^ _71909;
  wire _71911 = uncoded_block[1261] ^ uncoded_block[1294];
  wire _71912 = _67134 ^ _71911;
  wire _71913 = _71910 ^ _71912;
  wire _71914 = uncoded_block[1341] ^ uncoded_block[1439];
  wire _71915 = _71914 ^ _65987;
  wire _71916 = uncoded_block[1505] ^ uncoded_block[1628];
  wire _71917 = _71916 ^ uncoded_block[1704];
  wire _71918 = _71915 ^ _71917;
  wire _71919 = _71913 ^ _71918;
  wire _71920 = _71907 ^ _71919;
  wire _71921 = uncoded_block[11] ^ uncoded_block[105];
  wire _71922 = uncoded_block[115] ^ uncoded_block[181];
  wire _71923 = _71921 ^ _71922;
  wire _71924 = uncoded_block[238] ^ uncoded_block[296];
  wire _71925 = uncoded_block[385] ^ uncoded_block[418];
  wire _71926 = _71924 ^ _71925;
  wire _71927 = _71923 ^ _71926;
  wire _71928 = uncoded_block[500] ^ uncoded_block[508];
  wire _71929 = uncoded_block[583] ^ uncoded_block[643];
  wire _71930 = _71928 ^ _71929;
  wire _71931 = uncoded_block[689] ^ uncoded_block[730];
  wire _71932 = uncoded_block[826] ^ uncoded_block[839];
  wire _71933 = _71931 ^ _71932;
  wire _71934 = _71930 ^ _71933;
  wire _71935 = _71927 ^ _71934;
  wire _71936 = uncoded_block[893] ^ uncoded_block[950];
  wire _71937 = uncoded_block[1029] ^ uncoded_block[1108];
  wire _71938 = _71936 ^ _71937;
  wire _71939 = uncoded_block[1147] ^ uncoded_block[1184];
  wire _71940 = uncoded_block[1299] ^ uncoded_block[1376];
  wire _71941 = _71939 ^ _71940;
  wire _71942 = _71938 ^ _71941;
  wire _71943 = uncoded_block[1471] ^ uncoded_block[1523];
  wire _71944 = uncoded_block[1548] ^ uncoded_block[1595];
  wire _71945 = _71943 ^ _71944;
  wire _71946 = uncoded_block[1644] ^ uncoded_block[1683];
  wire _71947 = _71946 ^ uncoded_block[1717];
  wire _71948 = _71945 ^ _71947;
  wire _71949 = _71942 ^ _71948;
  wire _71950 = _71935 ^ _71949;
  wire _71951 = uncoded_block[14] ^ uncoded_block[86];
  wire _71952 = _71951 ^ _70240;
  wire _71953 = uncoded_block[267] ^ uncoded_block[317];
  wire _71954 = _71953 ^ _56452;
  wire _71955 = _71952 ^ _71954;
  wire _71956 = uncoded_block[464] ^ uncoded_block[530];
  wire _71957 = _71956 ^ _70254;
  wire _71958 = uncoded_block[769] ^ uncoded_block[811];
  wire _71959 = uncoded_block[832] ^ uncoded_block[939];
  wire _71960 = _71958 ^ _71959;
  wire _71961 = _71957 ^ _71960;
  wire _71962 = _71955 ^ _71961;
  wire _71963 = uncoded_block[970] ^ uncoded_block[1043];
  wire _71964 = uncoded_block[1080] ^ uncoded_block[1149];
  wire _71965 = _71963 ^ _71964;
  wire _71966 = uncoded_block[1204] ^ uncoded_block[1274];
  wire _71967 = uncoded_block[1312] ^ uncoded_block[1454];
  wire _71968 = _71966 ^ _71967;
  wire _71969 = _71965 ^ _71968;
  wire _71970 = _57765 ^ _21338;
  wire _71971 = uncoded_block[1533] ^ uncoded_block[1663];
  wire _71972 = _71971 ^ uncoded_block[1714];
  wire _71973 = _71970 ^ _71972;
  wire _71974 = _71969 ^ _71973;
  wire _71975 = _71962 ^ _71974;
  wire _71976 = uncoded_block[15] ^ uncoded_block[93];
  wire _71977 = uncoded_block[151] ^ uncoded_block[200];
  wire _71978 = _71976 ^ _71977;
  wire _71979 = uncoded_block[265] ^ uncoded_block[284];
  wire _71980 = uncoded_block[354] ^ uncoded_block[410];
  wire _71981 = _71979 ^ _71980;
  wire _71982 = _71978 ^ _71981;
  wire _71983 = uncoded_block[488] ^ uncoded_block[525];
  wire _71984 = uncoded_block[614] ^ uncoded_block[642];
  wire _71985 = _71983 ^ _71984;
  wire _71986 = uncoded_block[706] ^ uncoded_block[802];
  wire _71987 = uncoded_block[852] ^ uncoded_block[888];
  wire _71988 = _71986 ^ _71987;
  wire _71989 = _71985 ^ _71988;
  wire _71990 = _71982 ^ _71989;
  wire _71991 = uncoded_block[956] ^ uncoded_block[1022];
  wire _71992 = uncoded_block[1062] ^ uncoded_block[1131];
  wire _71993 = _71991 ^ _71992;
  wire _71994 = uncoded_block[1197] ^ uncoded_block[1236];
  wire _71995 = uncoded_block[1326] ^ uncoded_block[1366];
  wire _71996 = _71994 ^ _71995;
  wire _71997 = _71993 ^ _71996;
  wire _71998 = uncoded_block[1538] ^ uncoded_block[1553];
  wire _71999 = uncoded_block[1573] ^ uncoded_block[1604];
  wire _72000 = _71998 ^ _71999;
  wire _72001 = uncoded_block[1642] ^ uncoded_block[1650];
  wire _72002 = _72001 ^ uncoded_block[1712];
  wire _72003 = _72000 ^ _72002;
  wire _72004 = _71997 ^ _72003;
  wire _72005 = _71990 ^ _72004;
  wire _72006 = uncoded_block[19] ^ uncoded_block[76];
  wire _72007 = uncoded_block[126] ^ uncoded_block[198];
  wire _72008 = _72006 ^ _72007;
  wire _72009 = _49516 ^ _67184;
  wire _72010 = _72008 ^ _72009;
  wire _72011 = uncoded_block[467] ^ uncoded_block[540];
  wire _72012 = _72011 ^ _67197;
  wire _72013 = uncoded_block[715] ^ uncoded_block[750];
  wire _72014 = uncoded_block[793] ^ uncoded_block[834];
  wire _72015 = _72013 ^ _72014;
  wire _72016 = _72012 ^ _72015;
  wire _72017 = _72010 ^ _72016;
  wire _72018 = uncoded_block[925] ^ uncoded_block[968];
  wire _72019 = uncoded_block[1026] ^ uncoded_block[1096];
  wire _72020 = _72018 ^ _72019;
  wire _72021 = uncoded_block[1140] ^ uncoded_block[1238];
  wire _72022 = uncoded_block[1290] ^ uncoded_block[1355];
  wire _72023 = _72021 ^ _72022;
  wire _72024 = _72020 ^ _72023;
  wire _72025 = uncoded_block[1395] ^ uncoded_block[1558];
  wire _72026 = _72025 ^ _67232;
  wire _72027 = _67554 ^ uncoded_block[1691];
  wire _72028 = _72026 ^ _72027;
  wire _72029 = _72024 ^ _72028;
  wire _72030 = _72017 ^ _72029;
  wire _72031 = uncoded_block[21] ^ uncoded_block[65];
  wire _72032 = uncoded_block[142] ^ uncoded_block[180];
  wire _72033 = _72031 ^ _72032;
  wire _72034 = uncoded_block[260] ^ uncoded_block[316];
  wire _72035 = uncoded_block[370] ^ uncoded_block[419];
  wire _72036 = _72034 ^ _72035;
  wire _72037 = _72033 ^ _72036;
  wire _72038 = uncoded_block[456] ^ uncoded_block[557];
  wire _72039 = uncoded_block[595] ^ uncoded_block[636];
  wire _72040 = _72038 ^ _72039;
  wire _72041 = uncoded_block[693] ^ uncoded_block[748];
  wire _72042 = uncoded_block[809] ^ uncoded_block[876];
  wire _72043 = _72041 ^ _72042;
  wire _72044 = _72040 ^ _72043;
  wire _72045 = _72037 ^ _72044;
  wire _72046 = uncoded_block[900] ^ uncoded_block[988];
  wire _72047 = uncoded_block[1020] ^ uncoded_block[1077];
  wire _72048 = _72046 ^ _72047;
  wire _72049 = uncoded_block[1125] ^ uncoded_block[1199];
  wire _72050 = uncoded_block[1229] ^ uncoded_block[1324];
  wire _72051 = _72049 ^ _72050;
  wire _72052 = _72048 ^ _72051;
  wire _72053 = uncoded_block[1368] ^ uncoded_block[1406];
  wire _72054 = uncoded_block[1447] ^ uncoded_block[1575];
  wire _72055 = _72053 ^ _72054;
  wire _72056 = uncoded_block[1596] ^ uncoded_block[1633];
  wire _72057 = _72056 ^ uncoded_block[1665];
  wire _72058 = _72055 ^ _72057;
  wire _72059 = _72052 ^ _72058;
  wire _72060 = _72045 ^ _72059;
  wire _72061 = uncoded_block[23] ^ uncoded_block[63];
  wire _72062 = uncoded_block[134] ^ uncoded_block[190];
  wire _72063 = _72061 ^ _72062;
  wire _72064 = uncoded_block[234] ^ uncoded_block[303];
  wire _72065 = uncoded_block[352] ^ uncoded_block[443];
  wire _72066 = _72064 ^ _72065;
  wire _72067 = _72063 ^ _72066;
  wire _72068 = uncoded_block[460] ^ uncoded_block[547];
  wire _72069 = _72068 ^ _65368;
  wire _72070 = uncoded_block[678] ^ uncoded_block[732];
  wire _72071 = uncoded_block[814] ^ uncoded_block[875];
  wire _72072 = _72070 ^ _72071;
  wire _72073 = _72069 ^ _72072;
  wire _72074 = _72067 ^ _72073;
  wire _72075 = uncoded_block[932] ^ uncoded_block[995];
  wire _72076 = uncoded_block[1031] ^ uncoded_block[1145];
  wire _72077 = _72075 ^ _72076;
  wire _72078 = uncoded_block[1176] ^ uncoded_block[1250];
  wire _72079 = uncoded_block[1444] ^ uncoded_block[1487];
  wire _72080 = _72078 ^ _72079;
  wire _72081 = _72077 ^ _72080;
  wire _72082 = uncoded_block[1535] ^ uncoded_block[1552];
  wire _72083 = _65406 ^ _72082;
  wire _72084 = uncoded_block[1566] ^ uncoded_block[1623];
  wire _72085 = _72084 ^ uncoded_block[1684];
  wire _72086 = _72083 ^ _72085;
  wire _72087 = _72081 ^ _72086;
  wire _72088 = _72074 ^ _72087;
  wire _72089 = uncoded_block[25] ^ uncoded_block[78];
  wire _72090 = uncoded_block[164] ^ uncoded_block[224];
  wire _72091 = _72089 ^ _72090;
  wire _72092 = uncoded_block[231] ^ uncoded_block[311];
  wire _72093 = uncoded_block[340] ^ uncoded_block[413];
  wire _72094 = _72092 ^ _72093;
  wire _72095 = _72091 ^ _72094;
  wire _72096 = uncoded_block[471] ^ uncoded_block[545];
  wire _72097 = uncoded_block[581] ^ uncoded_block[647];
  wire _72098 = _72096 ^ _72097;
  wire _72099 = uncoded_block[698] ^ uncoded_block[765];
  wire _72100 = uncoded_block[790] ^ uncoded_block[848];
  wire _72101 = _72099 ^ _72100;
  wire _72102 = _72098 ^ _72101;
  wire _72103 = _72095 ^ _72102;
  wire _72104 = uncoded_block[919] ^ uncoded_block[967];
  wire _72105 = uncoded_block[1013] ^ uncoded_block[1064];
  wire _72106 = _72104 ^ _72105;
  wire _72107 = uncoded_block[1138] ^ uncoded_block[1209];
  wire _72108 = uncoded_block[1219] ^ uncoded_block[1266];
  wire _72109 = _72107 ^ _72108;
  wire _72110 = _72106 ^ _72109;
  wire _72111 = uncoded_block[1327] ^ uncoded_block[1408];
  wire _72112 = uncoded_block[1456] ^ uncoded_block[1579];
  wire _72113 = _72111 ^ _72112;
  wire _72114 = uncoded_block[1622] ^ uncoded_block[1661];
  wire _72115 = _72114 ^ uncoded_block[1715];
  wire _72116 = _72113 ^ _72115;
  wire _72117 = _72110 ^ _72116;
  wire _72118 = _72103 ^ _72117;
  wire _72119 = uncoded_block[26] ^ uncoded_block[103];
  wire _72120 = uncoded_block[145] ^ uncoded_block[195];
  wire _72121 = _72119 ^ _72120;
  wire _72122 = uncoded_block[242] ^ uncoded_block[324];
  wire _72123 = uncoded_block[378] ^ uncoded_block[432];
  wire _72124 = _72122 ^ _72123;
  wire _72125 = _72121 ^ _72124;
  wire _72126 = uncoded_block[489] ^ uncoded_block[516];
  wire _72127 = uncoded_block[613] ^ uncoded_block[646];
  wire _72128 = _72126 ^ _72127;
  wire _72129 = uncoded_block[786] ^ uncoded_block[831];
  wire _72130 = _68137 ^ _72129;
  wire _72131 = _72128 ^ _72130;
  wire _72132 = _72125 ^ _72131;
  wire _72133 = uncoded_block[984] ^ uncoded_block[1030];
  wire _72134 = _68146 ^ _72133;
  wire _72135 = uncoded_block[1070] ^ uncoded_block[1123];
  wire _72136 = uncoded_block[1191] ^ uncoded_block[1270];
  wire _72137 = _72135 ^ _72136;
  wire _72138 = _72134 ^ _72137;
  wire _72139 = uncoded_block[1298] ^ uncoded_block[1369];
  wire _72140 = uncoded_block[1385] ^ uncoded_block[1478];
  wire _72141 = _72139 ^ _72140;
  wire _72142 = uncoded_block[1613] ^ uncoded_block[1687];
  wire _72143 = _72142 ^ uncoded_block[1697];
  wire _72144 = _72141 ^ _72143;
  wire _72145 = _72138 ^ _72144;
  wire _72146 = _72132 ^ _72145;
  wire _72147 = uncoded_block[40] ^ uncoded_block[84];
  wire _72148 = _72147 ^ _66423;
  wire _72149 = uncoded_block[374] ^ uncoded_block[391];
  wire _72150 = _66989 ^ _72149;
  wire _72151 = _72148 ^ _72150;
  wire _72152 = uncoded_block[395] ^ uncoded_block[496];
  wire _72153 = uncoded_block[544] ^ uncoded_block[590];
  wire _72154 = _72152 ^ _72153;
  wire _72155 = uncoded_block[772] ^ uncoded_block[827];
  wire _72156 = _67006 ^ _72155;
  wire _72157 = _72154 ^ _72156;
  wire _72158 = _72151 ^ _72157;
  wire _72159 = uncoded_block[863] ^ uncoded_block[913];
  wire _72160 = uncoded_block[965] ^ uncoded_block[1009];
  wire _72161 = _72159 ^ _72160;
  wire _72162 = uncoded_block[1076] ^ uncoded_block[1146];
  wire _72163 = uncoded_block[1200] ^ uncoded_block[1253];
  wire _72164 = _72162 ^ _72163;
  wire _72165 = _72161 ^ _72164;
  wire _72166 = uncoded_block[1300] ^ uncoded_block[1361];
  wire _72167 = uncoded_block[1392] ^ uncoded_block[1437];
  wire _72168 = _72166 ^ _72167;
  wire _72169 = uncoded_block[1593] ^ uncoded_block[1616];
  wire _72170 = _72169 ^ uncoded_block[1680];
  wire _72171 = _72168 ^ _72170;
  wire _72172 = _72165 ^ _72171;
  wire _72173 = _72158 ^ _72172;
  wire _72174 = uncoded_block[41] ^ uncoded_block[106];
  wire _72175 = uncoded_block[124] ^ uncoded_block[174];
  wire _72176 = _72174 ^ _72175;
  wire _72177 = uncoded_block[270] ^ uncoded_block[332];
  wire _72178 = uncoded_block[348] ^ uncoded_block[408];
  wire _72179 = _72177 ^ _72178;
  wire _72180 = _72176 ^ _72179;
  wire _72181 = _65494 ^ _65501;
  wire _72182 = uncoded_block[699] ^ uncoded_block[761];
  wire _72183 = _72182 ^ _65509;
  wire _72184 = _72181 ^ _72183;
  wire _72185 = _72180 ^ _72184;
  wire _72186 = uncoded_block[912] ^ uncoded_block[997];
  wire _72187 = uncoded_block[1041] ^ uncoded_block[1086];
  wire _72188 = _72186 ^ _72187;
  wire _72189 = uncoded_block[1143] ^ uncoded_block[1188];
  wire _72190 = uncoded_block[1257] ^ uncoded_block[1286];
  wire _72191 = _72189 ^ _72190;
  wire _72192 = _72188 ^ _72191;
  wire _72193 = uncoded_block[1365] ^ uncoded_block[1460];
  wire _72194 = uncoded_block[1475] ^ uncoded_block[1547];
  wire _72195 = _72193 ^ _72194;
  wire _72196 = uncoded_block[1609] ^ uncoded_block[1653];
  wire _72197 = _72196 ^ uncoded_block[1694];
  wire _72198 = _72195 ^ _72197;
  wire _72199 = _72192 ^ _72198;
  wire _72200 = _72185 ^ _72199;
  wire _72201 = uncoded_block[49] ^ uncoded_block[112];
  wire _72202 = uncoded_block[210] ^ uncoded_block[256];
  wire _72203 = _72201 ^ _72202;
  wire _72204 = uncoded_block[318] ^ uncoded_block[381];
  wire _72205 = uncoded_block[417] ^ uncoded_block[485];
  wire _72206 = _72204 ^ _72205;
  wire _72207 = _72203 ^ _72206;
  wire _72208 = uncoded_block[528] ^ uncoded_block[601];
  wire _72209 = uncoded_block[627] ^ uncoded_block[694];
  wire _72210 = _72208 ^ _72209;
  wire _72211 = uncoded_block[741] ^ uncoded_block[791];
  wire _72212 = uncoded_block[861] ^ uncoded_block[897];
  wire _72213 = _72211 ^ _72212;
  wire _72214 = _72210 ^ _72213;
  wire _72215 = _72207 ^ _72214;
  wire _72216 = uncoded_block[979] ^ uncoded_block[1148];
  wire _72217 = uncoded_block[1195] ^ uncoded_block[1260];
  wire _72218 = _72216 ^ _72217;
  wire _72219 = uncoded_block[1350] ^ uncoded_block[1424];
  wire _72220 = uncoded_block[1442] ^ uncoded_block[1485];
  wire _72221 = _72219 ^ _72220;
  wire _72222 = _72218 ^ _72221;
  wire _72223 = uncoded_block[1529] ^ uncoded_block[1556];
  wire _72224 = _23190 ^ _72223;
  wire _72225 = uncoded_block[1578] ^ uncoded_block[1676];
  wire _72226 = _72225 ^ uncoded_block[1690];
  wire _72227 = _72224 ^ _72226;
  wire _72228 = _72222 ^ _72227;
  wire _72229 = _72215 ^ _72228;
  wire _72230 = uncoded_block[1] ^ uncoded_block[100];
  wire _72231 = uncoded_block[148] ^ uncoded_block[178];
  wire _72232 = _72230 ^ _72231;
  wire _72233 = uncoded_block[248] ^ uncoded_block[315];
  wire _72234 = uncoded_block[365] ^ uncoded_block[416];
  wire _72235 = _72233 ^ _72234;
  wire _72236 = _72232 ^ _72235;
  wire _72237 = uncoded_block[483] ^ uncoded_block[522];
  wire _72238 = uncoded_block[607] ^ uncoded_block[624];
  wire _72239 = _72237 ^ _72238;
  wire _72240 = uncoded_block[697] ^ uncoded_block[769];
  wire _72241 = uncoded_block[804] ^ uncoded_block[861];
  wire _72242 = _72240 ^ _72241;
  wire _72243 = _72239 ^ _72242;
  wire _72244 = _72236 ^ _72243;
  wire _72245 = uncoded_block[934] ^ uncoded_block[998];
  wire _72246 = uncoded_block[1030] ^ uncoded_block[1083];
  wire _72247 = _72245 ^ _72246;
  wire _72248 = uncoded_block[1209] ^ uncoded_block[1231];
  wire _72249 = _67530 ^ _72248;
  wire _72250 = _72247 ^ _72249;
  wire _72251 = uncoded_block[1299] ^ uncoded_block[1338];
  wire _72252 = uncoded_block[1395] ^ uncoded_block[1474];
  wire _72253 = _72251 ^ _72252;
  wire _72254 = uncoded_block[1494] ^ uncoded_block[1591];
  wire _72255 = _72254 ^ uncoded_block[1710];
  wire _72256 = _72253 ^ _72255;
  wire _72257 = _72250 ^ _72256;
  wire _72258 = _72244 ^ _72257;
  wire _72259 = uncoded_block[6] ^ uncoded_block[105];
  wire _72260 = uncoded_block[153] ^ uncoded_block[184];
  wire _72261 = _72259 ^ _72260;
  wire _72262 = uncoded_block[252] ^ uncoded_block[321];
  wire _72263 = uncoded_block[371] ^ uncoded_block[422];
  wire _72264 = _72262 ^ _72263;
  wire _72265 = _72261 ^ _72264;
  wire _72266 = uncoded_block[487] ^ uncoded_block[527];
  wire _72267 = uncoded_block[612] ^ uncoded_block[628];
  wire _72268 = _72266 ^ _72267;
  wire _72269 = uncoded_block[703] ^ uncoded_block[774];
  wire _72270 = uncoded_block[809] ^ uncoded_block[866];
  wire _72271 = _72269 ^ _72270;
  wire _72272 = _72268 ^ _72271;
  wire _72273 = _72265 ^ _72272;
  wire _72274 = uncoded_block[1035] ^ uncoded_block[1088];
  wire _72275 = _1300 ^ _72274;
  wire _72276 = uncoded_block[1152] ^ uncoded_block[1214];
  wire _72277 = _72276 ^ _62416;
  wire _72278 = _72275 ^ _72277;
  wire _72279 = uncoded_block[1303] ^ uncoded_block[1344];
  wire _72280 = uncoded_block[1400] ^ uncoded_block[1561];
  wire _72281 = _72279 ^ _72280;
  wire _72282 = uncoded_block[1594] ^ uncoded_block[1611];
  wire _72283 = _72282 ^ uncoded_block[1651];
  wire _72284 = _72281 ^ _72283;
  wire _72285 = _72278 ^ _72284;
  wire _72286 = _72273 ^ _72285;
  wire _72287 = uncoded_block[11] ^ uncoded_block[108];
  wire _72288 = uncoded_block[158] ^ uncoded_block[187];
  wire _72289 = _72287 ^ _72288;
  wire _72290 = uncoded_block[256] ^ uncoded_block[325];
  wire _72291 = uncoded_block[376] ^ uncoded_block[426];
  wire _72292 = _72290 ^ _72291;
  wire _72293 = _72289 ^ _72292;
  wire _72294 = uncoded_block[492] ^ uncoded_block[532];
  wire _72295 = uncoded_block[562] ^ uncoded_block[631];
  wire _72296 = _72294 ^ _72295;
  wire _72297 = uncoded_block[707] ^ uncoded_block[724];
  wire _72298 = uncoded_block[814] ^ uncoded_block[869];
  wire _72299 = _72297 ^ _72298;
  wire _72300 = _72296 ^ _72299;
  wire _72301 = _72293 ^ _72300;
  wire _72302 = uncoded_block[888] ^ uncoded_block[949];
  wire _72303 = uncoded_block[1040] ^ uncoded_block[1091];
  wire _72304 = _72302 ^ _72303;
  wire _72305 = uncoded_block[1156] ^ uncoded_block[1217];
  wire _72306 = uncoded_block[1240] ^ uncoded_block[1276];
  wire _72307 = _72305 ^ _72306;
  wire _72308 = _72304 ^ _72307;
  wire _72309 = uncoded_block[1306] ^ uncoded_block[1349];
  wire _72310 = uncoded_block[1405] ^ uncoded_block[1565];
  wire _72311 = _72309 ^ _72310;
  wire _72312 = uncoded_block[1598] ^ uncoded_block[1614];
  wire _72313 = _72312 ^ uncoded_block[1714];
  wire _72314 = _72311 ^ _72313;
  wire _72315 = _72308 ^ _72314;
  wire _72316 = _72301 ^ _72315;
  wire _72317 = uncoded_block[12] ^ uncoded_block[54];
  wire _72318 = uncoded_block[160] ^ uncoded_block[189];
  wire _72319 = _72317 ^ _72318;
  wire _72320 = uncoded_block[258] ^ uncoded_block[327];
  wire _72321 = uncoded_block[378] ^ uncoded_block[428];
  wire _72322 = _72320 ^ _72321;
  wire _72323 = _72319 ^ _72322;
  wire _72324 = uncoded_block[494] ^ uncoded_block[534];
  wire _72325 = uncoded_block[564] ^ uncoded_block[633];
  wire _72326 = _72324 ^ _72325;
  wire _72327 = uncoded_block[709] ^ uncoded_block[725];
  wire _72328 = uncoded_block[816] ^ uncoded_block[871];
  wire _72329 = _72327 ^ _72328;
  wire _72330 = _72326 ^ _72329;
  wire _72331 = _72323 ^ _72330;
  wire _72332 = uncoded_block[890] ^ uncoded_block[951];
  wire _72333 = uncoded_block[1042] ^ uncoded_block[1093];
  wire _72334 = _72332 ^ _72333;
  wire _72335 = uncoded_block[1158] ^ uncoded_block[1241];
  wire _72336 = uncoded_block[1308] ^ uncoded_block[1351];
  wire _72337 = _72335 ^ _72336;
  wire _72338 = _72334 ^ _72337;
  wire _72339 = uncoded_block[1407] ^ uncoded_block[1516];
  wire _72340 = _72339 ^ _68960;
  wire _72341 = uncoded_block[1616] ^ uncoded_block[1655];
  wire _72342 = _72341 ^ uncoded_block[1715];
  wire _72343 = _72340 ^ _72342;
  wire _72344 = _72338 ^ _72343;
  wire _72345 = _72331 ^ _72344;
  wire _72346 = uncoded_block[15] ^ uncoded_block[57];
  wire _72347 = uncoded_block[163] ^ uncoded_block[191];
  wire _72348 = _72346 ^ _72347;
  wire _72349 = uncoded_block[261] ^ uncoded_block[329];
  wire _72350 = uncoded_block[381] ^ uncoded_block[431];
  wire _72351 = _72349 ^ _72350;
  wire _72352 = _72348 ^ _72351;
  wire _72353 = uncoded_block[497] ^ uncoded_block[537];
  wire _72354 = uncoded_block[567] ^ uncoded_block[636];
  wire _72355 = _72353 ^ _72354;
  wire _72356 = uncoded_block[711] ^ uncoded_block[728];
  wire _72357 = uncoded_block[819] ^ uncoded_block[874];
  wire _72358 = _72356 ^ _72357;
  wire _72359 = _72355 ^ _72358;
  wire _72360 = _72352 ^ _72359;
  wire _72361 = uncoded_block[893] ^ uncoded_block[954];
  wire _72362 = uncoded_block[1045] ^ uncoded_block[1095];
  wire _72363 = _72361 ^ _72362;
  wire _72364 = uncoded_block[1161] ^ uncoded_block[1243];
  wire _72365 = uncoded_block[1280] ^ uncoded_block[1310];
  wire _72366 = _72364 ^ _72365;
  wire _72367 = _72363 ^ _72366;
  wire _72368 = uncoded_block[1354] ^ uncoded_block[1410];
  wire _72369 = uncoded_block[1517] ^ uncoded_block[1570];
  wire _72370 = _72368 ^ _72369;
  wire _72371 = uncoded_block[1602] ^ uncoded_block[1619];
  wire _72372 = _72371 ^ uncoded_block[1657];
  wire _72373 = _72370 ^ _72372;
  wire _72374 = _72367 ^ _72373;
  wire _72375 = _72360 ^ _72374;
  wire _72376 = uncoded_block[17] ^ uncoded_block[59];
  wire _72377 = uncoded_block[165] ^ uncoded_block[193];
  wire _72378 = _72376 ^ _72377;
  wire _72379 = uncoded_block[263] ^ uncoded_block[331];
  wire _72380 = uncoded_block[383] ^ uncoded_block[433];
  wire _72381 = _72379 ^ _72380;
  wire _72382 = _72378 ^ _72381;
  wire _72383 = uncoded_block[499] ^ uncoded_block[539];
  wire _72384 = uncoded_block[569] ^ uncoded_block[638];
  wire _72385 = _72383 ^ _72384;
  wire _72386 = uncoded_block[713] ^ uncoded_block[730];
  wire _72387 = uncoded_block[820] ^ uncoded_block[876];
  wire _72388 = _72386 ^ _72387;
  wire _72389 = _72385 ^ _72388;
  wire _72390 = _72382 ^ _72389;
  wire _72391 = uncoded_block[895] ^ uncoded_block[956];
  wire _72392 = uncoded_block[1047] ^ uncoded_block[1097];
  wire _72393 = _72391 ^ _72392;
  wire _72394 = uncoded_block[1163] ^ uncoded_block[1170];
  wire _72395 = uncoded_block[1245] ^ uncoded_block[1282];
  wire _72396 = _72394 ^ _72395;
  wire _72397 = _72393 ^ _72396;
  wire _72398 = uncoded_block[1312] ^ uncoded_block[1355];
  wire _72399 = uncoded_block[1572] ^ uncoded_block[1603];
  wire _72400 = _72398 ^ _72399;
  wire _72401 = uncoded_block[1621] ^ uncoded_block[1658];
  wire _72402 = _72401 ^ uncoded_block[1688];
  wire _72403 = _72400 ^ _72402;
  wire _72404 = _72397 ^ _72403;
  wire _72405 = _72390 ^ _72404;
  wire _72406 = uncoded_block[19] ^ uncoded_block[61];
  wire _72407 = uncoded_block[167] ^ uncoded_block[194];
  wire _72408 = _72406 ^ _72407;
  wire _72409 = uncoded_block[265] ^ uncoded_block[280];
  wire _72410 = uncoded_block[385] ^ uncoded_block[435];
  wire _72411 = _72409 ^ _72410;
  wire _72412 = _72408 ^ _72411;
  wire _72413 = uncoded_block[501] ^ uncoded_block[541];
  wire _72414 = uncoded_block[570] ^ uncoded_block[640];
  wire _72415 = _72413 ^ _72414;
  wire _72416 = uncoded_block[822] ^ uncoded_block[877];
  wire _72417 = _61308 ^ _72416;
  wire _72418 = _72415 ^ _72417;
  wire _72419 = _72412 ^ _72418;
  wire _72420 = uncoded_block[897] ^ uncoded_block[958];
  wire _72421 = uncoded_block[1049] ^ uncoded_block[1098];
  wire _72422 = _72420 ^ _72421;
  wire _72423 = uncoded_block[1172] ^ uncoded_block[1247];
  wire _72424 = _72423 ^ _61357;
  wire _72425 = _72422 ^ _72424;
  wire _72426 = uncoded_block[1357] ^ uncoded_block[1413];
  wire _72427 = uncoded_block[1510] ^ uncoded_block[1605];
  wire _72428 = _72426 ^ _72427;
  wire _72429 = uncoded_block[1623] ^ uncoded_block[1660];
  wire _72430 = _72429 ^ uncoded_block[1689];
  wire _72431 = _72428 ^ _72430;
  wire _72432 = _72425 ^ _72431;
  wire _72433 = _72419 ^ _72432;
  wire _72434 = uncoded_block[21] ^ uncoded_block[63];
  wire _72435 = uncoded_block[169] ^ uncoded_block[196];
  wire _72436 = _72434 ^ _72435;
  wire _72437 = uncoded_block[387] ^ uncoded_block[437];
  wire _72438 = _62475 ^ _72437;
  wire _72439 = _72436 ^ _72438;
  wire _72440 = uncoded_block[503] ^ uncoded_block[543];
  wire _72441 = uncoded_block[572] ^ uncoded_block[642];
  wire _72442 = _72440 ^ _72441;
  wire _72443 = uncoded_block[716] ^ uncoded_block[733];
  wire _72444 = uncoded_block[824] ^ uncoded_block[879];
  wire _72445 = _72443 ^ _72444;
  wire _72446 = _72442 ^ _72445;
  wire _72447 = _72439 ^ _72446;
  wire _72448 = uncoded_block[899] ^ uncoded_block[960];
  wire _72449 = uncoded_block[1051] ^ uncoded_block[1100];
  wire _72450 = _72448 ^ _72449;
  wire _72451 = uncoded_block[1174] ^ uncoded_block[1249];
  wire _72452 = _72451 ^ _67654;
  wire _72453 = _72450 ^ _72452;
  wire _72454 = uncoded_block[1358] ^ uncoded_block[1415];
  wire _72455 = uncoded_block[1458] ^ uncoded_block[1512];
  wire _72456 = _72454 ^ _72455;
  wire _72457 = _67664 ^ uncoded_block[1690];
  wire _72458 = _72456 ^ _72457;
  wire _72459 = _72453 ^ _72458;
  wire _72460 = _72447 ^ _72459;
  wire _72461 = uncoded_block[26] ^ uncoded_block[68];
  wire _72462 = uncoded_block[114] ^ uncoded_block[199];
  wire _72463 = _72461 ^ _72462;
  wire _72464 = uncoded_block[271] ^ uncoded_block[333];
  wire _72465 = uncoded_block[440] ^ uncoded_block[451];
  wire _72466 = _72464 ^ _72465;
  wire _72467 = _72463 ^ _72466;
  wire _72468 = uncoded_block[548] ^ uncoded_block[577];
  wire _72469 = uncoded_block[647] ^ uncoded_block[719];
  wire _72470 = _72468 ^ _72469;
  wire _72471 = uncoded_block[737] ^ uncoded_block[827];
  wire _72472 = uncoded_block[884] ^ uncoded_block[904];
  wire _72473 = _72471 ^ _72472;
  wire _72474 = _72470 ^ _72473;
  wire _72475 = _72467 ^ _72474;
  wire _72476 = uncoded_block[964] ^ uncoded_block[1056];
  wire _72477 = _72476 ^ _63680;
  wire _72478 = uncoded_block[1177] ^ uncoded_block[1254];
  wire _72479 = uncoded_block[1320] ^ uncoded_block[1363];
  wire _72480 = _72478 ^ _72479;
  wire _72481 = _72477 ^ _72480;
  wire _72482 = uncoded_block[1384] ^ uncoded_block[1419];
  wire _72483 = uncoded_block[1463] ^ uncoded_block[1556];
  wire _72484 = _72482 ^ _72483;
  wire _72485 = uncoded_block[1628] ^ uncoded_block[1664];
  wire _72486 = _72485 ^ uncoded_block[1693];
  wire _72487 = _72484 ^ _72486;
  wire _72488 = _72481 ^ _72487;
  wire _72489 = _72475 ^ _72488;
  wire _72490 = uncoded_block[28] ^ uncoded_block[70];
  wire _72491 = uncoded_block[116] ^ uncoded_block[201];
  wire _72492 = _72490 ^ _72491;
  wire _72493 = uncoded_block[334] ^ uncoded_block[442];
  wire _72494 = _66340 ^ _72493;
  wire _72495 = _72492 ^ _72494;
  wire _72496 = uncoded_block[453] ^ uncoded_block[550];
  wire _72497 = uncoded_block[578] ^ uncoded_block[649];
  wire _72498 = _72496 ^ _72497;
  wire _72499 = uncoded_block[829] ^ uncoded_block[886];
  wire _72500 = _66028 ^ _72499;
  wire _72501 = _72498 ^ _72500;
  wire _72502 = _72495 ^ _72501;
  wire _72503 = uncoded_block[906] ^ uncoded_block[966];
  wire _72504 = uncoded_block[1058] ^ uncoded_block[1106];
  wire _72505 = _72503 ^ _72504;
  wire _72506 = uncoded_block[1115] ^ uncoded_block[1179];
  wire _72507 = uncoded_block[1255] ^ uncoded_block[1322];
  wire _72508 = _72506 ^ _72507;
  wire _72509 = _72505 ^ _72508;
  wire _72510 = uncoded_block[1364] ^ uncoded_block[1386];
  wire _72511 = uncoded_block[1421] ^ uncoded_block[1465];
  wire _72512 = _72510 ^ _72511;
  wire _72513 = uncoded_block[1558] ^ uncoded_block[1666];
  wire _72514 = _72513 ^ uncoded_block[1694];
  wire _72515 = _72512 ^ _72514;
  wire _72516 = _72509 ^ _72515;
  wire _72517 = _72502 ^ _72516;
  wire _72518 = uncoded_block[36] ^ uncoded_block[78];
  wire _72519 = uncoded_block[123] ^ uncoded_block[207];
  wire _72520 = _72518 ^ _72519;
  wire _72521 = uncoded_block[225] ^ uncoded_block[293];
  wire _72522 = uncoded_block[341] ^ uncoded_block[393];
  wire _72523 = _72521 ^ _72522;
  wire _72524 = _72520 ^ _72523;
  wire _72525 = uncoded_block[461] ^ uncoded_block[557];
  wire _72526 = uncoded_block[585] ^ uncoded_block[654];
  wire _72527 = _72525 ^ _72526;
  wire _72528 = uncoded_block[674] ^ uncoded_block[746];
  wire _72529 = _72528 ^ _65443;
  wire _72530 = _72527 ^ _72529;
  wire _72531 = _72524 ^ _72530;
  wire _72532 = uncoded_block[1008] ^ uncoded_block[1061];
  wire _72533 = _65514 ^ _72532;
  wire _72534 = uncoded_block[1122] ^ uncoded_block[1186];
  wire _72535 = uncoded_block[1262] ^ uncoded_block[1371];
  wire _72536 = _72534 ^ _72535;
  wire _72537 = _72533 ^ _72536;
  wire _72538 = uncoded_block[1428] ^ uncoded_block[1448];
  wire _72539 = uncoded_block[1480] ^ uncoded_block[1527];
  wire _72540 = _72538 ^ _72539;
  wire _72541 = uncoded_block[1537] ^ uncoded_block[1635];
  wire _72542 = _72541 ^ uncoded_block[1698];
  wire _72543 = _72540 ^ _72542;
  wire _72544 = _72537 ^ _72543;
  wire _72545 = _72531 ^ _72544;
  wire _72546 = uncoded_block[41] ^ uncoded_block[83];
  wire _72547 = uncoded_block[129] ^ uncoded_block[213];
  wire _72548 = _72546 ^ _72547;
  wire _72549 = uncoded_block[231] ^ uncoded_block[299];
  wire _72550 = uncoded_block[347] ^ uncoded_block[399];
  wire _72551 = _72549 ^ _72550;
  wire _72552 = _72548 ^ _72551;
  wire _72553 = uncoded_block[590] ^ uncoded_block[660];
  wire _72554 = _67737 ^ _72553;
  wire _72555 = uncoded_block[679] ^ uncoded_block[751];
  wire _72556 = uncoded_block[788] ^ uncoded_block[843];
  wire _72557 = _72555 ^ _72556;
  wire _72558 = _72554 ^ _72557;
  wire _72559 = _72552 ^ _72558;
  wire _72560 = uncoded_block[918] ^ uncoded_block[980];
  wire _72561 = uncoded_block[1067] ^ uncoded_block[1128];
  wire _72562 = _72560 ^ _72561;
  wire _72563 = uncoded_block[1192] ^ uncoded_block[1268];
  wire _72564 = uncoded_block[1284] ^ uncoded_block[1377];
  wire _72565 = _72563 ^ _72564;
  wire _72566 = _72562 ^ _72565;
  wire _72567 = uncoded_block[1433] ^ uncoded_block[1453];
  wire _72568 = _72567 ^ _67770;
  wire _72569 = uncoded_block[1639] ^ uncoded_block[1672];
  wire _72570 = _72569 ^ uncoded_block[1703];
  wire _72571 = _72568 ^ _72570;
  wire _72572 = _72566 ^ _72571;
  wire _72573 = _72559 ^ _72572;
  wire _72574 = uncoded_block[44] ^ uncoded_block[86];
  wire _72575 = uncoded_block[132] ^ uncoded_block[215];
  wire _72576 = _72574 ^ _72575;
  wire _72577 = uncoded_block[234] ^ uncoded_block[300];
  wire _72578 = uncoded_block[350] ^ uncoded_block[391];
  wire _72579 = _72577 ^ _72578;
  wire _72580 = _72576 ^ _72579;
  wire _72581 = uncoded_block[401] ^ uncoded_block[468];
  wire _72582 = uncoded_block[509] ^ uncoded_block[592];
  wire _72583 = _72581 ^ _72582;
  wire _72584 = uncoded_block[754] ^ uncoded_block[791];
  wire _72585 = _66930 ^ _72584;
  wire _72586 = _72583 ^ _72585;
  wire _72587 = _72580 ^ _72586;
  wire _72588 = uncoded_block[846] ^ uncoded_block[921];
  wire _72589 = uncoded_block[982] ^ uncoded_block[1016];
  wire _72590 = _72588 ^ _72589;
  wire _72591 = uncoded_block[1069] ^ uncoded_block[1130];
  wire _72592 = uncoded_block[1193] ^ uncoded_block[1271];
  wire _72593 = _72591 ^ _72592;
  wire _72594 = _72590 ^ _72593;
  wire _72595 = uncoded_block[1285] ^ uncoded_block[1379];
  wire _72596 = uncoded_block[1435] ^ uncoded_block[1543];
  wire _72597 = _72595 ^ _72596;
  wire _72598 = uncoded_block[1579] ^ uncoded_block[1642];
  wire _72599 = _72598 ^ uncoded_block[1675];
  wire _72600 = _72597 ^ _72599;
  wire _72601 = _72594 ^ _72600;
  wire _72602 = _72587 ^ _72601;
  wire _72603 = uncoded_block[46] ^ uncoded_block[87];
  wire _72604 = uncoded_block[134] ^ uncoded_block[217];
  wire _72605 = _72603 ^ _72604;
  wire _72606 = uncoded_block[235] ^ uncoded_block[301];
  wire _72607 = uncoded_block[351] ^ uncoded_block[403];
  wire _72608 = _72606 ^ _72607;
  wire _72609 = _72605 ^ _72608;
  wire _72610 = uncoded_block[470] ^ uncoded_block[510];
  wire _72611 = uncoded_block[594] ^ uncoded_block[664];
  wire _72612 = _72610 ^ _72611;
  wire _72613 = uncoded_block[683] ^ uncoded_block[722];
  wire _72614 = uncoded_block[756] ^ uncoded_block[792];
  wire _72615 = _72613 ^ _72614;
  wire _72616 = _72612 ^ _72615;
  wire _72617 = _72609 ^ _72616;
  wire _72618 = uncoded_block[848] ^ uncoded_block[922];
  wire _72619 = uncoded_block[984] ^ uncoded_block[1018];
  wire _72620 = _72618 ^ _72619;
  wire _72621 = uncoded_block[1071] ^ uncoded_block[1132];
  wire _72622 = uncoded_block[1195] ^ uncoded_block[1273];
  wire _72623 = _72621 ^ _72622;
  wire _72624 = _72620 ^ _72623;
  wire _72625 = uncoded_block[1286] ^ uncoded_block[1381];
  wire _72626 = uncoded_block[1437] ^ uncoded_block[1545];
  wire _72627 = _72625 ^ _72626;
  wire _72628 = uncoded_block[1580] ^ uncoded_block[1677];
  wire _72629 = _72628 ^ uncoded_block[1705];
  wire _72630 = _72627 ^ _72629;
  wire _72631 = _72624 ^ _72630;
  wire _72632 = _72617 ^ _72631;
  wire _72633 = uncoded_block[47] ^ uncoded_block[88];
  wire _72634 = uncoded_block[135] ^ uncoded_block[218];
  wire _72635 = _72633 ^ _72634;
  wire _72636 = uncoded_block[236] ^ uncoded_block[302];
  wire _72637 = uncoded_block[352] ^ uncoded_block[404];
  wire _72638 = _72636 ^ _72637;
  wire _72639 = _72635 ^ _72638;
  wire _72640 = uncoded_block[471] ^ uncoded_block[511];
  wire _72641 = uncoded_block[595] ^ uncoded_block[665];
  wire _72642 = _72640 ^ _72641;
  wire _72643 = uncoded_block[684] ^ uncoded_block[757];
  wire _72644 = _72643 ^ _67878;
  wire _72645 = _72642 ^ _72644;
  wire _72646 = _72639 ^ _72645;
  wire _72647 = uncoded_block[849] ^ uncoded_block[923];
  wire _72648 = _72647 ^ _67887;
  wire _72649 = uncoded_block[1072] ^ uncoded_block[1133];
  wire _72650 = uncoded_block[1196] ^ uncoded_block[1274];
  wire _72651 = _72649 ^ _72650;
  wire _72652 = _72648 ^ _72651;
  wire _72653 = uncoded_block[1287] ^ uncoded_block[1382];
  wire _72654 = uncoded_block[1438] ^ uncoded_block[1546];
  wire _72655 = _72653 ^ _72654;
  wire _72656 = uncoded_block[1581] ^ uncoded_block[1644];
  wire _72657 = _72656 ^ uncoded_block[1706];
  wire _72658 = _72655 ^ _72657;
  wire _72659 = _72652 ^ _72658;
  wire _72660 = _72646 ^ _72659;
  wire _72661 = uncoded_block[48] ^ uncoded_block[89];
  wire _72662 = uncoded_block[136] ^ uncoded_block[219];
  wire _72663 = _72661 ^ _72662;
  wire _72664 = uncoded_block[237] ^ uncoded_block[303];
  wire _72665 = uncoded_block[353] ^ uncoded_block[405];
  wire _72666 = _72664 ^ _72665;
  wire _72667 = _72663 ^ _72666;
  wire _72668 = uncoded_block[472] ^ uncoded_block[512];
  wire _72669 = uncoded_block[596] ^ uncoded_block[666];
  wire _72670 = _72668 ^ _72669;
  wire _72671 = uncoded_block[685] ^ uncoded_block[758];
  wire _72672 = uncoded_block[794] ^ uncoded_block[830];
  wire _72673 = _72671 ^ _72672;
  wire _72674 = _72670 ^ _72673;
  wire _72675 = _72667 ^ _72674;
  wire _72676 = uncoded_block[850] ^ uncoded_block[924];
  wire _72677 = uncoded_block[986] ^ uncoded_block[1020];
  wire _72678 = _72676 ^ _72677;
  wire _72679 = uncoded_block[1073] ^ uncoded_block[1134];
  wire _72680 = uncoded_block[1197] ^ uncoded_block[1275];
  wire _72681 = _72679 ^ _72680;
  wire _72682 = _72678 ^ _72681;
  wire _72683 = uncoded_block[1288] ^ uncoded_block[1383];
  wire _72684 = uncoded_block[1439] ^ uncoded_block[1547];
  wire _72685 = _72683 ^ _72684;
  wire _72686 = uncoded_block[1582] ^ uncoded_block[1645];
  wire _72687 = _72686 ^ uncoded_block[1678];
  wire _72688 = _72685 ^ _72687;
  wire _72689 = _72682 ^ _72688;
  wire _72690 = _72675 ^ _72689;
  wire _72691 = uncoded_block[53] ^ uncoded_block[110];
  wire _72692 = uncoded_block[170] ^ uncoded_block[224];
  wire _72693 = _72691 ^ _72692;
  wire _72694 = uncoded_block[279] ^ uncoded_block[332];
  wire _72695 = uncoded_block[447] ^ uncoded_block[505];
  wire _72696 = _72694 ^ _72695;
  wire _72697 = _72693 ^ _72696;
  wire _72698 = uncoded_block[616] ^ uncoded_block[668];
  wire _72699 = _72698 ^ _743;
  wire _72700 = _72699 ^ _45099;
  wire _72701 = _72697 ^ _72700;
  wire _72702 = _4614 ^ _66111;
  wire _72703 = _66112 ^ _66116;
  wire _72704 = _72702 ^ _72703;
  wire _72705 = uncoded_block[1575] ^ uncoded_block[1607];
  wire _72706 = _66117 ^ _72705;
  wire _72707 = uncoded_block[1648] ^ uncoded_block[1687];
  wire _72708 = _72707 ^ uncoded_block[1718];
  wire _72709 = _72706 ^ _72708;
  wire _72710 = _72704 ^ _72709;
  wire _72711 = _72701 ^ _72710;
  wire _72712 = _4001 ^ _11344;
  wire _72713 = _72712 ^ _58345;
  wire _72714 = _60128 ^ _72713;
  wire _72715 = _15590 ^ _4008;
  wire _72716 = _72715 ^ _24;
  wire _72717 = _72716 ^ _60138;
  wire _72718 = _72714 ^ _72717;
  wire _72719 = _4735 ^ _13558;
  wire _72720 = _33894 ^ _903;
  wire _72721 = _72719 ^ _72720;
  wire _72722 = _60141 ^ _72721;
  wire _72723 = _60145 ^ _15608;
  wire _72724 = _46546 ^ _4034;
  wire _72725 = _72724 ^ _38310;
  wire _72726 = _72723 ^ _72725;
  wire _72727 = _72722 ^ _72726;
  wire _72728 = _72718 ^ _72727;
  wire _72729 = _9729 ^ _56659;
  wire _72730 = _69347 ^ _72729;
  wire _72731 = _69346 ^ _72730;
  wire _72732 = _68467 ^ _58373;
  wire _72733 = _4053 ^ _8589;
  wire _72734 = _72733 ^ _32646;
  wire _72735 = _72732 ^ _72734;
  wire _72736 = _72731 ^ _72735;
  wire _72737 = _20979 ^ _941;
  wire _72738 = _72737 ^ _36332;
  wire _72739 = _947 ^ _89;
  wire _72740 = _18583 ^ _6805;
  wire _72741 = _72739 ^ _72740;
  wire _72742 = _72738 ^ _72741;
  wire _72743 = _12479 ^ _6806;
  wire _72744 = _72743 ^ _14625;
  wire _72745 = _14626 ^ _29639;
  wire _72746 = _72744 ^ _72745;
  wire _72747 = _72742 ^ _72746;
  wire _72748 = _72736 ^ _72747;
  wire _72749 = _72728 ^ _72748;
  wire _72750 = _1776 ^ _44461;
  wire _72751 = _9756 ^ _6179;
  wire _72752 = _72751 ^ _60181;
  wire _72753 = _72750 ^ _72752;
  wire _72754 = _60185 ^ _21935;
  wire _72755 = _60184 ^ _72754;
  wire _72756 = _72753 ^ _72755;
  wire _72757 = _21942 ^ _3346;
  wire _72758 = _72757 ^ _23322;
  wire _72759 = _3352 ^ _1825;
  wire _72760 = _4129 ^ _6218;
  wire _72761 = _72759 ^ _72760;
  wire _72762 = _72758 ^ _72761;
  wire _72763 = _69378 ^ _72762;
  wire _72764 = _72756 ^ _72763;
  wire _72765 = _35170 ^ _168;
  wire _72766 = _72765 ^ _49225;
  wire _72767 = _69388 ^ _72766;
  wire _72768 = _55530 ^ _46607;
  wire _72769 = _29677 ^ _72768;
  wire _72770 = _10907 ^ _12006;
  wire _72771 = _72770 ^ _30137;
  wire _72772 = _72769 ^ _72771;
  wire _72773 = _72767 ^ _72772;
  wire _72774 = _60214 ^ _60218;
  wire _72775 = _4163 ^ _4874;
  wire _72776 = _197 ^ _34771;
  wire _72777 = _72775 ^ _72776;
  wire _72778 = _72774 ^ _72777;
  wire _72779 = uncoded_block[439] ^ uncoded_block[445];
  wire _72780 = _10352 ^ _72779;
  wire _72781 = _72780 ^ _3412;
  wire _72782 = _69403 ^ _4189;
  wire _72783 = _50820 ^ _72782;
  wire _72784 = _72781 ^ _72783;
  wire _72785 = _72778 ^ _72784;
  wire _72786 = _72773 ^ _72785;
  wire _72787 = _72764 ^ _72786;
  wire _72788 = _72749 ^ _72787;
  wire _72789 = _15212 ^ _13135;
  wire _72790 = _58444 ^ _72789;
  wire _72791 = _17198 ^ _1094;
  wire _72792 = _1097 ^ _1892;
  wire _72793 = _72791 ^ _72792;
  wire _72794 = _72790 ^ _72793;
  wire _72795 = _33579 ^ _68544;
  wire _72796 = _72795 ^ _68547;
  wire _72797 = _72794 ^ _72796;
  wire _72798 = _58461 ^ _52792;
  wire _72799 = _68552 ^ _72798;
  wire _72800 = _1130 ^ _18684;
  wire _72801 = _265 ^ _2696;
  wire _72802 = _72800 ^ _72801;
  wire _72803 = _19656 ^ _1938;
  wire _72804 = _17721 ^ _5646;
  wire _72805 = _72803 ^ _72804;
  wire _72806 = _72802 ^ _72805;
  wire _72807 = _72799 ^ _72806;
  wire _72808 = _72797 ^ _72807;
  wire _72809 = _8152 ^ _16734;
  wire _72810 = _13713 ^ _6960;
  wire _72811 = _72809 ^ _72810;
  wire _72812 = _2719 ^ _6966;
  wire _72813 = _12071 ^ _16740;
  wire _72814 = _72812 ^ _72813;
  wire _72815 = _72811 ^ _72814;
  wire _72816 = _36018 ^ _40796;
  wire _72817 = _64518 ^ _7582;
  wire _72818 = _72817 ^ _54723;
  wire _72819 = _72816 ^ _72818;
  wire _72820 = _72815 ^ _72819;
  wire _72821 = _1968 ^ _19191;
  wire _72822 = _31938 ^ _72821;
  wire _72823 = _18716 ^ _325;
  wire _72824 = _72823 ^ _31519;
  wire _72825 = _72822 ^ _72824;
  wire _72826 = _5685 ^ _1192;
  wire _72827 = _69448 ^ _72826;
  wire _72828 = _19201 ^ _5002;
  wire _72829 = _72828 ^ _69456;
  wire _72830 = _72827 ^ _72829;
  wire _72831 = _72825 ^ _72830;
  wire _72832 = _72820 ^ _72831;
  wire _72833 = _72808 ^ _72832;
  wire _72834 = _68584 ^ _352;
  wire _72835 = _72834 ^ _20666;
  wire _72836 = _2003 ^ _3556;
  wire _72837 = _38457 ^ _72836;
  wire _72838 = _72835 ^ _72837;
  wire _72839 = _69460 ^ _10470;
  wire _72840 = _72839 ^ _15800;
  wire _72841 = _68596 ^ _68598;
  wire _72842 = _72840 ^ _72841;
  wire _72843 = _72838 ^ _72842;
  wire _72844 = _47445 ^ _69469;
  wire _72845 = uncoded_block[801] ^ uncoded_block[805];
  wire _72846 = _72845 ^ _16791;
  wire _72847 = _53744 ^ _5045;
  wire _72848 = _72846 ^ _72847;
  wire _72849 = _72844 ^ _72848;
  wire _72850 = _69475 ^ _2813;
  wire _72851 = _57415 ^ _60301;
  wire _72852 = _72850 ^ _72851;
  wire _72853 = _72849 ^ _72852;
  wire _72854 = _72843 ^ _72853;
  wire _72855 = _19725 ^ _68610;
  wire _72856 = _72855 ^ _40472;
  wire _72857 = _14303 ^ _45348;
  wire _72858 = _72856 ^ _72857;
  wire _72859 = _61870 ^ _7660;
  wire _72860 = _11060 ^ _3616;
  wire _72861 = _72859 ^ _72860;
  wire _72862 = _49819 ^ _7665;
  wire _72863 = _25266 ^ _72862;
  wire _72864 = _72861 ^ _72863;
  wire _72865 = _72858 ^ _72864;
  wire _72866 = _42399 ^ _8260;
  wire _72867 = _72866 ^ _12170;
  wire _72868 = _453 ^ _58542;
  wire _72869 = _8842 ^ _2090;
  wire _72870 = _72868 ^ _72869;
  wire _72871 = _72867 ^ _72870;
  wire _72872 = _53214 ^ _55304;
  wire _72873 = _68635 ^ _5790;
  wire _72874 = _72873 ^ _55311;
  wire _72875 = _72872 ^ _72874;
  wire _72876 = _72871 ^ _72875;
  wire _72877 = _72865 ^ _72876;
  wire _72878 = _72854 ^ _72877;
  wire _72879 = _72833 ^ _72878;
  wire _72880 = _72788 ^ _72879;
  wire _72881 = _8859 ^ _10543;
  wire _72882 = _13277 ^ _7691;
  wire _72883 = _72881 ^ _72882;
  wire _72884 = _38929 ^ _11661;
  wire _72885 = _25295 ^ _9996;
  wire _72886 = _72884 ^ _72885;
  wire _72887 = _72883 ^ _72886;
  wire _72888 = _68647 ^ _43472;
  wire _72889 = _72888 ^ _69522;
  wire _72890 = _72887 ^ _72889;
  wire _72891 = _5163 ^ _1373;
  wire _72892 = _68657 ^ _72891;
  wire _72893 = _69526 ^ _72892;
  wire _72894 = _18822 ^ _68662;
  wire _72895 = _58577 ^ _68664;
  wire _72896 = _72894 ^ _72895;
  wire _72897 = _72893 ^ _72896;
  wire _72898 = _72890 ^ _72897;
  wire _72899 = _58584 ^ _60366;
  wire _72900 = _69536 ^ _72899;
  wire _72901 = _5188 ^ _27105;
  wire _72902 = _29877 ^ _72901;
  wire _72903 = _40539 ^ _2967;
  wire _72904 = _34961 ^ _592;
  wire _72905 = _72903 ^ _72904;
  wire _72906 = _72902 ^ _72905;
  wire _72907 = _72900 ^ _72906;
  wire _72908 = _23538 ^ _22180;
  wire _72909 = _8951 ^ _2974;
  wire _72910 = _2210 ^ _14912;
  wire _72911 = _72909 ^ _72910;
  wire _72912 = _72908 ^ _72911;
  wire _72913 = _5215 ^ _7168;
  wire _72914 = _17905 ^ _72913;
  wire _72915 = _1436 ^ _18400;
  wire _72916 = _72915 ^ _69552;
  wire _72917 = _72914 ^ _72916;
  wire _72918 = _72912 ^ _72917;
  wire _72919 = _72907 ^ _72918;
  wire _72920 = _72898 ^ _72919;
  wire _72921 = _5902 ^ _4514;
  wire _72922 = _69558 ^ _72921;
  wire _72923 = _29906 ^ _2244;
  wire _72924 = _72923 ^ _1464;
  wire _72925 = _72922 ^ _72924;
  wire _72926 = _3795 ^ _27568;
  wire _72927 = _19368 ^ _14428;
  wire _72928 = _72926 ^ _72927;
  wire _72929 = _72925 ^ _72928;
  wire _72930 = _68704 ^ _1479;
  wire _72931 = _72930 ^ _22667;
  wire _72932 = _7805 ^ _3032;
  wire _72933 = _72932 ^ _60398;
  wire _72934 = _72931 ^ _72933;
  wire _72935 = _9564 ^ _18434;
  wire _72936 = _72935 ^ _16943;
  wire _72937 = _6588 ^ _12861;
  wire _72938 = _72937 ^ _43175;
  wire _72939 = _72936 ^ _72938;
  wire _72940 = _72934 ^ _72939;
  wire _72941 = _72929 ^ _72940;
  wire _72942 = _18444 ^ _24511;
  wire _72943 = _58635 ^ _72942;
  wire _72944 = _1516 ^ _3066;
  wire _72945 = _72944 ^ _60413;
  wire _72946 = _72943 ^ _72945;
  wire _72947 = _68731 ^ _68733;
  wire _72948 = _69585 ^ _72947;
  wire _72949 = _72946 ^ _72948;
  wire _72950 = _68735 ^ _68739;
  wire _72951 = _1550 ^ _3097;
  wire _72952 = _41757 ^ _19887;
  wire _72953 = _72951 ^ _72952;
  wire _72954 = _72950 ^ _72953;
  wire _72955 = _2352 ^ _52995;
  wire _72956 = _32960 ^ _72955;
  wire _72957 = _72956 ^ _69600;
  wire _72958 = _72954 ^ _72957;
  wire _72959 = _72949 ^ _72958;
  wire _72960 = _72941 ^ _72959;
  wire _72961 = _72920 ^ _72960;
  wire _72962 = _60440 ^ _68757;
  wire _72963 = _69606 ^ _72962;
  wire _72964 = _9072 ^ _781;
  wire _72965 = _782 ^ _13479;
  wire _72966 = _72964 ^ _72965;
  wire _72967 = _40243 ^ _25454;
  wire _72968 = _17013 ^ _1621;
  wire _72969 = _72967 ^ _72968;
  wire _72970 = _72966 ^ _72969;
  wire _72971 = _72963 ^ _72970;
  wire _72972 = _68768 ^ _27649;
  wire _72973 = _33421 ^ _72972;
  wire _72974 = _2404 ^ _42177;
  wire _72975 = _6689 ^ _34255;
  wire _72976 = _72974 ^ _72975;
  wire _72977 = _72973 ^ _72976;
  wire _72978 = _72977 ^ _68779;
  wire _72979 = _72971 ^ _72978;
  wire _72980 = _844 ^ _22773;
  wire _72981 = _68786 ^ _72980;
  wire _72982 = _68784 ^ _72981;
  wire _72983 = _72982 ^ _68792;
  wire _72984 = _72979 ^ _72983;
  wire _72985 = _72961 ^ _72984;
  wire _72986 = _72880 ^ _72985;
  assign coded_block = {_865, _1682, _2452, _3208, _3992, _4709, _5421, _6079, _6723, _7346, _7952, _8543, _9133, _9687, _10222, _10786, _11339, _11886, _12414, _12982, _13533, _14037, _14558, _15072, _15581, _16071, _16559, _17055, _17557, _18055, _18538, _18998, _19492, _19958, _20446, _20931, _21406, _21860, _22324, _22784, _23245, _23685, _24146, _24601, _25048, _25494, _25935, _26378, _26844, _27240, _27679, _27994, _28432, _28745, _29175, _29585, _30033, _30477, _30914, _31354, _31775, _32200, _32607, _33030, _33452, _33876, _34276, _34672, _35093, _35484, _35864, _36286, _36706, _37109, _37515, _37907, _38288, _38693, _39096, _39486, _39878, _40280, _40661, _41025, _41431, _41818, _42202, _42578, _42849, _43256, _43629, _44011, _44414, _44788, _45146, _45539, _45926, _46147, _46523, _46912, _47282, _47659, _48041, _48410, _48789, _49147, _49501, _49624, _49998, _50379, _50717, _51107, _51480, _51799, _52102, _52350, _52676, _53048, _53367, _53570, _53951, _54223, _54577, _54961, _55138, _55447, _55820, _56172, _56403, _56635, _56961, _57253, _57588, _57800, _58045, _58341, _58711, _58983, _59248, _59401, _59664, _59919, _60125, _60477, _60614, _60737, _60930, _61066, _61251, _61396, _61567, _61760, _61986, _62127, _62350, _62453, _62610, _62816, _63024, _63162, _63402, _63552, _63761, _63996, _64154, _64332, _64456, _64627, _64776, _64859, _65050, _65290, _65345, _65418, _65475, _65546, _65603, _65660, _65741, _65874, _65928, _65999, _66076, _66128, _66220, _66277, _66328, _66419, _66474, _66532, _66586, _66641, _66695, _66749, _66845, _66902, _66977, _67060, _67168, _67239, _67341, _67393, _67465, _67562, _67618, _67670, _67723, _67780, _67857, _67911, _67967, _68050, _68106, _68185, _68244, _68296, _68353, _68435, _68796, _68875, _68974, _69031, _69084, _69160, _69214, _69260, _69328, _69640, _69713, _69765, _69819, _69893, _69962, _70035, _70112, _70183, _70236, _70288, _70316, _70345, _70370, _70398, _70426, _70453, _70480, _70506, _70535, _70565, _70594, _70624, _70653, _70683, _70713, _70742, _70769, _70796, _70825, _70855, _70880, _70906, _70936, _70962, _70991, _71017, _71046, _71074, _71101, _71130, _71160, _71189, _71219, _71248, _71276, _71305, _71332, _71360, _71388, _71418, _71445, _71471, _71499, _71528, _71555, _71583, _71609, _71639, _71669, _71697, _71725, _71755, _71783, _71810, _71833, _71863, _71892, _71920, _71950, _71975, _72005, _72030, _72060, _72088, _72118, _72146, _72173, _72200, _72229, _72258, _72286, _72316, _72345, _72375, _72405, _72433, _72460, _72489, _72517, _72545, _72573, _72602, _72632, _72660, _72690, _72711, _72986, uncoded_block[1722], uncoded_block[1721], uncoded_block[1720], uncoded_block[1719], uncoded_block[1718], uncoded_block[1717], uncoded_block[1716], uncoded_block[1715], uncoded_block[1714], uncoded_block[1713], uncoded_block[1712], uncoded_block[1711], uncoded_block[1710], uncoded_block[1709], uncoded_block[1708], uncoded_block[1707], uncoded_block[1706], uncoded_block[1705], uncoded_block[1704], uncoded_block[1703], uncoded_block[1702], uncoded_block[1701], uncoded_block[1700], uncoded_block[1699], uncoded_block[1698], uncoded_block[1697], uncoded_block[1696], uncoded_block[1695], uncoded_block[1694], uncoded_block[1693], uncoded_block[1692], uncoded_block[1691], uncoded_block[1690], uncoded_block[1689], uncoded_block[1688], uncoded_block[1687], uncoded_block[1686], uncoded_block[1685], uncoded_block[1684], uncoded_block[1683], uncoded_block[1682], uncoded_block[1681], uncoded_block[1680], uncoded_block[1679], uncoded_block[1678], uncoded_block[1677], uncoded_block[1676], uncoded_block[1675], uncoded_block[1674], uncoded_block[1673], uncoded_block[1672], uncoded_block[1671], uncoded_block[1670], uncoded_block[1669], uncoded_block[1668], uncoded_block[1667], uncoded_block[1666], uncoded_block[1665], uncoded_block[1664], uncoded_block[1663], uncoded_block[1662], uncoded_block[1661], uncoded_block[1660], uncoded_block[1659], uncoded_block[1658], uncoded_block[1657], uncoded_block[1656], uncoded_block[1655], uncoded_block[1654], uncoded_block[1653], uncoded_block[1652], uncoded_block[1651], uncoded_block[1650], uncoded_block[1649], uncoded_block[1648], uncoded_block[1647], uncoded_block[1646], uncoded_block[1645], uncoded_block[1644], uncoded_block[1643], uncoded_block[1642], uncoded_block[1641], uncoded_block[1640], uncoded_block[1639], uncoded_block[1638], uncoded_block[1637], uncoded_block[1636], uncoded_block[1635], uncoded_block[1634], uncoded_block[1633], uncoded_block[1632], uncoded_block[1631], uncoded_block[1630], uncoded_block[1629], uncoded_block[1628], uncoded_block[1627], uncoded_block[1626], uncoded_block[1625], uncoded_block[1624], uncoded_block[1623], uncoded_block[1622], uncoded_block[1621], uncoded_block[1620], uncoded_block[1619], uncoded_block[1618], uncoded_block[1617], uncoded_block[1616], uncoded_block[1615], uncoded_block[1614], uncoded_block[1613], uncoded_block[1612], uncoded_block[1611], uncoded_block[1610], uncoded_block[1609], uncoded_block[1608], uncoded_block[1607], uncoded_block[1606], uncoded_block[1605], uncoded_block[1604], uncoded_block[1603], uncoded_block[1602], uncoded_block[1601], uncoded_block[1600], uncoded_block[1599], uncoded_block[1598], uncoded_block[1597], uncoded_block[1596], uncoded_block[1595], uncoded_block[1594], uncoded_block[1593], uncoded_block[1592], uncoded_block[1591], uncoded_block[1590], uncoded_block[1589], uncoded_block[1588], uncoded_block[1587], uncoded_block[1586], uncoded_block[1585], uncoded_block[1584], uncoded_block[1583], uncoded_block[1582], uncoded_block[1581], uncoded_block[1580], uncoded_block[1579], uncoded_block[1578], uncoded_block[1577], uncoded_block[1576], uncoded_block[1575], uncoded_block[1574], uncoded_block[1573], uncoded_block[1572], uncoded_block[1571], uncoded_block[1570], uncoded_block[1569], uncoded_block[1568], uncoded_block[1567], uncoded_block[1566], uncoded_block[1565], uncoded_block[1564], uncoded_block[1563], uncoded_block[1562], uncoded_block[1561], uncoded_block[1560], uncoded_block[1559], uncoded_block[1558], uncoded_block[1557], uncoded_block[1556], uncoded_block[1555], uncoded_block[1554], uncoded_block[1553], uncoded_block[1552], uncoded_block[1551], uncoded_block[1550], uncoded_block[1549], uncoded_block[1548], uncoded_block[1547], uncoded_block[1546], uncoded_block[1545], uncoded_block[1544], uncoded_block[1543], uncoded_block[1542], uncoded_block[1541], uncoded_block[1540], uncoded_block[1539], uncoded_block[1538], uncoded_block[1537], uncoded_block[1536], uncoded_block[1535], uncoded_block[1534], uncoded_block[1533], uncoded_block[1532], uncoded_block[1531], uncoded_block[1530], uncoded_block[1529], uncoded_block[1528], uncoded_block[1527], uncoded_block[1526], uncoded_block[1525], uncoded_block[1524], uncoded_block[1523], uncoded_block[1522], uncoded_block[1521], uncoded_block[1520], uncoded_block[1519], uncoded_block[1518], uncoded_block[1517], uncoded_block[1516], uncoded_block[1515], uncoded_block[1514], uncoded_block[1513], uncoded_block[1512], uncoded_block[1511], uncoded_block[1510], uncoded_block[1509], uncoded_block[1508], uncoded_block[1507], uncoded_block[1506], uncoded_block[1505], uncoded_block[1504], uncoded_block[1503], uncoded_block[1502], uncoded_block[1501], uncoded_block[1500], uncoded_block[1499], uncoded_block[1498], uncoded_block[1497], uncoded_block[1496], uncoded_block[1495], uncoded_block[1494], uncoded_block[1493], uncoded_block[1492], uncoded_block[1491], uncoded_block[1490], uncoded_block[1489], uncoded_block[1488], uncoded_block[1487], uncoded_block[1486], uncoded_block[1485], uncoded_block[1484], uncoded_block[1483], uncoded_block[1482], uncoded_block[1481], uncoded_block[1480], uncoded_block[1479], uncoded_block[1478], uncoded_block[1477], uncoded_block[1476], uncoded_block[1475], uncoded_block[1474], uncoded_block[1473], uncoded_block[1472], uncoded_block[1471], uncoded_block[1470], uncoded_block[1469], uncoded_block[1468], uncoded_block[1467], uncoded_block[1466], uncoded_block[1465], uncoded_block[1464], uncoded_block[1463], uncoded_block[1462], uncoded_block[1461], uncoded_block[1460], uncoded_block[1459], uncoded_block[1458], uncoded_block[1457], uncoded_block[1456], uncoded_block[1455], uncoded_block[1454], uncoded_block[1453], uncoded_block[1452], uncoded_block[1451], uncoded_block[1450], uncoded_block[1449], uncoded_block[1448], uncoded_block[1447], uncoded_block[1446], uncoded_block[1445], uncoded_block[1444], uncoded_block[1443], uncoded_block[1442], uncoded_block[1441], uncoded_block[1440], uncoded_block[1439], uncoded_block[1438], uncoded_block[1437], uncoded_block[1436], uncoded_block[1435], uncoded_block[1434], uncoded_block[1433], uncoded_block[1432], uncoded_block[1431], uncoded_block[1430], uncoded_block[1429], uncoded_block[1428], uncoded_block[1427], uncoded_block[1426], uncoded_block[1425], uncoded_block[1424], uncoded_block[1423], uncoded_block[1422], uncoded_block[1421], uncoded_block[1420], uncoded_block[1419], uncoded_block[1418], uncoded_block[1417], uncoded_block[1416], uncoded_block[1415], uncoded_block[1414], uncoded_block[1413], uncoded_block[1412], uncoded_block[1411], uncoded_block[1410], uncoded_block[1409], uncoded_block[1408], uncoded_block[1407], uncoded_block[1406], uncoded_block[1405], uncoded_block[1404], uncoded_block[1403], uncoded_block[1402], uncoded_block[1401], uncoded_block[1400], uncoded_block[1399], uncoded_block[1398], uncoded_block[1397], uncoded_block[1396], uncoded_block[1395], uncoded_block[1394], uncoded_block[1393], uncoded_block[1392], uncoded_block[1391], uncoded_block[1390], uncoded_block[1389], uncoded_block[1388], uncoded_block[1387], uncoded_block[1386], uncoded_block[1385], uncoded_block[1384], uncoded_block[1383], uncoded_block[1382], uncoded_block[1381], uncoded_block[1380], uncoded_block[1379], uncoded_block[1378], uncoded_block[1377], uncoded_block[1376], uncoded_block[1375], uncoded_block[1374], uncoded_block[1373], uncoded_block[1372], uncoded_block[1371], uncoded_block[1370], uncoded_block[1369], uncoded_block[1368], uncoded_block[1367], uncoded_block[1366], uncoded_block[1365], uncoded_block[1364], uncoded_block[1363], uncoded_block[1362], uncoded_block[1361], uncoded_block[1360], uncoded_block[1359], uncoded_block[1358], uncoded_block[1357], uncoded_block[1356], uncoded_block[1355], uncoded_block[1354], uncoded_block[1353], uncoded_block[1352], uncoded_block[1351], uncoded_block[1350], uncoded_block[1349], uncoded_block[1348], uncoded_block[1347], uncoded_block[1346], uncoded_block[1345], uncoded_block[1344], uncoded_block[1343], uncoded_block[1342], uncoded_block[1341], uncoded_block[1340], uncoded_block[1339], uncoded_block[1338], uncoded_block[1337], uncoded_block[1336], uncoded_block[1335], uncoded_block[1334], uncoded_block[1333], uncoded_block[1332], uncoded_block[1331], uncoded_block[1330], uncoded_block[1329], uncoded_block[1328], uncoded_block[1327], uncoded_block[1326], uncoded_block[1325], uncoded_block[1324], uncoded_block[1323], uncoded_block[1322], uncoded_block[1321], uncoded_block[1320], uncoded_block[1319], uncoded_block[1318], uncoded_block[1317], uncoded_block[1316], uncoded_block[1315], uncoded_block[1314], uncoded_block[1313], uncoded_block[1312], uncoded_block[1311], uncoded_block[1310], uncoded_block[1309], uncoded_block[1308], uncoded_block[1307], uncoded_block[1306], uncoded_block[1305], uncoded_block[1304], uncoded_block[1303], uncoded_block[1302], uncoded_block[1301], uncoded_block[1300], uncoded_block[1299], uncoded_block[1298], uncoded_block[1297], uncoded_block[1296], uncoded_block[1295], uncoded_block[1294], uncoded_block[1293], uncoded_block[1292], uncoded_block[1291], uncoded_block[1290], uncoded_block[1289], uncoded_block[1288], uncoded_block[1287], uncoded_block[1286], uncoded_block[1285], uncoded_block[1284], uncoded_block[1283], uncoded_block[1282], uncoded_block[1281], uncoded_block[1280], uncoded_block[1279], uncoded_block[1278], uncoded_block[1277], uncoded_block[1276], uncoded_block[1275], uncoded_block[1274], uncoded_block[1273], uncoded_block[1272], uncoded_block[1271], uncoded_block[1270], uncoded_block[1269], uncoded_block[1268], uncoded_block[1267], uncoded_block[1266], uncoded_block[1265], uncoded_block[1264], uncoded_block[1263], uncoded_block[1262], uncoded_block[1261], uncoded_block[1260], uncoded_block[1259], uncoded_block[1258], uncoded_block[1257], uncoded_block[1256], uncoded_block[1255], uncoded_block[1254], uncoded_block[1253], uncoded_block[1252], uncoded_block[1251], uncoded_block[1250], uncoded_block[1249], uncoded_block[1248], uncoded_block[1247], uncoded_block[1246], uncoded_block[1245], uncoded_block[1244], uncoded_block[1243], uncoded_block[1242], uncoded_block[1241], uncoded_block[1240], uncoded_block[1239], uncoded_block[1238], uncoded_block[1237], uncoded_block[1236], uncoded_block[1235], uncoded_block[1234], uncoded_block[1233], uncoded_block[1232], uncoded_block[1231], uncoded_block[1230], uncoded_block[1229], uncoded_block[1228], uncoded_block[1227], uncoded_block[1226], uncoded_block[1225], uncoded_block[1224], uncoded_block[1223], uncoded_block[1222], uncoded_block[1221], uncoded_block[1220], uncoded_block[1219], uncoded_block[1218], uncoded_block[1217], uncoded_block[1216], uncoded_block[1215], uncoded_block[1214], uncoded_block[1213], uncoded_block[1212], uncoded_block[1211], uncoded_block[1210], uncoded_block[1209], uncoded_block[1208], uncoded_block[1207], uncoded_block[1206], uncoded_block[1205], uncoded_block[1204], uncoded_block[1203], uncoded_block[1202], uncoded_block[1201], uncoded_block[1200], uncoded_block[1199], uncoded_block[1198], uncoded_block[1197], uncoded_block[1196], uncoded_block[1195], uncoded_block[1194], uncoded_block[1193], uncoded_block[1192], uncoded_block[1191], uncoded_block[1190], uncoded_block[1189], uncoded_block[1188], uncoded_block[1187], uncoded_block[1186], uncoded_block[1185], uncoded_block[1184], uncoded_block[1183], uncoded_block[1182], uncoded_block[1181], uncoded_block[1180], uncoded_block[1179], uncoded_block[1178], uncoded_block[1177], uncoded_block[1176], uncoded_block[1175], uncoded_block[1174], uncoded_block[1173], uncoded_block[1172], uncoded_block[1171], uncoded_block[1170], uncoded_block[1169], uncoded_block[1168], uncoded_block[1167], uncoded_block[1166], uncoded_block[1165], uncoded_block[1164], uncoded_block[1163], uncoded_block[1162], uncoded_block[1161], uncoded_block[1160], uncoded_block[1159], uncoded_block[1158], uncoded_block[1157], uncoded_block[1156], uncoded_block[1155], uncoded_block[1154], uncoded_block[1153], uncoded_block[1152], uncoded_block[1151], uncoded_block[1150], uncoded_block[1149], uncoded_block[1148], uncoded_block[1147], uncoded_block[1146], uncoded_block[1145], uncoded_block[1144], uncoded_block[1143], uncoded_block[1142], uncoded_block[1141], uncoded_block[1140], uncoded_block[1139], uncoded_block[1138], uncoded_block[1137], uncoded_block[1136], uncoded_block[1135], uncoded_block[1134], uncoded_block[1133], uncoded_block[1132], uncoded_block[1131], uncoded_block[1130], uncoded_block[1129], uncoded_block[1128], uncoded_block[1127], uncoded_block[1126], uncoded_block[1125], uncoded_block[1124], uncoded_block[1123], uncoded_block[1122], uncoded_block[1121], uncoded_block[1120], uncoded_block[1119], uncoded_block[1118], uncoded_block[1117], uncoded_block[1116], uncoded_block[1115], uncoded_block[1114], uncoded_block[1113], uncoded_block[1112], uncoded_block[1111], uncoded_block[1110], uncoded_block[1109], uncoded_block[1108], uncoded_block[1107], uncoded_block[1106], uncoded_block[1105], uncoded_block[1104], uncoded_block[1103], uncoded_block[1102], uncoded_block[1101], uncoded_block[1100], uncoded_block[1099], uncoded_block[1098], uncoded_block[1097], uncoded_block[1096], uncoded_block[1095], uncoded_block[1094], uncoded_block[1093], uncoded_block[1092], uncoded_block[1091], uncoded_block[1090], uncoded_block[1089], uncoded_block[1088], uncoded_block[1087], uncoded_block[1086], uncoded_block[1085], uncoded_block[1084], uncoded_block[1083], uncoded_block[1082], uncoded_block[1081], uncoded_block[1080], uncoded_block[1079], uncoded_block[1078], uncoded_block[1077], uncoded_block[1076], uncoded_block[1075], uncoded_block[1074], uncoded_block[1073], uncoded_block[1072], uncoded_block[1071], uncoded_block[1070], uncoded_block[1069], uncoded_block[1068], uncoded_block[1067], uncoded_block[1066], uncoded_block[1065], uncoded_block[1064], uncoded_block[1063], uncoded_block[1062], uncoded_block[1061], uncoded_block[1060], uncoded_block[1059], uncoded_block[1058], uncoded_block[1057], uncoded_block[1056], uncoded_block[1055], uncoded_block[1054], uncoded_block[1053], uncoded_block[1052], uncoded_block[1051], uncoded_block[1050], uncoded_block[1049], uncoded_block[1048], uncoded_block[1047], uncoded_block[1046], uncoded_block[1045], uncoded_block[1044], uncoded_block[1043], uncoded_block[1042], uncoded_block[1041], uncoded_block[1040], uncoded_block[1039], uncoded_block[1038], uncoded_block[1037], uncoded_block[1036], uncoded_block[1035], uncoded_block[1034], uncoded_block[1033], uncoded_block[1032], uncoded_block[1031], uncoded_block[1030], uncoded_block[1029], uncoded_block[1028], uncoded_block[1027], uncoded_block[1026], uncoded_block[1025], uncoded_block[1024], uncoded_block[1023], uncoded_block[1022], uncoded_block[1021], uncoded_block[1020], uncoded_block[1019], uncoded_block[1018], uncoded_block[1017], uncoded_block[1016], uncoded_block[1015], uncoded_block[1014], uncoded_block[1013], uncoded_block[1012], uncoded_block[1011], uncoded_block[1010], uncoded_block[1009], uncoded_block[1008], uncoded_block[1007], uncoded_block[1006], uncoded_block[1005], uncoded_block[1004], uncoded_block[1003], uncoded_block[1002], uncoded_block[1001], uncoded_block[1000], uncoded_block[999], uncoded_block[998], uncoded_block[997], uncoded_block[996], uncoded_block[995], uncoded_block[994], uncoded_block[993], uncoded_block[992], uncoded_block[991], uncoded_block[990], uncoded_block[989], uncoded_block[988], uncoded_block[987], uncoded_block[986], uncoded_block[985], uncoded_block[984], uncoded_block[983], uncoded_block[982], uncoded_block[981], uncoded_block[980], uncoded_block[979], uncoded_block[978], uncoded_block[977], uncoded_block[976], uncoded_block[975], uncoded_block[974], uncoded_block[973], uncoded_block[972], uncoded_block[971], uncoded_block[970], uncoded_block[969], uncoded_block[968], uncoded_block[967], uncoded_block[966], uncoded_block[965], uncoded_block[964], uncoded_block[963], uncoded_block[962], uncoded_block[961], uncoded_block[960], uncoded_block[959], uncoded_block[958], uncoded_block[957], uncoded_block[956], uncoded_block[955], uncoded_block[954], uncoded_block[953], uncoded_block[952], uncoded_block[951], uncoded_block[950], uncoded_block[949], uncoded_block[948], uncoded_block[947], uncoded_block[946], uncoded_block[945], uncoded_block[944], uncoded_block[943], uncoded_block[942], uncoded_block[941], uncoded_block[940], uncoded_block[939], uncoded_block[938], uncoded_block[937], uncoded_block[936], uncoded_block[935], uncoded_block[934], uncoded_block[933], uncoded_block[932], uncoded_block[931], uncoded_block[930], uncoded_block[929], uncoded_block[928], uncoded_block[927], uncoded_block[926], uncoded_block[925], uncoded_block[924], uncoded_block[923], uncoded_block[922], uncoded_block[921], uncoded_block[920], uncoded_block[919], uncoded_block[918], uncoded_block[917], uncoded_block[916], uncoded_block[915], uncoded_block[914], uncoded_block[913], uncoded_block[912], uncoded_block[911], uncoded_block[910], uncoded_block[909], uncoded_block[908], uncoded_block[907], uncoded_block[906], uncoded_block[905], uncoded_block[904], uncoded_block[903], uncoded_block[902], uncoded_block[901], uncoded_block[900], uncoded_block[899], uncoded_block[898], uncoded_block[897], uncoded_block[896], uncoded_block[895], uncoded_block[894], uncoded_block[893], uncoded_block[892], uncoded_block[891], uncoded_block[890], uncoded_block[889], uncoded_block[888], uncoded_block[887], uncoded_block[886], uncoded_block[885], uncoded_block[884], uncoded_block[883], uncoded_block[882], uncoded_block[881], uncoded_block[880], uncoded_block[879], uncoded_block[878], uncoded_block[877], uncoded_block[876], uncoded_block[875], uncoded_block[874], uncoded_block[873], uncoded_block[872], uncoded_block[871], uncoded_block[870], uncoded_block[869], uncoded_block[868], uncoded_block[867], uncoded_block[866], uncoded_block[865], uncoded_block[864], uncoded_block[863], uncoded_block[862], uncoded_block[861], uncoded_block[860], uncoded_block[859], uncoded_block[858], uncoded_block[857], uncoded_block[856], uncoded_block[855], uncoded_block[854], uncoded_block[853], uncoded_block[852], uncoded_block[851], uncoded_block[850], uncoded_block[849], uncoded_block[848], uncoded_block[847], uncoded_block[846], uncoded_block[845], uncoded_block[844], uncoded_block[843], uncoded_block[842], uncoded_block[841], uncoded_block[840], uncoded_block[839], uncoded_block[838], uncoded_block[837], uncoded_block[836], uncoded_block[835], uncoded_block[834], uncoded_block[833], uncoded_block[832], uncoded_block[831], uncoded_block[830], uncoded_block[829], uncoded_block[828], uncoded_block[827], uncoded_block[826], uncoded_block[825], uncoded_block[824], uncoded_block[823], uncoded_block[822], uncoded_block[821], uncoded_block[820], uncoded_block[819], uncoded_block[818], uncoded_block[817], uncoded_block[816], uncoded_block[815], uncoded_block[814], uncoded_block[813], uncoded_block[812], uncoded_block[811], uncoded_block[810], uncoded_block[809], uncoded_block[808], uncoded_block[807], uncoded_block[806], uncoded_block[805], uncoded_block[804], uncoded_block[803], uncoded_block[802], uncoded_block[801], uncoded_block[800], uncoded_block[799], uncoded_block[798], uncoded_block[797], uncoded_block[796], uncoded_block[795], uncoded_block[794], uncoded_block[793], uncoded_block[792], uncoded_block[791], uncoded_block[790], uncoded_block[789], uncoded_block[788], uncoded_block[787], uncoded_block[786], uncoded_block[785], uncoded_block[784], uncoded_block[783], uncoded_block[782], uncoded_block[781], uncoded_block[780], uncoded_block[779], uncoded_block[778], uncoded_block[777], uncoded_block[776], uncoded_block[775], uncoded_block[774], uncoded_block[773], uncoded_block[772], uncoded_block[771], uncoded_block[770], uncoded_block[769], uncoded_block[768], uncoded_block[767], uncoded_block[766], uncoded_block[765], uncoded_block[764], uncoded_block[763], uncoded_block[762], uncoded_block[761], uncoded_block[760], uncoded_block[759], uncoded_block[758], uncoded_block[757], uncoded_block[756], uncoded_block[755], uncoded_block[754], uncoded_block[753], uncoded_block[752], uncoded_block[751], uncoded_block[750], uncoded_block[749], uncoded_block[748], uncoded_block[747], uncoded_block[746], uncoded_block[745], uncoded_block[744], uncoded_block[743], uncoded_block[742], uncoded_block[741], uncoded_block[740], uncoded_block[739], uncoded_block[738], uncoded_block[737], uncoded_block[736], uncoded_block[735], uncoded_block[734], uncoded_block[733], uncoded_block[732], uncoded_block[731], uncoded_block[730], uncoded_block[729], uncoded_block[728], uncoded_block[727], uncoded_block[726], uncoded_block[725], uncoded_block[724], uncoded_block[723], uncoded_block[722], uncoded_block[721], uncoded_block[720], uncoded_block[719], uncoded_block[718], uncoded_block[717], uncoded_block[716], uncoded_block[715], uncoded_block[714], uncoded_block[713], uncoded_block[712], uncoded_block[711], uncoded_block[710], uncoded_block[709], uncoded_block[708], uncoded_block[707], uncoded_block[706], uncoded_block[705], uncoded_block[704], uncoded_block[703], uncoded_block[702], uncoded_block[701], uncoded_block[700], uncoded_block[699], uncoded_block[698], uncoded_block[697], uncoded_block[696], uncoded_block[695], uncoded_block[694], uncoded_block[693], uncoded_block[692], uncoded_block[691], uncoded_block[690], uncoded_block[689], uncoded_block[688], uncoded_block[687], uncoded_block[686], uncoded_block[685], uncoded_block[684], uncoded_block[683], uncoded_block[682], uncoded_block[681], uncoded_block[680], uncoded_block[679], uncoded_block[678], uncoded_block[677], uncoded_block[676], uncoded_block[675], uncoded_block[674], uncoded_block[673], uncoded_block[672], uncoded_block[671], uncoded_block[670], uncoded_block[669], uncoded_block[668], uncoded_block[667], uncoded_block[666], uncoded_block[665], uncoded_block[664], uncoded_block[663], uncoded_block[662], uncoded_block[661], uncoded_block[660], uncoded_block[659], uncoded_block[658], uncoded_block[657], uncoded_block[656], uncoded_block[655], uncoded_block[654], uncoded_block[653], uncoded_block[652], uncoded_block[651], uncoded_block[650], uncoded_block[649], uncoded_block[648], uncoded_block[647], uncoded_block[646], uncoded_block[645], uncoded_block[644], uncoded_block[643], uncoded_block[642], uncoded_block[641], uncoded_block[640], uncoded_block[639], uncoded_block[638], uncoded_block[637], uncoded_block[636], uncoded_block[635], uncoded_block[634], uncoded_block[633], uncoded_block[632], uncoded_block[631], uncoded_block[630], uncoded_block[629], uncoded_block[628], uncoded_block[627], uncoded_block[626], uncoded_block[625], uncoded_block[624], uncoded_block[623], uncoded_block[622], uncoded_block[621], uncoded_block[620], uncoded_block[619], uncoded_block[618], uncoded_block[617], uncoded_block[616], uncoded_block[615], uncoded_block[614], uncoded_block[613], uncoded_block[612], uncoded_block[611], uncoded_block[610], uncoded_block[609], uncoded_block[608], uncoded_block[607], uncoded_block[606], uncoded_block[605], uncoded_block[604], uncoded_block[603], uncoded_block[602], uncoded_block[601], uncoded_block[600], uncoded_block[599], uncoded_block[598], uncoded_block[597], uncoded_block[596], uncoded_block[595], uncoded_block[594], uncoded_block[593], uncoded_block[592], uncoded_block[591], uncoded_block[590], uncoded_block[589], uncoded_block[588], uncoded_block[587], uncoded_block[586], uncoded_block[585], uncoded_block[584], uncoded_block[583], uncoded_block[582], uncoded_block[581], uncoded_block[580], uncoded_block[579], uncoded_block[578], uncoded_block[577], uncoded_block[576], uncoded_block[575], uncoded_block[574], uncoded_block[573], uncoded_block[572], uncoded_block[571], uncoded_block[570], uncoded_block[569], uncoded_block[568], uncoded_block[567], uncoded_block[566], uncoded_block[565], uncoded_block[564], uncoded_block[563], uncoded_block[562], uncoded_block[561], uncoded_block[560], uncoded_block[559], uncoded_block[558], uncoded_block[557], uncoded_block[556], uncoded_block[555], uncoded_block[554], uncoded_block[553], uncoded_block[552], uncoded_block[551], uncoded_block[550], uncoded_block[549], uncoded_block[548], uncoded_block[547], uncoded_block[546], uncoded_block[545], uncoded_block[544], uncoded_block[543], uncoded_block[542], uncoded_block[541], uncoded_block[540], uncoded_block[539], uncoded_block[538], uncoded_block[537], uncoded_block[536], uncoded_block[535], uncoded_block[534], uncoded_block[533], uncoded_block[532], uncoded_block[531], uncoded_block[530], uncoded_block[529], uncoded_block[528], uncoded_block[527], uncoded_block[526], uncoded_block[525], uncoded_block[524], uncoded_block[523], uncoded_block[522], uncoded_block[521], uncoded_block[520], uncoded_block[519], uncoded_block[518], uncoded_block[517], uncoded_block[516], uncoded_block[515], uncoded_block[514], uncoded_block[513], uncoded_block[512], uncoded_block[511], uncoded_block[510], uncoded_block[509], uncoded_block[508], uncoded_block[507], uncoded_block[506], uncoded_block[505], uncoded_block[504], uncoded_block[503], uncoded_block[502], uncoded_block[501], uncoded_block[500], uncoded_block[499], uncoded_block[498], uncoded_block[497], uncoded_block[496], uncoded_block[495], uncoded_block[494], uncoded_block[493], uncoded_block[492], uncoded_block[491], uncoded_block[490], uncoded_block[489], uncoded_block[488], uncoded_block[487], uncoded_block[486], uncoded_block[485], uncoded_block[484], uncoded_block[483], uncoded_block[482], uncoded_block[481], uncoded_block[480], uncoded_block[479], uncoded_block[478], uncoded_block[477], uncoded_block[476], uncoded_block[475], uncoded_block[474], uncoded_block[473], uncoded_block[472], uncoded_block[471], uncoded_block[470], uncoded_block[469], uncoded_block[468], uncoded_block[467], uncoded_block[466], uncoded_block[465], uncoded_block[464], uncoded_block[463], uncoded_block[462], uncoded_block[461], uncoded_block[460], uncoded_block[459], uncoded_block[458], uncoded_block[457], uncoded_block[456], uncoded_block[455], uncoded_block[454], uncoded_block[453], uncoded_block[452], uncoded_block[451], uncoded_block[450], uncoded_block[449], uncoded_block[448], uncoded_block[447], uncoded_block[446], uncoded_block[445], uncoded_block[444], uncoded_block[443], uncoded_block[442], uncoded_block[441], uncoded_block[440], uncoded_block[439], uncoded_block[438], uncoded_block[437], uncoded_block[436], uncoded_block[435], uncoded_block[434], uncoded_block[433], uncoded_block[432], uncoded_block[431], uncoded_block[430], uncoded_block[429], uncoded_block[428], uncoded_block[427], uncoded_block[426], uncoded_block[425], uncoded_block[424], uncoded_block[423], uncoded_block[422], uncoded_block[421], uncoded_block[420], uncoded_block[419], uncoded_block[418], uncoded_block[417], uncoded_block[416], uncoded_block[415], uncoded_block[414], uncoded_block[413], uncoded_block[412], uncoded_block[411], uncoded_block[410], uncoded_block[409], uncoded_block[408], uncoded_block[407], uncoded_block[406], uncoded_block[405], uncoded_block[404], uncoded_block[403], uncoded_block[402], uncoded_block[401], uncoded_block[400], uncoded_block[399], uncoded_block[398], uncoded_block[397], uncoded_block[396], uncoded_block[395], uncoded_block[394], uncoded_block[393], uncoded_block[392], uncoded_block[391], uncoded_block[390], uncoded_block[389], uncoded_block[388], uncoded_block[387], uncoded_block[386], uncoded_block[385], uncoded_block[384], uncoded_block[383], uncoded_block[382], uncoded_block[381], uncoded_block[380], uncoded_block[379], uncoded_block[378], uncoded_block[377], uncoded_block[376], uncoded_block[375], uncoded_block[374], uncoded_block[373], uncoded_block[372], uncoded_block[371], uncoded_block[370], uncoded_block[369], uncoded_block[368], uncoded_block[367], uncoded_block[366], uncoded_block[365], uncoded_block[364], uncoded_block[363], uncoded_block[362], uncoded_block[361], uncoded_block[360], uncoded_block[359], uncoded_block[358], uncoded_block[357], uncoded_block[356], uncoded_block[355], uncoded_block[354], uncoded_block[353], uncoded_block[352], uncoded_block[351], uncoded_block[350], uncoded_block[349], uncoded_block[348], uncoded_block[347], uncoded_block[346], uncoded_block[345], uncoded_block[344], uncoded_block[343], uncoded_block[342], uncoded_block[341], uncoded_block[340], uncoded_block[339], uncoded_block[338], uncoded_block[337], uncoded_block[336], uncoded_block[335], uncoded_block[334], uncoded_block[333], uncoded_block[332], uncoded_block[331], uncoded_block[330], uncoded_block[329], uncoded_block[328], uncoded_block[327], uncoded_block[326], uncoded_block[325], uncoded_block[324], uncoded_block[323], uncoded_block[322], uncoded_block[321], uncoded_block[320], uncoded_block[319], uncoded_block[318], uncoded_block[317], uncoded_block[316], uncoded_block[315], uncoded_block[314], uncoded_block[313], uncoded_block[312], uncoded_block[311], uncoded_block[310], uncoded_block[309], uncoded_block[308], uncoded_block[307], uncoded_block[306], uncoded_block[305], uncoded_block[304], uncoded_block[303], uncoded_block[302], uncoded_block[301], uncoded_block[300], uncoded_block[299], uncoded_block[298], uncoded_block[297], uncoded_block[296], uncoded_block[295], uncoded_block[294], uncoded_block[293], uncoded_block[292], uncoded_block[291], uncoded_block[290], uncoded_block[289], uncoded_block[288], uncoded_block[287], uncoded_block[286], uncoded_block[285], uncoded_block[284], uncoded_block[283], uncoded_block[282], uncoded_block[281], uncoded_block[280], uncoded_block[279], uncoded_block[278], uncoded_block[277], uncoded_block[276], uncoded_block[275], uncoded_block[274], uncoded_block[273], uncoded_block[272], uncoded_block[271], uncoded_block[270], uncoded_block[269], uncoded_block[268], uncoded_block[267], uncoded_block[266], uncoded_block[265], uncoded_block[264], uncoded_block[263], uncoded_block[262], uncoded_block[261], uncoded_block[260], uncoded_block[259], uncoded_block[258], uncoded_block[257], uncoded_block[256], uncoded_block[255], uncoded_block[254], uncoded_block[253], uncoded_block[252], uncoded_block[251], uncoded_block[250], uncoded_block[249], uncoded_block[248], uncoded_block[247], uncoded_block[246], uncoded_block[245], uncoded_block[244], uncoded_block[243], uncoded_block[242], uncoded_block[241], uncoded_block[240], uncoded_block[239], uncoded_block[238], uncoded_block[237], uncoded_block[236], uncoded_block[235], uncoded_block[234], uncoded_block[233], uncoded_block[232], uncoded_block[231], uncoded_block[230], uncoded_block[229], uncoded_block[228], uncoded_block[227], uncoded_block[226], uncoded_block[225], uncoded_block[224], uncoded_block[223], uncoded_block[222], uncoded_block[221], uncoded_block[220], uncoded_block[219], uncoded_block[218], uncoded_block[217], uncoded_block[216], uncoded_block[215], uncoded_block[214], uncoded_block[213], uncoded_block[212], uncoded_block[211], uncoded_block[210], uncoded_block[209], uncoded_block[208], uncoded_block[207], uncoded_block[206], uncoded_block[205], uncoded_block[204], uncoded_block[203], uncoded_block[202], uncoded_block[201], uncoded_block[200], uncoded_block[199], uncoded_block[198], uncoded_block[197], uncoded_block[196], uncoded_block[195], uncoded_block[194], uncoded_block[193], uncoded_block[192], uncoded_block[191], uncoded_block[190], uncoded_block[189], uncoded_block[188], uncoded_block[187], uncoded_block[186], uncoded_block[185], uncoded_block[184], uncoded_block[183], uncoded_block[182], uncoded_block[181], uncoded_block[180], uncoded_block[179], uncoded_block[178], uncoded_block[177], uncoded_block[176], uncoded_block[175], uncoded_block[174], uncoded_block[173], uncoded_block[172], uncoded_block[171], uncoded_block[170], uncoded_block[169], uncoded_block[168], uncoded_block[167], uncoded_block[166], uncoded_block[165], uncoded_block[164], uncoded_block[163], uncoded_block[162], uncoded_block[161], uncoded_block[160], uncoded_block[159], uncoded_block[158], uncoded_block[157], uncoded_block[156], uncoded_block[155], uncoded_block[154], uncoded_block[153], uncoded_block[152], uncoded_block[151], uncoded_block[150], uncoded_block[149], uncoded_block[148], uncoded_block[147], uncoded_block[146], uncoded_block[145], uncoded_block[144], uncoded_block[143], uncoded_block[142], uncoded_block[141], uncoded_block[140], uncoded_block[139], uncoded_block[138], uncoded_block[137], uncoded_block[136], uncoded_block[135], uncoded_block[134], uncoded_block[133], uncoded_block[132], uncoded_block[131], uncoded_block[130], uncoded_block[129], uncoded_block[128], uncoded_block[127], uncoded_block[126], uncoded_block[125], uncoded_block[124], uncoded_block[123], uncoded_block[122], uncoded_block[121], uncoded_block[120], uncoded_block[119], uncoded_block[118], uncoded_block[117], uncoded_block[116], uncoded_block[115], uncoded_block[114], uncoded_block[113], uncoded_block[112], uncoded_block[111], uncoded_block[110], uncoded_block[109], uncoded_block[108], uncoded_block[107], uncoded_block[106], uncoded_block[105], uncoded_block[104], uncoded_block[103], uncoded_block[102], uncoded_block[101], uncoded_block[100], uncoded_block[99], uncoded_block[98], uncoded_block[97], uncoded_block[96], uncoded_block[95], uncoded_block[94], uncoded_block[93], uncoded_block[92], uncoded_block[91], uncoded_block[90], uncoded_block[89], uncoded_block[88], uncoded_block[87], uncoded_block[86], uncoded_block[85], uncoded_block[84], uncoded_block[83], uncoded_block[82], uncoded_block[81], uncoded_block[80], uncoded_block[79], uncoded_block[78], uncoded_block[77], uncoded_block[76], uncoded_block[75], uncoded_block[74], uncoded_block[73], uncoded_block[72], uncoded_block[71], uncoded_block[70], uncoded_block[69], uncoded_block[68], uncoded_block[67], uncoded_block[66], uncoded_block[65], uncoded_block[64], uncoded_block[63], uncoded_block[62], uncoded_block[61], uncoded_block[60], uncoded_block[59], uncoded_block[58], uncoded_block[57], uncoded_block[56], uncoded_block[55], uncoded_block[54], uncoded_block[53], uncoded_block[52], uncoded_block[51], uncoded_block[50], uncoded_block[49], uncoded_block[48], uncoded_block[47], uncoded_block[46], uncoded_block[45], uncoded_block[44], uncoded_block[43], uncoded_block[42], uncoded_block[41], uncoded_block[40], uncoded_block[39], uncoded_block[38], uncoded_block[37], uncoded_block[36], uncoded_block[35], uncoded_block[34], uncoded_block[33], uncoded_block[32], uncoded_block[31], uncoded_block[30], uncoded_block[29], uncoded_block[28], uncoded_block[27], uncoded_block[26], uncoded_block[25], uncoded_block[24], uncoded_block[23], uncoded_block[22], uncoded_block[21], uncoded_block[20], uncoded_block[19], uncoded_block[18], uncoded_block[17], uncoded_block[16], uncoded_block[15], uncoded_block[14], uncoded_block[13], uncoded_block[12], uncoded_block[11], uncoded_block[10], uncoded_block[9], uncoded_block[8], uncoded_block[7], uncoded_block[6], uncoded_block[5], uncoded_block[4], uncoded_block[3], uncoded_block[2], uncoded_block[1], uncoded_block[0]};
endmodule
