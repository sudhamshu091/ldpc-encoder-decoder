module ldpc_decoder
  ( reset
  , clock
  , load
  , coded_block
  , decoded
  , decoded_block
  );
  input  reset;
  input  clock;
  input  load;
  input  [2047:0] coded_block;
  output decoded;
  output [2047:0] decoded_block;
  reg  r2047;
  reg  r2046;
  reg  r2045;
  reg  r2044;
  reg  r2043;
  reg  r2042;
  reg  r2041;
  reg  r2040;
  reg  r2039;
  reg  r2038;
  reg  r2037;
  reg  r2036;
  reg  r2035;
  reg  r2034;
  reg  r2033;
  reg  r2032;
  reg  r2031;
  reg  r2030;
  reg  r2029;
  reg  r2028;
  reg  r2027;
  reg  r2026;
  reg  r2025;
  reg  r2024;
  reg  r2023;
  reg  r2022;
  reg  r2021;
  reg  r2020;
  reg  r2019;
  reg  r2018;
  reg  r2017;
  reg  r2016;
  reg  r2015;
  reg  r2014;
  reg  r2013;
  reg  r2012;
  reg  r2011;
  reg  r2010;
  reg  r2009;
  reg  r2008;
  reg  r2007;
  reg  r2006;
  reg  r2005;
  reg  r2004;
  reg  r2003;
  reg  r2002;
  reg  r2001;
  reg  r2000;
  reg  r1999;
  reg  r1998;
  reg  r1997;
  reg  r1996;
  reg  r1995;
  reg  r1994;
  reg  r1993;
  reg  r1992;
  reg  r1991;
  reg  r1990;
  reg  r1989;
  reg  r1988;
  reg  r1987;
  reg  r1986;
  reg  r1985;
  reg  r1984;
  reg  r1983;
  reg  r1982;
  reg  r1981;
  reg  r1980;
  reg  r1979;
  reg  r1978;
  reg  r1977;
  reg  r1976;
  reg  r1975;
  reg  r1974;
  reg  r1973;
  reg  r1972;
  reg  r1971;
  reg  r1970;
  reg  r1969;
  reg  r1968;
  reg  r1967;
  reg  r1966;
  reg  r1965;
  reg  r1964;
  reg  r1963;
  reg  r1962;
  reg  r1961;
  reg  r1960;
  reg  r1959;
  reg  r1958;
  reg  r1957;
  reg  r1956;
  reg  r1955;
  reg  r1954;
  reg  r1953;
  reg  r1952;
  reg  r1951;
  reg  r1950;
  reg  r1949;
  reg  r1948;
  reg  r1947;
  reg  r1946;
  reg  r1945;
  reg  r1944;
  reg  r1943;
  reg  r1942;
  reg  r1941;
  reg  r1940;
  reg  r1939;
  reg  r1938;
  reg  r1937;
  reg  r1936;
  reg  r1935;
  reg  r1934;
  reg  r1933;
  reg  r1932;
  reg  r1931;
  reg  r1930;
  reg  r1929;
  reg  r1928;
  reg  r1927;
  reg  r1926;
  reg  r1925;
  reg  r1924;
  reg  r1923;
  reg  r1922;
  reg  r1921;
  reg  r1920;
  reg  r1919;
  reg  r1918;
  reg  r1917;
  reg  r1916;
  reg  r1915;
  reg  r1914;
  reg  r1913;
  reg  r1912;
  reg  r1911;
  reg  r1910;
  reg  r1909;
  reg  r1908;
  reg  r1907;
  reg  r1906;
  reg  r1905;
  reg  r1904;
  reg  r1903;
  reg  r1902;
  reg  r1901;
  reg  r1900;
  reg  r1899;
  reg  r1898;
  reg  r1897;
  reg  r1896;
  reg  r1895;
  reg  r1894;
  reg  r1893;
  reg  r1892;
  reg  r1891;
  reg  r1890;
  reg  r1889;
  reg  r1888;
  reg  r1887;
  reg  r1886;
  reg  r1885;
  reg  r1884;
  reg  r1883;
  reg  r1882;
  reg  r1881;
  reg  r1880;
  reg  r1879;
  reg  r1878;
  reg  r1877;
  reg  r1876;
  reg  r1875;
  reg  r1874;
  reg  r1873;
  reg  r1872;
  reg  r1871;
  reg  r1870;
  reg  r1869;
  reg  r1868;
  reg  r1867;
  reg  r1866;
  reg  r1865;
  reg  r1864;
  reg  r1863;
  reg  r1862;
  reg  r1861;
  reg  r1860;
  reg  r1859;
  reg  r1858;
  reg  r1857;
  reg  r1856;
  reg  r1855;
  reg  r1854;
  reg  r1853;
  reg  r1852;
  reg  r1851;
  reg  r1850;
  reg  r1849;
  reg  r1848;
  reg  r1847;
  reg  r1846;
  reg  r1845;
  reg  r1844;
  reg  r1843;
  reg  r1842;
  reg  r1841;
  reg  r1840;
  reg  r1839;
  reg  r1838;
  reg  r1837;
  reg  r1836;
  reg  r1835;
  reg  r1834;
  reg  r1833;
  reg  r1832;
  reg  r1831;
  reg  r1830;
  reg  r1829;
  reg  r1828;
  reg  r1827;
  reg  r1826;
  reg  r1825;
  reg  r1824;
  reg  r1823;
  reg  r1822;
  reg  r1821;
  reg  r1820;
  reg  r1819;
  reg  r1818;
  reg  r1817;
  reg  r1816;
  reg  r1815;
  reg  r1814;
  reg  r1813;
  reg  r1812;
  reg  r1811;
  reg  r1810;
  reg  r1809;
  reg  r1808;
  reg  r1807;
  reg  r1806;
  reg  r1805;
  reg  r1804;
  reg  r1803;
  reg  r1802;
  reg  r1801;
  reg  r1800;
  reg  r1799;
  reg  r1798;
  reg  r1797;
  reg  r1796;
  reg  r1795;
  reg  r1794;
  reg  r1793;
  reg  r1792;
  reg  r1791;
  reg  r1790;
  reg  r1789;
  reg  r1788;
  reg  r1787;
  reg  r1786;
  reg  r1785;
  reg  r1784;
  reg  r1783;
  reg  r1782;
  reg  r1781;
  reg  r1780;
  reg  r1779;
  reg  r1778;
  reg  r1777;
  reg  r1776;
  reg  r1775;
  reg  r1774;
  reg  r1773;
  reg  r1772;
  reg  r1771;
  reg  r1770;
  reg  r1769;
  reg  r1768;
  reg  r1767;
  reg  r1766;
  reg  r1765;
  reg  r1764;
  reg  r1763;
  reg  r1762;
  reg  r1761;
  reg  r1760;
  reg  r1759;
  reg  r1758;
  reg  r1757;
  reg  r1756;
  reg  r1755;
  reg  r1754;
  reg  r1753;
  reg  r1752;
  reg  r1751;
  reg  r1750;
  reg  r1749;
  reg  r1748;
  reg  r1747;
  reg  r1746;
  reg  r1745;
  reg  r1744;
  reg  r1743;
  reg  r1742;
  reg  r1741;
  reg  r1740;
  reg  r1739;
  reg  r1738;
  reg  r1737;
  reg  r1736;
  reg  r1735;
  reg  r1734;
  reg  r1733;
  reg  r1732;
  reg  r1731;
  reg  r1730;
  reg  r1729;
  reg  r1728;
  reg  r1727;
  reg  r1726;
  reg  r1725;
  reg  r1724;
  reg  r1723;
  reg  r1722;
  reg  r1721;
  reg  r1720;
  reg  r1719;
  reg  r1718;
  reg  r1717;
  reg  r1716;
  reg  r1715;
  reg  r1714;
  reg  r1713;
  reg  r1712;
  reg  r1711;
  reg  r1710;
  reg  r1709;
  reg  r1708;
  reg  r1707;
  reg  r1706;
  reg  r1705;
  reg  r1704;
  reg  r1703;
  reg  r1702;
  reg  r1701;
  reg  r1700;
  reg  r1699;
  reg  r1698;
  reg  r1697;
  reg  r1696;
  reg  r1695;
  reg  r1694;
  reg  r1693;
  reg  r1692;
  reg  r1691;
  reg  r1690;
  reg  r1689;
  reg  r1688;
  reg  r1687;
  reg  r1686;
  reg  r1685;
  reg  r1684;
  reg  r1683;
  reg  r1682;
  reg  r1681;
  reg  r1680;
  reg  r1679;
  reg  r1678;
  reg  r1677;
  reg  r1676;
  reg  r1675;
  reg  r1674;
  reg  r1673;
  reg  r1672;
  reg  r1671;
  reg  r1670;
  reg  r1669;
  reg  r1668;
  reg  r1667;
  reg  r1666;
  reg  r1665;
  reg  r1664;
  reg  r1663;
  reg  r1662;
  reg  r1661;
  reg  r1660;
  reg  r1659;
  reg  r1658;
  reg  r1657;
  reg  r1656;
  reg  r1655;
  reg  r1654;
  reg  r1653;
  reg  r1652;
  reg  r1651;
  reg  r1650;
  reg  r1649;
  reg  r1648;
  reg  r1647;
  reg  r1646;
  reg  r1645;
  reg  r1644;
  reg  r1643;
  reg  r1642;
  reg  r1641;
  reg  r1640;
  reg  r1639;
  reg  r1638;
  reg  r1637;
  reg  r1636;
  reg  r1635;
  reg  r1634;
  reg  r1633;
  reg  r1632;
  reg  r1631;
  reg  r1630;
  reg  r1629;
  reg  r1628;
  reg  r1627;
  reg  r1626;
  reg  r1625;
  reg  r1624;
  reg  r1623;
  reg  r1622;
  reg  r1621;
  reg  r1620;
  reg  r1619;
  reg  r1618;
  reg  r1617;
  reg  r1616;
  reg  r1615;
  reg  r1614;
  reg  r1613;
  reg  r1612;
  reg  r1611;
  reg  r1610;
  reg  r1609;
  reg  r1608;
  reg  r1607;
  reg  r1606;
  reg  r1605;
  reg  r1604;
  reg  r1603;
  reg  r1602;
  reg  r1601;
  reg  r1600;
  reg  r1599;
  reg  r1598;
  reg  r1597;
  reg  r1596;
  reg  r1595;
  reg  r1594;
  reg  r1593;
  reg  r1592;
  reg  r1591;
  reg  r1590;
  reg  r1589;
  reg  r1588;
  reg  r1587;
  reg  r1586;
  reg  r1585;
  reg  r1584;
  reg  r1583;
  reg  r1582;
  reg  r1581;
  reg  r1580;
  reg  r1579;
  reg  r1578;
  reg  r1577;
  reg  r1576;
  reg  r1575;
  reg  r1574;
  reg  r1573;
  reg  r1572;
  reg  r1571;
  reg  r1570;
  reg  r1569;
  reg  r1568;
  reg  r1567;
  reg  r1566;
  reg  r1565;
  reg  r1564;
  reg  r1563;
  reg  r1562;
  reg  r1561;
  reg  r1560;
  reg  r1559;
  reg  r1558;
  reg  r1557;
  reg  r1556;
  reg  r1555;
  reg  r1554;
  reg  r1553;
  reg  r1552;
  reg  r1551;
  reg  r1550;
  reg  r1549;
  reg  r1548;
  reg  r1547;
  reg  r1546;
  reg  r1545;
  reg  r1544;
  reg  r1543;
  reg  r1542;
  reg  r1541;
  reg  r1540;
  reg  r1539;
  reg  r1538;
  reg  r1537;
  reg  r1536;
  reg  r1535;
  reg  r1534;
  reg  r1533;
  reg  r1532;
  reg  r1531;
  reg  r1530;
  reg  r1529;
  reg  r1528;
  reg  r1527;
  reg  r1526;
  reg  r1525;
  reg  r1524;
  reg  r1523;
  reg  r1522;
  reg  r1521;
  reg  r1520;
  reg  r1519;
  reg  r1518;
  reg  r1517;
  reg  r1516;
  reg  r1515;
  reg  r1514;
  reg  r1513;
  reg  r1512;
  reg  r1511;
  reg  r1510;
  reg  r1509;
  reg  r1508;
  reg  r1507;
  reg  r1506;
  reg  r1505;
  reg  r1504;
  reg  r1503;
  reg  r1502;
  reg  r1501;
  reg  r1500;
  reg  r1499;
  reg  r1498;
  reg  r1497;
  reg  r1496;
  reg  r1495;
  reg  r1494;
  reg  r1493;
  reg  r1492;
  reg  r1491;
  reg  r1490;
  reg  r1489;
  reg  r1488;
  reg  r1487;
  reg  r1486;
  reg  r1485;
  reg  r1484;
  reg  r1483;
  reg  r1482;
  reg  r1481;
  reg  r1480;
  reg  r1479;
  reg  r1478;
  reg  r1477;
  reg  r1476;
  reg  r1475;
  reg  r1474;
  reg  r1473;
  reg  r1472;
  reg  r1471;
  reg  r1470;
  reg  r1469;
  reg  r1468;
  reg  r1467;
  reg  r1466;
  reg  r1465;
  reg  r1464;
  reg  r1463;
  reg  r1462;
  reg  r1461;
  reg  r1460;
  reg  r1459;
  reg  r1458;
  reg  r1457;
  reg  r1456;
  reg  r1455;
  reg  r1454;
  reg  r1453;
  reg  r1452;
  reg  r1451;
  reg  r1450;
  reg  r1449;
  reg  r1448;
  reg  r1447;
  reg  r1446;
  reg  r1445;
  reg  r1444;
  reg  r1443;
  reg  r1442;
  reg  r1441;
  reg  r1440;
  reg  r1439;
  reg  r1438;
  reg  r1437;
  reg  r1436;
  reg  r1435;
  reg  r1434;
  reg  r1433;
  reg  r1432;
  reg  r1431;
  reg  r1430;
  reg  r1429;
  reg  r1428;
  reg  r1427;
  reg  r1426;
  reg  r1425;
  reg  r1424;
  reg  r1423;
  reg  r1422;
  reg  r1421;
  reg  r1420;
  reg  r1419;
  reg  r1418;
  reg  r1417;
  reg  r1416;
  reg  r1415;
  reg  r1414;
  reg  r1413;
  reg  r1412;
  reg  r1411;
  reg  r1410;
  reg  r1409;
  reg  r1408;
  reg  r1407;
  reg  r1406;
  reg  r1405;
  reg  r1404;
  reg  r1403;
  reg  r1402;
  reg  r1401;
  reg  r1400;
  reg  r1399;
  reg  r1398;
  reg  r1397;
  reg  r1396;
  reg  r1395;
  reg  r1394;
  reg  r1393;
  reg  r1392;
  reg  r1391;
  reg  r1390;
  reg  r1389;
  reg  r1388;
  reg  r1387;
  reg  r1386;
  reg  r1385;
  reg  r1384;
  reg  r1383;
  reg  r1382;
  reg  r1381;
  reg  r1380;
  reg  r1379;
  reg  r1378;
  reg  r1377;
  reg  r1376;
  reg  r1375;
  reg  r1374;
  reg  r1373;
  reg  r1372;
  reg  r1371;
  reg  r1370;
  reg  r1369;
  reg  r1368;
  reg  r1367;
  reg  r1366;
  reg  r1365;
  reg  r1364;
  reg  r1363;
  reg  r1362;
  reg  r1361;
  reg  r1360;
  reg  r1359;
  reg  r1358;
  reg  r1357;
  reg  r1356;
  reg  r1355;
  reg  r1354;
  reg  r1353;
  reg  r1352;
  reg  r1351;
  reg  r1350;
  reg  r1349;
  reg  r1348;
  reg  r1347;
  reg  r1346;
  reg  r1345;
  reg  r1344;
  reg  r1343;
  reg  r1342;
  reg  r1341;
  reg  r1340;
  reg  r1339;
  reg  r1338;
  reg  r1337;
  reg  r1336;
  reg  r1335;
  reg  r1334;
  reg  r1333;
  reg  r1332;
  reg  r1331;
  reg  r1330;
  reg  r1329;
  reg  r1328;
  reg  r1327;
  reg  r1326;
  reg  r1325;
  reg  r1324;
  reg  r1323;
  reg  r1322;
  reg  r1321;
  reg  r1320;
  reg  r1319;
  reg  r1318;
  reg  r1317;
  reg  r1316;
  reg  r1315;
  reg  r1314;
  reg  r1313;
  reg  r1312;
  reg  r1311;
  reg  r1310;
  reg  r1309;
  reg  r1308;
  reg  r1307;
  reg  r1306;
  reg  r1305;
  reg  r1304;
  reg  r1303;
  reg  r1302;
  reg  r1301;
  reg  r1300;
  reg  r1299;
  reg  r1298;
  reg  r1297;
  reg  r1296;
  reg  r1295;
  reg  r1294;
  reg  r1293;
  reg  r1292;
  reg  r1291;
  reg  r1290;
  reg  r1289;
  reg  r1288;
  reg  r1287;
  reg  r1286;
  reg  r1285;
  reg  r1284;
  reg  r1283;
  reg  r1282;
  reg  r1281;
  reg  r1280;
  reg  r1279;
  reg  r1278;
  reg  r1277;
  reg  r1276;
  reg  r1275;
  reg  r1274;
  reg  r1273;
  reg  r1272;
  reg  r1271;
  reg  r1270;
  reg  r1269;
  reg  r1268;
  reg  r1267;
  reg  r1266;
  reg  r1265;
  reg  r1264;
  reg  r1263;
  reg  r1262;
  reg  r1261;
  reg  r1260;
  reg  r1259;
  reg  r1258;
  reg  r1257;
  reg  r1256;
  reg  r1255;
  reg  r1254;
  reg  r1253;
  reg  r1252;
  reg  r1251;
  reg  r1250;
  reg  r1249;
  reg  r1248;
  reg  r1247;
  reg  r1246;
  reg  r1245;
  reg  r1244;
  reg  r1243;
  reg  r1242;
  reg  r1241;
  reg  r1240;
  reg  r1239;
  reg  r1238;
  reg  r1237;
  reg  r1236;
  reg  r1235;
  reg  r1234;
  reg  r1233;
  reg  r1232;
  reg  r1231;
  reg  r1230;
  reg  r1229;
  reg  r1228;
  reg  r1227;
  reg  r1226;
  reg  r1225;
  reg  r1224;
  reg  r1223;
  reg  r1222;
  reg  r1221;
  reg  r1220;
  reg  r1219;
  reg  r1218;
  reg  r1217;
  reg  r1216;
  reg  r1215;
  reg  r1214;
  reg  r1213;
  reg  r1212;
  reg  r1211;
  reg  r1210;
  reg  r1209;
  reg  r1208;
  reg  r1207;
  reg  r1206;
  reg  r1205;
  reg  r1204;
  reg  r1203;
  reg  r1202;
  reg  r1201;
  reg  r1200;
  reg  r1199;
  reg  r1198;
  reg  r1197;
  reg  r1196;
  reg  r1195;
  reg  r1194;
  reg  r1193;
  reg  r1192;
  reg  r1191;
  reg  r1190;
  reg  r1189;
  reg  r1188;
  reg  r1187;
  reg  r1186;
  reg  r1185;
  reg  r1184;
  reg  r1183;
  reg  r1182;
  reg  r1181;
  reg  r1180;
  reg  r1179;
  reg  r1178;
  reg  r1177;
  reg  r1176;
  reg  r1175;
  reg  r1174;
  reg  r1173;
  reg  r1172;
  reg  r1171;
  reg  r1170;
  reg  r1169;
  reg  r1168;
  reg  r1167;
  reg  r1166;
  reg  r1165;
  reg  r1164;
  reg  r1163;
  reg  r1162;
  reg  r1161;
  reg  r1160;
  reg  r1159;
  reg  r1158;
  reg  r1157;
  reg  r1156;
  reg  r1155;
  reg  r1154;
  reg  r1153;
  reg  r1152;
  reg  r1151;
  reg  r1150;
  reg  r1149;
  reg  r1148;
  reg  r1147;
  reg  r1146;
  reg  r1145;
  reg  r1144;
  reg  r1143;
  reg  r1142;
  reg  r1141;
  reg  r1140;
  reg  r1139;
  reg  r1138;
  reg  r1137;
  reg  r1136;
  reg  r1135;
  reg  r1134;
  reg  r1133;
  reg  r1132;
  reg  r1131;
  reg  r1130;
  reg  r1129;
  reg  r1128;
  reg  r1127;
  reg  r1126;
  reg  r1125;
  reg  r1124;
  reg  r1123;
  reg  r1122;
  reg  r1121;
  reg  r1120;
  reg  r1119;
  reg  r1118;
  reg  r1117;
  reg  r1116;
  reg  r1115;
  reg  r1114;
  reg  r1113;
  reg  r1112;
  reg  r1111;
  reg  r1110;
  reg  r1109;
  reg  r1108;
  reg  r1107;
  reg  r1106;
  reg  r1105;
  reg  r1104;
  reg  r1103;
  reg  r1102;
  reg  r1101;
  reg  r1100;
  reg  r1099;
  reg  r1098;
  reg  r1097;
  reg  r1096;
  reg  r1095;
  reg  r1094;
  reg  r1093;
  reg  r1092;
  reg  r1091;
  reg  r1090;
  reg  r1089;
  reg  r1088;
  reg  r1087;
  reg  r1086;
  reg  r1085;
  reg  r1084;
  reg  r1083;
  reg  r1082;
  reg  r1081;
  reg  r1080;
  reg  r1079;
  reg  r1078;
  reg  r1077;
  reg  r1076;
  reg  r1075;
  reg  r1074;
  reg  r1073;
  reg  r1072;
  reg  r1071;
  reg  r1070;
  reg  r1069;
  reg  r1068;
  reg  r1067;
  reg  r1066;
  reg  r1065;
  reg  r1064;
  reg  r1063;
  reg  r1062;
  reg  r1061;
  reg  r1060;
  reg  r1059;
  reg  r1058;
  reg  r1057;
  reg  r1056;
  reg  r1055;
  reg  r1054;
  reg  r1053;
  reg  r1052;
  reg  r1051;
  reg  r1050;
  reg  r1049;
  reg  r1048;
  reg  r1047;
  reg  r1046;
  reg  r1045;
  reg  r1044;
  reg  r1043;
  reg  r1042;
  reg  r1041;
  reg  r1040;
  reg  r1039;
  reg  r1038;
  reg  r1037;
  reg  r1036;
  reg  r1035;
  reg  r1034;
  reg  r1033;
  reg  r1032;
  reg  r1031;
  reg  r1030;
  reg  r1029;
  reg  r1028;
  reg  r1027;
  reg  r1026;
  reg  r1025;
  reg  r1024;
  reg  r1023;
  reg  r1022;
  reg  r1021;
  reg  r1020;
  reg  r1019;
  reg  r1018;
  reg  r1017;
  reg  r1016;
  reg  r1015;
  reg  r1014;
  reg  r1013;
  reg  r1012;
  reg  r1011;
  reg  r1010;
  reg  r1009;
  reg  r1008;
  reg  r1007;
  reg  r1006;
  reg  r1005;
  reg  r1004;
  reg  r1003;
  reg  r1002;
  reg  r1001;
  reg  r1000;
  reg  r999;
  reg  r998;
  reg  r997;
  reg  r996;
  reg  r995;
  reg  r994;
  reg  r993;
  reg  r992;
  reg  r991;
  reg  r990;
  reg  r989;
  reg  r988;
  reg  r987;
  reg  r986;
  reg  r985;
  reg  r984;
  reg  r983;
  reg  r982;
  reg  r981;
  reg  r980;
  reg  r979;
  reg  r978;
  reg  r977;
  reg  r976;
  reg  r975;
  reg  r974;
  reg  r973;
  reg  r972;
  reg  r971;
  reg  r970;
  reg  r969;
  reg  r968;
  reg  r967;
  reg  r966;
  reg  r965;
  reg  r964;
  reg  r963;
  reg  r962;
  reg  r961;
  reg  r960;
  reg  r959;
  reg  r958;
  reg  r957;
  reg  r956;
  reg  r955;
  reg  r954;
  reg  r953;
  reg  r952;
  reg  r951;
  reg  r950;
  reg  r949;
  reg  r948;
  reg  r947;
  reg  r946;
  reg  r945;
  reg  r944;
  reg  r943;
  reg  r942;
  reg  r941;
  reg  r940;
  reg  r939;
  reg  r938;
  reg  r937;
  reg  r936;
  reg  r935;
  reg  r934;
  reg  r933;
  reg  r932;
  reg  r931;
  reg  r930;
  reg  r929;
  reg  r928;
  reg  r927;
  reg  r926;
  reg  r925;
  reg  r924;
  reg  r923;
  reg  r922;
  reg  r921;
  reg  r920;
  reg  r919;
  reg  r918;
  reg  r917;
  reg  r916;
  reg  r915;
  reg  r914;
  reg  r913;
  reg  r912;
  reg  r911;
  reg  r910;
  reg  r909;
  reg  r908;
  reg  r907;
  reg  r906;
  reg  r905;
  reg  r904;
  reg  r903;
  reg  r902;
  reg  r901;
  reg  r900;
  reg  r899;
  reg  r898;
  reg  r897;
  reg  r896;
  reg  r895;
  reg  r894;
  reg  r893;
  reg  r892;
  reg  r891;
  reg  r890;
  reg  r889;
  reg  r888;
  reg  r887;
  reg  r886;
  reg  r885;
  reg  r884;
  reg  r883;
  reg  r882;
  reg  r881;
  reg  r880;
  reg  r879;
  reg  r878;
  reg  r877;
  reg  r876;
  reg  r875;
  reg  r874;
  reg  r873;
  reg  r872;
  reg  r871;
  reg  r870;
  reg  r869;
  reg  r868;
  reg  r867;
  reg  r866;
  reg  r865;
  reg  r864;
  reg  r863;
  reg  r862;
  reg  r861;
  reg  r860;
  reg  r859;
  reg  r858;
  reg  r857;
  reg  r856;
  reg  r855;
  reg  r854;
  reg  r853;
  reg  r852;
  reg  r851;
  reg  r850;
  reg  r849;
  reg  r848;
  reg  r847;
  reg  r846;
  reg  r845;
  reg  r844;
  reg  r843;
  reg  r842;
  reg  r841;
  reg  r840;
  reg  r839;
  reg  r838;
  reg  r837;
  reg  r836;
  reg  r835;
  reg  r834;
  reg  r833;
  reg  r832;
  reg  r831;
  reg  r830;
  reg  r829;
  reg  r828;
  reg  r827;
  reg  r826;
  reg  r825;
  reg  r824;
  reg  r823;
  reg  r822;
  reg  r821;
  reg  r820;
  reg  r819;
  reg  r818;
  reg  r817;
  reg  r816;
  reg  r815;
  reg  r814;
  reg  r813;
  reg  r812;
  reg  r811;
  reg  r810;
  reg  r809;
  reg  r808;
  reg  r807;
  reg  r806;
  reg  r805;
  reg  r804;
  reg  r803;
  reg  r802;
  reg  r801;
  reg  r800;
  reg  r799;
  reg  r798;
  reg  r797;
  reg  r796;
  reg  r795;
  reg  r794;
  reg  r793;
  reg  r792;
  reg  r791;
  reg  r790;
  reg  r789;
  reg  r788;
  reg  r787;
  reg  r786;
  reg  r785;
  reg  r784;
  reg  r783;
  reg  r782;
  reg  r781;
  reg  r780;
  reg  r779;
  reg  r778;
  reg  r777;
  reg  r776;
  reg  r775;
  reg  r774;
  reg  r773;
  reg  r772;
  reg  r771;
  reg  r770;
  reg  r769;
  reg  r768;
  reg  r767;
  reg  r766;
  reg  r765;
  reg  r764;
  reg  r763;
  reg  r762;
  reg  r761;
  reg  r760;
  reg  r759;
  reg  r758;
  reg  r757;
  reg  r756;
  reg  r755;
  reg  r754;
  reg  r753;
  reg  r752;
  reg  r751;
  reg  r750;
  reg  r749;
  reg  r748;
  reg  r747;
  reg  r746;
  reg  r745;
  reg  r744;
  reg  r743;
  reg  r742;
  reg  r741;
  reg  r740;
  reg  r739;
  reg  r738;
  reg  r737;
  reg  r736;
  reg  r735;
  reg  r734;
  reg  r733;
  reg  r732;
  reg  r731;
  reg  r730;
  reg  r729;
  reg  r728;
  reg  r727;
  reg  r726;
  reg  r725;
  reg  r724;
  reg  r723;
  reg  r722;
  reg  r721;
  reg  r720;
  reg  r719;
  reg  r718;
  reg  r717;
  reg  r716;
  reg  r715;
  reg  r714;
  reg  r713;
  reg  r712;
  reg  r711;
  reg  r710;
  reg  r709;
  reg  r708;
  reg  r707;
  reg  r706;
  reg  r705;
  reg  r704;
  reg  r703;
  reg  r702;
  reg  r701;
  reg  r700;
  reg  r699;
  reg  r698;
  reg  r697;
  reg  r696;
  reg  r695;
  reg  r694;
  reg  r693;
  reg  r692;
  reg  r691;
  reg  r690;
  reg  r689;
  reg  r688;
  reg  r687;
  reg  r686;
  reg  r685;
  reg  r684;
  reg  r683;
  reg  r682;
  reg  r681;
  reg  r680;
  reg  r679;
  reg  r678;
  reg  r677;
  reg  r676;
  reg  r675;
  reg  r674;
  reg  r673;
  reg  r672;
  reg  r671;
  reg  r670;
  reg  r669;
  reg  r668;
  reg  r667;
  reg  r666;
  reg  r665;
  reg  r664;
  reg  r663;
  reg  r662;
  reg  r661;
  reg  r660;
  reg  r659;
  reg  r658;
  reg  r657;
  reg  r656;
  reg  r655;
  reg  r654;
  reg  r653;
  reg  r652;
  reg  r651;
  reg  r650;
  reg  r649;
  reg  r648;
  reg  r647;
  reg  r646;
  reg  r645;
  reg  r644;
  reg  r643;
  reg  r642;
  reg  r641;
  reg  r640;
  reg  r639;
  reg  r638;
  reg  r637;
  reg  r636;
  reg  r635;
  reg  r634;
  reg  r633;
  reg  r632;
  reg  r631;
  reg  r630;
  reg  r629;
  reg  r628;
  reg  r627;
  reg  r626;
  reg  r625;
  reg  r624;
  reg  r623;
  reg  r622;
  reg  r621;
  reg  r620;
  reg  r619;
  reg  r618;
  reg  r617;
  reg  r616;
  reg  r615;
  reg  r614;
  reg  r613;
  reg  r612;
  reg  r611;
  reg  r610;
  reg  r609;
  reg  r608;
  reg  r607;
  reg  r606;
  reg  r605;
  reg  r604;
  reg  r603;
  reg  r602;
  reg  r601;
  reg  r600;
  reg  r599;
  reg  r598;
  reg  r597;
  reg  r596;
  reg  r595;
  reg  r594;
  reg  r593;
  reg  r592;
  reg  r591;
  reg  r590;
  reg  r589;
  reg  r588;
  reg  r587;
  reg  r586;
  reg  r585;
  reg  r584;
  reg  r583;
  reg  r582;
  reg  r581;
  reg  r580;
  reg  r579;
  reg  r578;
  reg  r577;
  reg  r576;
  reg  r575;
  reg  r574;
  reg  r573;
  reg  r572;
  reg  r571;
  reg  r570;
  reg  r569;
  reg  r568;
  reg  r567;
  reg  r566;
  reg  r565;
  reg  r564;
  reg  r563;
  reg  r562;
  reg  r561;
  reg  r560;
  reg  r559;
  reg  r558;
  reg  r557;
  reg  r556;
  reg  r555;
  reg  r554;
  reg  r553;
  reg  r552;
  reg  r551;
  reg  r550;
  reg  r549;
  reg  r548;
  reg  r547;
  reg  r546;
  reg  r545;
  reg  r544;
  reg  r543;
  reg  r542;
  reg  r541;
  reg  r540;
  reg  r539;
  reg  r538;
  reg  r537;
  reg  r536;
  reg  r535;
  reg  r534;
  reg  r533;
  reg  r532;
  reg  r531;
  reg  r530;
  reg  r529;
  reg  r528;
  reg  r527;
  reg  r526;
  reg  r525;
  reg  r524;
  reg  r523;
  reg  r522;
  reg  r521;
  reg  r520;
  reg  r519;
  reg  r518;
  reg  r517;
  reg  r516;
  reg  r515;
  reg  r514;
  reg  r513;
  reg  r512;
  reg  r511;
  reg  r510;
  reg  r509;
  reg  r508;
  reg  r507;
  reg  r506;
  reg  r505;
  reg  r504;
  reg  r503;
  reg  r502;
  reg  r501;
  reg  r500;
  reg  r499;
  reg  r498;
  reg  r497;
  reg  r496;
  reg  r495;
  reg  r494;
  reg  r493;
  reg  r492;
  reg  r491;
  reg  r490;
  reg  r489;
  reg  r488;
  reg  r487;
  reg  r486;
  reg  r485;
  reg  r484;
  reg  r483;
  reg  r482;
  reg  r481;
  reg  r480;
  reg  r479;
  reg  r478;
  reg  r477;
  reg  r476;
  reg  r475;
  reg  r474;
  reg  r473;
  reg  r472;
  reg  r471;
  reg  r470;
  reg  r469;
  reg  r468;
  reg  r467;
  reg  r466;
  reg  r465;
  reg  r464;
  reg  r463;
  reg  r462;
  reg  r461;
  reg  r460;
  reg  r459;
  reg  r458;
  reg  r457;
  reg  r456;
  reg  r455;
  reg  r454;
  reg  r453;
  reg  r452;
  reg  r451;
  reg  r450;
  reg  r449;
  reg  r448;
  reg  r447;
  reg  r446;
  reg  r445;
  reg  r444;
  reg  r443;
  reg  r442;
  reg  r441;
  reg  r440;
  reg  r439;
  reg  r438;
  reg  r437;
  reg  r436;
  reg  r435;
  reg  r434;
  reg  r433;
  reg  r432;
  reg  r431;
  reg  r430;
  reg  r429;
  reg  r428;
  reg  r427;
  reg  r426;
  reg  r425;
  reg  r424;
  reg  r423;
  reg  r422;
  reg  r421;
  reg  r420;
  reg  r419;
  reg  r418;
  reg  r417;
  reg  r416;
  reg  r415;
  reg  r414;
  reg  r413;
  reg  r412;
  reg  r411;
  reg  r410;
  reg  r409;
  reg  r408;
  reg  r407;
  reg  r406;
  reg  r405;
  reg  r404;
  reg  r403;
  reg  r402;
  reg  r401;
  reg  r400;
  reg  r399;
  reg  r398;
  reg  r397;
  reg  r396;
  reg  r395;
  reg  r394;
  reg  r393;
  reg  r392;
  reg  r391;
  reg  r390;
  reg  r389;
  reg  r388;
  reg  r387;
  reg  r386;
  reg  r385;
  reg  r384;
  reg  r383;
  reg  r382;
  reg  r381;
  reg  r380;
  reg  r379;
  reg  r378;
  reg  r377;
  reg  r376;
  reg  r375;
  reg  r374;
  reg  r373;
  reg  r372;
  reg  r371;
  reg  r370;
  reg  r369;
  reg  r368;
  reg  r367;
  reg  r366;
  reg  r365;
  reg  r364;
  reg  r363;
  reg  r362;
  reg  r361;
  reg  r360;
  reg  r359;
  reg  r358;
  reg  r357;
  reg  r356;
  reg  r355;
  reg  r354;
  reg  r353;
  reg  r352;
  reg  r351;
  reg  r350;
  reg  r349;
  reg  r348;
  reg  r347;
  reg  r346;
  reg  r345;
  reg  r344;
  reg  r343;
  reg  r342;
  reg  r341;
  reg  r340;
  reg  r339;
  reg  r338;
  reg  r337;
  reg  r336;
  reg  r335;
  reg  r334;
  reg  r333;
  reg  r332;
  reg  r331;
  reg  r330;
  reg  r329;
  reg  r328;
  reg  r327;
  reg  r326;
  reg  r325;
  reg  r324;
  reg  r323;
  reg  r322;
  reg  r321;
  reg  r320;
  reg  r319;
  reg  r318;
  reg  r317;
  reg  r316;
  reg  r315;
  reg  r314;
  reg  r313;
  reg  r312;
  reg  r311;
  reg  r310;
  reg  r309;
  reg  r308;
  reg  r307;
  reg  r306;
  reg  r305;
  reg  r304;
  reg  r303;
  reg  r302;
  reg  r301;
  reg  r300;
  reg  r299;
  reg  r298;
  reg  r297;
  reg  r296;
  reg  r295;
  reg  r294;
  reg  r293;
  reg  r292;
  reg  r291;
  reg  r290;
  reg  r289;
  reg  r288;
  reg  r287;
  reg  r286;
  reg  r285;
  reg  r284;
  reg  r283;
  reg  r282;
  reg  r281;
  reg  r280;
  reg  r279;
  reg  r278;
  reg  r277;
  reg  r276;
  reg  r275;
  reg  r274;
  reg  r273;
  reg  r272;
  reg  r271;
  reg  r270;
  reg  r269;
  reg  r268;
  reg  r267;
  reg  r266;
  reg  r265;
  reg  r264;
  reg  r263;
  reg  r262;
  reg  r261;
  reg  r260;
  reg  r259;
  reg  r258;
  reg  r257;
  reg  r256;
  reg  r255;
  reg  r254;
  reg  r253;
  reg  r252;
  reg  r251;
  reg  r250;
  reg  r249;
  reg  r248;
  reg  r247;
  reg  r246;
  reg  r245;
  reg  r244;
  reg  r243;
  reg  r242;
  reg  r241;
  reg  r240;
  reg  r239;
  reg  r238;
  reg  r237;
  reg  r236;
  reg  r235;
  reg  r234;
  reg  r233;
  reg  r232;
  reg  r231;
  reg  r230;
  reg  r229;
  reg  r228;
  reg  r227;
  reg  r226;
  reg  r225;
  reg  r224;
  reg  r223;
  reg  r222;
  reg  r221;
  reg  r220;
  reg  r219;
  reg  r218;
  reg  r217;
  reg  r216;
  reg  r215;
  reg  r214;
  reg  r213;
  reg  r212;
  reg  r211;
  reg  r210;
  reg  r209;
  reg  r208;
  reg  r207;
  reg  r206;
  reg  r205;
  reg  r204;
  reg  r203;
  reg  r202;
  reg  r201;
  reg  r200;
  reg  r199;
  reg  r198;
  reg  r197;
  reg  r196;
  reg  r195;
  reg  r194;
  reg  r193;
  reg  r192;
  reg  r191;
  reg  r190;
  reg  r189;
  reg  r188;
  reg  r187;
  reg  r186;
  reg  r185;
  reg  r184;
  reg  r183;
  reg  r182;
  reg  r181;
  reg  r180;
  reg  r179;
  reg  r178;
  reg  r177;
  reg  r176;
  reg  r175;
  reg  r174;
  reg  r173;
  reg  r172;
  reg  r171;
  reg  r170;
  reg  r169;
  reg  r168;
  reg  r167;
  reg  r166;
  reg  r165;
  reg  r164;
  reg  r163;
  reg  r162;
  reg  r161;
  reg  r160;
  reg  r159;
  reg  r158;
  reg  r157;
  reg  r156;
  reg  r155;
  reg  r154;
  reg  r153;
  reg  r152;
  reg  r151;
  reg  r150;
  reg  r149;
  reg  r148;
  reg  r147;
  reg  r146;
  reg  r145;
  reg  r144;
  reg  r143;
  reg  r142;
  reg  r141;
  reg  r140;
  reg  r139;
  reg  r138;
  reg  r137;
  reg  r136;
  reg  r135;
  reg  r134;
  reg  r133;
  reg  r132;
  reg  r131;
  reg  r130;
  reg  r129;
  reg  r128;
  reg  r127;
  reg  r126;
  reg  r125;
  reg  r124;
  reg  r123;
  reg  r122;
  reg  r121;
  reg  r120;
  reg  r119;
  reg  r118;
  reg  r117;
  reg  r116;
  reg  r115;
  reg  r114;
  reg  r113;
  reg  r112;
  reg  r111;
  reg  r110;
  reg  r109;
  reg  r108;
  reg  r107;
  reg  r106;
  reg  r105;
  reg  r104;
  reg  r103;
  reg  r102;
  reg  r101;
  reg  r100;
  reg  r99;
  reg  r98;
  reg  r97;
  reg  r96;
  reg  r95;
  reg  r94;
  reg  r93;
  reg  r92;
  reg  r91;
  reg  r90;
  reg  r89;
  reg  r88;
  reg  r87;
  reg  r86;
  reg  r85;
  reg  r84;
  reg  r83;
  reg  r82;
  reg  r81;
  reg  r80;
  reg  r79;
  reg  r78;
  reg  r77;
  reg  r76;
  reg  r75;
  reg  r74;
  reg  r73;
  reg  r72;
  reg  r71;
  reg  r70;
  reg  r69;
  reg  r68;
  reg  r67;
  reg  r66;
  reg  r65;
  reg  r64;
  reg  r63;
  reg  r62;
  reg  r61;
  reg  r60;
  reg  r59;
  reg  r58;
  reg  r57;
  reg  r56;
  reg  r55;
  reg  r54;
  reg  r53;
  reg  r52;
  reg  r51;
  reg  r50;
  reg  r49;
  reg  r48;
  reg  r47;
  reg  r46;
  reg  r45;
  reg  r44;
  reg  r43;
  reg  r42;
  reg  r41;
  reg  r40;
  reg  r39;
  reg  r38;
  reg  r37;
  reg  r36;
  reg  r35;
  reg  r34;
  reg  r33;
  reg  r32;
  reg  r31;
  reg  r30;
  reg  r29;
  reg  r28;
  reg  r27;
  reg  r26;
  reg  r25;
  reg  r24;
  reg  r23;
  reg  r22;
  reg  r21;
  reg  r20;
  reg  r19;
  reg  r18;
  reg  r17;
  reg  r16;
  reg  r15;
  reg  r14;
  reg  r13;
  reg  r12;
  reg  r11;
  reg  r10;
  reg  r9;
  reg  r8;
  reg  r7;
  reg  r6;
  reg  r5;
  reg  r4;
  reg  r3;
  reg  r2;
  reg  r1;
  reg  r0;
  wire _0 = 1'd0;
  wire _1 = 1'd1;
  wire _2 = load & _1;
  wire _3 = _1 & _2;
  wire _4 = r53 ^ r110;
  wire _5 = r170 ^ r224;
  wire _6 = _4 ^ _5;
  wire _7 = r279 ^ r332;
  wire _8 = r447 ^ r505;
  wire _9 = _7 ^ _8;
  wire _10 = _6 ^ _9;
  wire _11 = r616 ^ r668;
  wire _12 = r1496 ^ r1497;
  wire _13 = _11 ^ _12;
  wire _14 = r1498 ^ r1499;
  wire _15 = r1500 ^ r1501;
  wire _16 = _14 ^ _15;
  wire _17 = _13 ^ _16;
  wire _18 = _10 ^ _17;
  wire _19 = r1502 ^ r1503;
  wire _20 = r1505 ^ r1509;
  wire _21 = _19 ^ _20;
  wire _22 = r1514 ^ r1519;
  wire _23 = r1525 ^ r1532;
  wire _24 = _22 ^ _23;
  wire _25 = _21 ^ _24;
  wire _26 = r1536 ^ r1552;
  wire _27 = r1575 ^ r1607;
  wire _28 = _26 ^ _27;
  wire _29 = r1648 ^ r1687;
  wire _30 = r1718 ^ r1724;
  wire _31 = _29 ^ _30;
  wire _32 = _28 ^ _31;
  wire _33 = _25 ^ _32;
  wire _34 = _18 ^ _33;
  wire _35 = r51 ^ r139;
  wire _36 = r223 ^ r241;
  wire _37 = _35 ^ _36;
  wire _38 = r307 ^ r356;
  wire _39 = r408 ^ r476;
  wire _40 = _38 ^ _39;
  wire _41 = _37 ^ _40;
  wire _42 = r515 ^ r600;
  wire _43 = r617 ^ r689;
  wire _44 = _42 ^ _43;
  wire _45 = r762 ^ r797;
  wire _46 = r854 ^ r927;
  wire _47 = _45 ^ _46;
  wire _48 = _44 ^ _47;
  wire _49 = _41 ^ _48;
  wire _50 = r990 ^ r1023;
  wire _51 = r1059 ^ r1077;
  wire _52 = _50 ^ _51;
  wire _53 = r1138 ^ r1200;
  wire _54 = r1292 ^ r1442;
  wire _55 = _53 ^ _54;
  wire _56 = _52 ^ _55;
  wire _57 = r1488 ^ r1522;
  wire _58 = r1535 ^ r1550;
  wire _59 = _57 ^ _58;
  wire _60 = r1585 ^ r1681;
  wire _61 = r1994 ^ r1996;
  wire _62 = _60 ^ _61;
  wire _63 = _59 ^ _62;
  wire _64 = _56 ^ _63;
  wire _65 = _49 ^ _64;
  wire _66 = _34 | _65;
  wire _67 = r50 ^ r92;
  wire _68 = r138 ^ r222;
  wire _69 = _67 ^ _68;
  wire _70 = r240 ^ r306;
  wire _71 = r355 ^ r407;
  wire _72 = _70 ^ _71;
  wire _73 = _69 ^ _72;
  wire _74 = r475 ^ r599;
  wire _75 = r688 ^ r761;
  wire _76 = _74 ^ _75;
  wire _77 = r853 ^ r989;
  wire _78 = r1003 ^ r1022;
  wire _79 = _77 ^ _78;
  wire _80 = _76 ^ _79;
  wire _81 = _73 ^ _80;
  wire _82 = r1076 ^ r1137;
  wire _83 = r1199 ^ r1291;
  wire _84 = _82 ^ _83;
  wire _85 = r1441 ^ r1521;
  wire _86 = r1534 ^ r1549;
  wire _87 = _85 ^ _86;
  wire _88 = _84 ^ _87;
  wire _89 = r1584 ^ r1707;
  wire _90 = r1808 ^ r1837;
  wire _91 = _89 ^ _90;
  wire _92 = r1904 ^ r1948;
  wire _93 = r2003 ^ r2007;
  wire _94 = _92 ^ _93;
  wire _95 = _91 ^ _94;
  wire _96 = _88 ^ _95;
  wire _97 = _81 ^ _96;
  wire _98 = r91 ^ r137;
  wire _99 = r221 ^ r239;
  wire _100 = _98 ^ _99;
  wire _101 = r305 ^ r474;
  wire _102 = r514 ^ r598;
  wire _103 = _101 ^ _102;
  wire _104 = _100 ^ _103;
  wire _105 = r687 ^ r760;
  wire _106 = r796 ^ r852;
  wire _107 = _105 ^ _106;
  wire _108 = r926 ^ r988;
  wire _109 = r1021 ^ r1075;
  wire _110 = _108 ^ _109;
  wire _111 = _107 ^ _110;
  wire _112 = _104 ^ _111;
  wire _113 = r1136 ^ r1290;
  wire _114 = r1440 ^ r1520;
  wire _115 = _113 ^ _114;
  wire _116 = r1533 ^ r1548;
  wire _117 = r1647 ^ r1680;
  wire _118 = _116 ^ _117;
  wire _119 = _115 ^ _118;
  wire _120 = r1801 ^ r1824;
  wire _121 = r1833 ^ r1845;
  wire _122 = _120 ^ _121;
  wire _123 = r1850 ^ r1919;
  wire _124 = r1940 ^ r1942;
  wire _125 = _123 ^ _124;
  wire _126 = _122 ^ _125;
  wire _127 = _119 ^ _126;
  wire _128 = _112 ^ _127;
  wire _129 = _97 | _128;
  wire _130 = _66 | _129;
  wire _131 = r49 ^ r90;
  wire _132 = r220 ^ r238;
  wire _133 = _131 ^ _132;
  wire _134 = r304 ^ r354;
  wire _135 = r406 ^ r473;
  wire _136 = _134 ^ _135;
  wire _137 = _133 ^ _136;
  wire _138 = r513 ^ r597;
  wire _139 = r667 ^ r686;
  wire _140 = _138 ^ _139;
  wire _141 = r759 ^ r795;
  wire _142 = r851 ^ r887;
  wire _143 = _141 ^ _142;
  wire _144 = _140 ^ _143;
  wire _145 = _137 ^ _144;
  wire _146 = r925 ^ r987;
  wire _147 = r1074 ^ r1135;
  wire _148 = _146 ^ _147;
  wire _149 = r1198 ^ r1289;
  wire _150 = r1583 ^ r1646;
  wire _151 = _149 ^ _150;
  wire _152 = _148 ^ _151;
  wire _153 = r1679 ^ r1747;
  wire _154 = r1892 ^ r1901;
  wire _155 = _153 ^ _154;
  wire _156 = r1907 ^ r1944;
  wire _157 = r1977 ^ r1978;
  wire _158 = _156 ^ _157;
  wire _159 = _155 ^ _158;
  wire _160 = _152 ^ _159;
  wire _161 = _145 ^ _160;
  wire _162 = r48 ^ r89;
  wire _163 = r136 ^ r219;
  wire _164 = _162 ^ _163;
  wire _165 = r237 ^ r303;
  wire _166 = r353 ^ r405;
  wire _167 = _165 ^ _166;
  wire _168 = _164 ^ _167;
  wire _169 = r472 ^ r512;
  wire _170 = r596 ^ r666;
  wire _171 = _169 ^ _170;
  wire _172 = r685 ^ r758;
  wire _173 = r794 ^ r830;
  wire _174 = _172 ^ _173;
  wire _175 = _171 ^ _174;
  wire _176 = _168 ^ _175;
  wire _177 = r850 ^ r924;
  wire _178 = r986 ^ r1020;
  wire _179 = _177 ^ _178;
  wire _180 = r1073 ^ r1134;
  wire _181 = r1197 ^ r1275;
  wire _182 = _180 ^ _181;
  wire _183 = _179 ^ _182;
  wire _184 = r1288 ^ r1383;
  wire _185 = r1439 ^ r1547;
  wire _186 = _184 ^ _185;
  wire _187 = r1582 ^ r1645;
  wire _188 = r1678 ^ r1725;
  wire _189 = _187 ^ _188;
  wire _190 = _186 ^ _189;
  wire _191 = _183 ^ _190;
  wire _192 = _176 ^ _191;
  wire _193 = _161 | _192;
  wire _194 = r47 ^ r88;
  wire _195 = r135 ^ r218;
  wire _196 = _194 ^ _195;
  wire _197 = r236 ^ r302;
  wire _198 = r352 ^ r404;
  wire _199 = _197 ^ _198;
  wire _200 = _196 ^ _199;
  wire _201 = r471 ^ r511;
  wire _202 = r595 ^ r665;
  wire _203 = _201 ^ _202;
  wire _204 = r684 ^ r757;
  wire _205 = r777 ^ r793;
  wire _206 = _204 ^ _205;
  wire _207 = _203 ^ _206;
  wire _208 = _200 ^ _207;
  wire _209 = r849 ^ r923;
  wire _210 = r985 ^ r1019;
  wire _211 = _209 ^ _210;
  wire _212 = r1072 ^ r1133;
  wire _213 = r1196 ^ r1274;
  wire _214 = _212 ^ _213;
  wire _215 = _211 ^ _214;
  wire _216 = r1287 ^ r1382;
  wire _217 = r1438 ^ r1546;
  wire _218 = _216 ^ _217;
  wire _219 = r1581 ^ r1644;
  wire _220 = r1706 ^ r1726;
  wire _221 = _219 ^ _220;
  wire _222 = _218 ^ _221;
  wire _223 = _215 ^ _222;
  wire _224 = _208 ^ _223;
  wire _225 = r46 ^ r87;
  wire _226 = r134 ^ r217;
  wire _227 = _225 ^ _226;
  wire _228 = r235 ^ r301;
  wire _229 = r351 ^ r403;
  wire _230 = _228 ^ _229;
  wire _231 = _227 ^ _230;
  wire _232 = r470 ^ r510;
  wire _233 = r594 ^ r664;
  wire _234 = _232 ^ _233;
  wire _235 = r683 ^ r722;
  wire _236 = r756 ^ r792;
  wire _237 = _235 ^ _236;
  wire _238 = _234 ^ _237;
  wire _239 = _231 ^ _238;
  wire _240 = r848 ^ r922;
  wire _241 = r984 ^ r1018;
  wire _242 = _240 ^ _241;
  wire _243 = r1071 ^ r1132;
  wire _244 = r1195 ^ r1273;
  wire _245 = _243 ^ _244;
  wire _246 = _242 ^ _245;
  wire _247 = r1286 ^ r1381;
  wire _248 = r1437 ^ r1545;
  wire _249 = _247 ^ _248;
  wire _250 = r1580 ^ r1677;
  wire _251 = r1705 ^ r1727;
  wire _252 = _250 ^ _251;
  wire _253 = _249 ^ _252;
  wire _254 = _246 ^ _253;
  wire _255 = _239 ^ _254;
  wire _256 = _224 | _255;
  wire _257 = _193 | _256;
  wire _258 = _130 | _257;
  wire _259 = r45 ^ r133;
  wire _260 = r216 ^ r402;
  wire _261 = _259 ^ _260;
  wire _262 = r469 ^ r593;
  wire _263 = r682 ^ r755;
  wire _264 = _262 ^ _263;
  wire _265 = _261 ^ _264;
  wire _266 = r847 ^ r983;
  wire _267 = r1017 ^ r1070;
  wire _268 = _266 ^ _267;
  wire _269 = r1131 ^ r1194;
  wire _270 = r1272 ^ r1380;
  wire _271 = _269 ^ _270;
  wire _272 = _268 ^ _271;
  wire _273 = _265 ^ _272;
  wire _274 = r1436 ^ r1544;
  wire _275 = r1643 ^ r1676;
  wire _276 = _274 ^ _275;
  wire _277 = r1788 ^ r1792;
  wire _278 = r1859 ^ r1886;
  wire _279 = _277 ^ _278;
  wire _280 = _276 ^ _279;
  wire _281 = r1891 ^ r1902;
  wire _282 = r1924 ^ r1965;
  wire _283 = _281 ^ _282;
  wire _284 = r1997 ^ r2019;
  wire _285 = r2037 ^ r2038;
  wire _286 = _284 ^ _285;
  wire _287 = _283 ^ _286;
  wire _288 = _280 ^ _287;
  wire _289 = _273 ^ _288;
  wire _290 = r44 ^ r86;
  wire _291 = r132 ^ r215;
  wire _292 = _290 ^ _291;
  wire _293 = r234 ^ r300;
  wire _294 = r350 ^ r391;
  wire _295 = _293 ^ _294;
  wire _296 = _292 ^ _295;
  wire _297 = r401 ^ r468;
  wire _298 = r509 ^ r592;
  wire _299 = _297 ^ _298;
  wire _300 = r663 ^ r681;
  wire _301 = r754 ^ r791;
  wire _302 = _300 ^ _301;
  wire _303 = _299 ^ _302;
  wire _304 = _296 ^ _303;
  wire _305 = r846 ^ r921;
  wire _306 = r982 ^ r1016;
  wire _307 = _305 ^ _306;
  wire _308 = r1069 ^ r1130;
  wire _309 = r1193 ^ r1271;
  wire _310 = _308 ^ _309;
  wire _311 = _307 ^ _310;
  wire _312 = r1285 ^ r1379;
  wire _313 = r1435 ^ r1543;
  wire _314 = _312 ^ _313;
  wire _315 = r1579 ^ r1642;
  wire _316 = r1675 ^ r1728;
  wire _317 = _315 ^ _316;
  wire _318 = _314 ^ _317;
  wire _319 = _311 ^ _318;
  wire _320 = _304 ^ _319;
  wire _321 = _289 | _320;
  wire _322 = r43 ^ r85;
  wire _323 = r131 ^ r233;
  wire _324 = _322 ^ _323;
  wire _325 = r349 ^ r467;
  wire _326 = r508 ^ r662;
  wire _327 = _325 ^ _326;
  wire _328 = _324 ^ _327;
  wire _329 = r753 ^ r790;
  wire _330 = r845 ^ r920;
  wire _331 = _329 ^ _330;
  wire _332 = r981 ^ r1015;
  wire _333 = r1270 ^ r1378;
  wire _334 = _332 ^ _333;
  wire _335 = _331 ^ _334;
  wire _336 = _328 ^ _335;
  wire _337 = r1455 ^ r1542;
  wire _338 = r1578 ^ r1641;
  wire _339 = _337 ^ _338;
  wire _340 = r1674 ^ r1704;
  wire _341 = r1830 ^ r1895;
  wire _342 = _340 ^ _341;
  wire _343 = _339 ^ _342;
  wire _344 = r1918 ^ r1971;
  wire _345 = r1981 ^ r1982;
  wire _346 = _344 ^ _345;
  wire _347 = r1993 ^ r2009;
  wire _348 = r2013 ^ r2014;
  wire _349 = _347 ^ _348;
  wire _350 = _346 ^ _349;
  wire _351 = _343 ^ _350;
  wire _352 = _336 ^ _351;
  wire _353 = r42 ^ r84;
  wire _354 = r130 ^ r214;
  wire _355 = _353 ^ _354;
  wire _356 = r232 ^ r348;
  wire _357 = r400 ^ r591;
  wire _358 = _356 ^ _357;
  wire _359 = _355 ^ _358;
  wire _360 = r661 ^ r680;
  wire _361 = r752 ^ r789;
  wire _362 = _360 ^ _361;
  wire _363 = r844 ^ r919;
  wire _364 = r1014 ^ r1068;
  wire _365 = _363 ^ _364;
  wire _366 = _362 ^ _365;
  wire _367 = _359 ^ _366;
  wire _368 = r1129 ^ r1269;
  wire _369 = r1434 ^ r1454;
  wire _370 = _368 ^ _369;
  wire _371 = r1541 ^ r1577;
  wire _372 = r1640 ^ r1673;
  wire _373 = _371 ^ _372;
  wire _374 = _370 ^ _373;
  wire _375 = r1764 ^ r1829;
  wire _376 = r1843 ^ r1860;
  wire _377 = _375 ^ _376;
  wire _378 = r1867 ^ r1914;
  wire _379 = r1946 ^ r1951;
  wire _380 = _378 ^ _379;
  wire _381 = _377 ^ _380;
  wire _382 = _374 ^ _381;
  wire _383 = _367 ^ _382;
  wire _384 = _352 | _383;
  wire _385 = _321 | _384;
  wire _386 = r41 ^ r83;
  wire _387 = r129 ^ r213;
  wire _388 = _386 ^ _387;
  wire _389 = r231 ^ r299;
  wire _390 = r347 ^ r399;
  wire _391 = _389 ^ _390;
  wire _392 = _388 ^ _391;
  wire _393 = r466 ^ r507;
  wire _394 = r590 ^ r660;
  wire _395 = _393 ^ _394;
  wire _396 = r679 ^ r751;
  wire _397 = r788 ^ r843;
  wire _398 = _396 ^ _397;
  wire _399 = _395 ^ _398;
  wire _400 = _392 ^ _399;
  wire _401 = r918 ^ r980;
  wire _402 = r1067 ^ r1128;
  wire _403 = _401 ^ _402;
  wire _404 = r1192 ^ r1268;
  wire _405 = r1284 ^ r1377;
  wire _406 = _404 ^ _405;
  wire _407 = _403 ^ _406;
  wire _408 = r1433 ^ r1453;
  wire _409 = r1487 ^ r1540;
  wire _410 = _408 ^ _409;
  wire _411 = r1639 ^ r1672;
  wire _412 = r1703 ^ r1729;
  wire _413 = _411 ^ _412;
  wire _414 = _410 ^ _413;
  wire _415 = _407 ^ _414;
  wire _416 = _400 ^ _415;
  wire _417 = r82 ^ r128;
  wire _418 = r212 ^ r230;
  wire _419 = _417 ^ _418;
  wire _420 = r298 ^ r346;
  wire _421 = r398 ^ r465;
  wire _422 = _420 ^ _421;
  wire _423 = _419 ^ _422;
  wire _424 = r506 ^ r589;
  wire _425 = r659 ^ r678;
  wire _426 = _424 ^ _425;
  wire _427 = r750 ^ r787;
  wire _428 = r842 ^ r917;
  wire _429 = _427 ^ _428;
  wire _430 = _426 ^ _429;
  wire _431 = _423 ^ _430;
  wire _432 = r979 ^ r1013;
  wire _433 = r1066 ^ r1127;
  wire _434 = _432 ^ _433;
  wire _435 = r1191 ^ r1267;
  wire _436 = r1283 ^ r1376;
  wire _437 = _435 ^ _436;
  wire _438 = _434 ^ _437;
  wire _439 = r1432 ^ r1452;
  wire _440 = r1576 ^ r1638;
  wire _441 = _439 ^ _440;
  wire _442 = r1671 ^ r1702;
  wire _443 = r1750 ^ r1810;
  wire _444 = _442 ^ _443;
  wire _445 = _441 ^ _444;
  wire _446 = _438 ^ _445;
  wire _447 = _431 ^ _446;
  wire _448 = _416 | _447;
  wire _449 = r40 ^ r81;
  wire _450 = r127 ^ r211;
  wire _451 = _449 ^ _450;
  wire _452 = r229 ^ r297;
  wire _453 = r345 ^ r397;
  wire _454 = _452 ^ _453;
  wire _455 = _451 ^ _454;
  wire _456 = r464 ^ r560;
  wire _457 = r588 ^ r658;
  wire _458 = _456 ^ _457;
  wire _459 = r677 ^ r749;
  wire _460 = r786 ^ r841;
  wire _461 = _459 ^ _460;
  wire _462 = _458 ^ _461;
  wire _463 = _455 ^ _462;
  wire _464 = r916 ^ r978;
  wire _465 = r1012 ^ r1065;
  wire _466 = _464 ^ _465;
  wire _467 = r1126 ^ r1190;
  wire _468 = r1266 ^ r1375;
  wire _469 = _467 ^ _468;
  wire _470 = _466 ^ _469;
  wire _471 = r1431 ^ r1451;
  wire _472 = r1486 ^ r1531;
  wire _473 = _471 ^ _472;
  wire _474 = r1539 ^ r1637;
  wire _475 = r1778 ^ r1811;
  wire _476 = _474 ^ _475;
  wire _477 = _473 ^ _476;
  wire _478 = _470 ^ _477;
  wire _479 = _463 ^ _478;
  wire _480 = r39 ^ r80;
  wire _481 = r126 ^ r210;
  wire _482 = _480 ^ _481;
  wire _483 = r228 ^ r296;
  wire _484 = r344 ^ r396;
  wire _485 = _483 ^ _484;
  wire _486 = _482 ^ _485;
  wire _487 = r559 ^ r657;
  wire _488 = r785 ^ r840;
  wire _489 = _487 ^ _488;
  wire _490 = r915 ^ r977;
  wire _491 = r1011 ^ r1064;
  wire _492 = _490 ^ _491;
  wire _493 = _489 ^ _492;
  wire _494 = _486 ^ _493;
  wire _495 = r1125 ^ r1189;
  wire _496 = r1265 ^ r1374;
  wire _497 = _495 ^ _496;
  wire _498 = r1450 ^ r1483;
  wire _499 = r1530 ^ r1701;
  wire _500 = _498 ^ _499;
  wire _501 = _497 ^ _500;
  wire _502 = r1753 ^ r1809;
  wire _503 = r1842 ^ r1910;
  wire _504 = _502 ^ _503;
  wire _505 = r1925 ^ r1937;
  wire _506 = r1953 ^ r1961;
  wire _507 = _505 ^ _506;
  wire _508 = _504 ^ _507;
  wire _509 = _501 ^ _508;
  wire _510 = _494 ^ _509;
  wire _511 = _479 | _510;
  wire _512 = _448 | _511;
  wire _513 = _385 | _512;
  wire _514 = _258 | _513;
  wire _515 = r38 ^ r125;
  wire _516 = r209 ^ r227;
  wire _517 = _515 ^ _516;
  wire _518 = r295 ^ r343;
  wire _519 = r395 ^ r463;
  wire _520 = _518 ^ _519;
  wire _521 = _517 ^ _520;
  wire _522 = r587 ^ r656;
  wire _523 = r676 ^ r748;
  wire _524 = _522 ^ _523;
  wire _525 = r839 ^ r976;
  wire _526 = r1010 ^ r1063;
  wire _527 = _525 ^ _526;
  wire _528 = _524 ^ _527;
  wire _529 = _521 ^ _528;
  wire _530 = r1124 ^ r1188;
  wire _531 = r1264 ^ r1373;
  wire _532 = _530 ^ _531;
  wire _533 = r1430 ^ r1482;
  wire _534 = r1529 ^ r1538;
  wire _535 = _533 ^ _534;
  wire _536 = _532 ^ _535;
  wire _537 = r1636 ^ r1670;
  wire _538 = r1700 ^ r1900;
  wire _539 = _537 ^ _538;
  wire _540 = r2006 ^ r2023;
  wire _541 = r2034 ^ r2036;
  wire _542 = _540 ^ _541;
  wire _543 = _539 ^ _542;
  wire _544 = _536 ^ _543;
  wire _545 = _529 ^ _544;
  wire _546 = r37 ^ r79;
  wire _547 = r124 ^ r208;
  wire _548 = _546 ^ _547;
  wire _549 = r226 ^ r294;
  wire _550 = r342 ^ r394;
  wire _551 = _549 ^ _550;
  wire _552 = _548 ^ _551;
  wire _553 = r462 ^ r558;
  wire _554 = r586 ^ r655;
  wire _555 = _553 ^ _554;
  wire _556 = r675 ^ r747;
  wire _557 = r784 ^ r838;
  wire _558 = _556 ^ _557;
  wire _559 = _555 ^ _558;
  wire _560 = _552 ^ _559;
  wire _561 = r914 ^ r975;
  wire _562 = r1009 ^ r1062;
  wire _563 = _561 ^ _562;
  wire _564 = r1123 ^ r1187;
  wire _565 = r1263 ^ r1372;
  wire _566 = _564 ^ _565;
  wire _567 = _563 ^ _566;
  wire _568 = r1429 ^ r1449;
  wire _569 = r1481 ^ r1528;
  wire _570 = _568 ^ _569;
  wire _571 = r1699 ^ r1786;
  wire _572 = r1807 ^ r1812;
  wire _573 = _571 ^ _572;
  wire _574 = _570 ^ _573;
  wire _575 = _567 ^ _574;
  wire _576 = _560 ^ _575;
  wire _577 = _545 | _576;
  wire _578 = r36 ^ r78;
  wire _579 = r123 ^ r207;
  wire _580 = _578 ^ _579;
  wire _581 = r225 ^ r293;
  wire _582 = r341 ^ r393;
  wire _583 = _581 ^ _582;
  wire _584 = _580 ^ _583;
  wire _585 = r461 ^ r557;
  wire _586 = r585 ^ r654;
  wire _587 = _585 ^ _586;
  wire _588 = r674 ^ r746;
  wire _589 = r783 ^ r837;
  wire _590 = _588 ^ _589;
  wire _591 = _587 ^ _590;
  wire _592 = _584 ^ _591;
  wire _593 = r913 ^ r974;
  wire _594 = r1008 ^ r1061;
  wire _595 = _593 ^ _594;
  wire _596 = r1122 ^ r1186;
  wire _597 = r1262 ^ r1371;
  wire _598 = _596 ^ _597;
  wire _599 = _595 ^ _598;
  wire _600 = r1428 ^ r1448;
  wire _601 = r1480 ^ r1527;
  wire _602 = _600 ^ _601;
  wire _603 = r1537 ^ r1635;
  wire _604 = r1698 ^ r1730;
  wire _605 = _603 ^ _604;
  wire _606 = _602 ^ _605;
  wire _607 = _599 ^ _606;
  wire _608 = _592 ^ _607;
  wire _609 = r35 ^ r77;
  wire _610 = r122 ^ r278;
  wire _611 = _609 ^ _610;
  wire _612 = r340 ^ r460;
  wire _613 = r556 ^ r584;
  wire _614 = _612 ^ _613;
  wire _615 = _611 ^ _614;
  wire _616 = r745 ^ r782;
  wire _617 = r836 ^ r912;
  wire _618 = _616 ^ _617;
  wire _619 = r973 ^ r1261;
  wire _620 = r1370 ^ r1447;
  wire _621 = _619 ^ _620;
  wire _622 = _618 ^ _621;
  wire _623 = _615 ^ _622;
  wire _624 = r1479 ^ r1526;
  wire _625 = r1634 ^ r1669;
  wire _626 = _624 ^ _625;
  wire _627 = r1697 ^ r1772;
  wire _628 = r1849 ^ r1884;
  wire _629 = _627 ^ _628;
  wire _630 = _626 ^ _629;
  wire _631 = r1885 ^ r1957;
  wire _632 = r1964 ^ r1986;
  wire _633 = _631 ^ _632;
  wire _634 = r1989 ^ r2028;
  wire _635 = r2041 ^ r2042;
  wire _636 = _634 ^ _635;
  wire _637 = _633 ^ _636;
  wire _638 = _630 ^ _637;
  wire _639 = _623 ^ _638;
  wire _640 = _608 | _639;
  wire _641 = _577 | _640;
  wire _642 = r34 ^ r76;
  wire _643 = r277 ^ r292;
  wire _644 = _642 ^ _643;
  wire _645 = r339 ^ r459;
  wire _646 = r555 ^ r583;
  wire _647 = _645 ^ _646;
  wire _648 = _644 ^ _647;
  wire _649 = r673 ^ r781;
  wire _650 = r911 ^ r972;
  wire _651 = _649 ^ _650;
  wire _652 = r1007 ^ r1121;
  wire _653 = r1185 ^ r1260;
  wire _654 = _652 ^ _653;
  wire _655 = _651 ^ _654;
  wire _656 = _648 ^ _655;
  wire _657 = r1328 ^ r1427;
  wire _658 = r1446 ^ r1478;
  wire _659 = _657 ^ _658;
  wire _660 = r1508 ^ r1633;
  wire _661 = r1696 ^ r1770;
  wire _662 = _660 ^ _661;
  wire _663 = _659 ^ _662;
  wire _664 = r1773 ^ r1787;
  wire _665 = r1844 ^ r1852;
  wire _666 = _664 ^ _665;
  wire _667 = r1854 ^ r1857;
  wire _668 = r1858 ^ r1876;
  wire _669 = _667 ^ _668;
  wire _670 = _666 ^ _669;
  wire _671 = _663 ^ _670;
  wire _672 = _656 ^ _671;
  wire _673 = r33 ^ r75;
  wire _674 = r121 ^ r206;
  wire _675 = _673 ^ _674;
  wire _676 = r276 ^ r291;
  wire _677 = r338 ^ r392;
  wire _678 = _676 ^ _677;
  wire _679 = _675 ^ _678;
  wire _680 = r458 ^ r554;
  wire _681 = r653 ^ r672;
  wire _682 = _680 ^ _681;
  wire _683 = r744 ^ r780;
  wire _684 = r835 ^ r910;
  wire _685 = _683 ^ _684;
  wire _686 = _682 ^ _685;
  wire _687 = _679 ^ _686;
  wire _688 = r971 ^ r1006;
  wire _689 = r1111 ^ r1120;
  wire _690 = _688 ^ _689;
  wire _691 = r1184 ^ r1259;
  wire _692 = r1327 ^ r1369;
  wire _693 = _691 ^ _692;
  wire _694 = _690 ^ _693;
  wire _695 = r1425 ^ r1426;
  wire _696 = r1445 ^ r1477;
  wire _697 = _695 ^ _696;
  wire _698 = r1632 ^ r1668;
  wire _699 = r1932 ^ r1934;
  wire _700 = _698 ^ _699;
  wire _701 = _697 ^ _700;
  wire _702 = _694 ^ _701;
  wire _703 = _687 ^ _702;
  wire _704 = _672 | _703;
  wire _705 = r32 ^ r74;
  wire _706 = r120 ^ r205;
  wire _707 = _705 ^ _706;
  wire _708 = r275 ^ r290;
  wire _709 = r337 ^ r446;
  wire _710 = _708 ^ _709;
  wire _711 = _707 ^ _710;
  wire _712 = r457 ^ r582;
  wire _713 = r671 ^ r743;
  wire _714 = _712 ^ _713;
  wire _715 = r834 ^ r970;
  wire _716 = r1119 ^ r1183;
  wire _717 = _715 ^ _716;
  wire _718 = _714 ^ _717;
  wire _719 = _711 ^ _718;
  wire _720 = r1258 ^ r1326;
  wire _721 = r1368 ^ r1390;
  wire _722 = _720 ^ _721;
  wire _723 = r1424 ^ r1507;
  wire _724 = r1631 ^ r1765;
  wire _725 = _723 ^ _724;
  wire _726 = _722 ^ _725;
  wire _727 = r1793 ^ r1795;
  wire _728 = r1882 ^ r1903;
  wire _729 = _727 ^ _728;
  wire _730 = r1941 ^ r1987;
  wire _731 = r2032 ^ r2035;
  wire _732 = _730 ^ _731;
  wire _733 = _729 ^ _732;
  wire _734 = _726 ^ _733;
  wire _735 = _719 ^ _734;
  wire _736 = r31 ^ r73;
  wire _737 = r119 ^ r204;
  wire _738 = _736 ^ _737;
  wire _739 = r274 ^ r289;
  wire _740 = r336 ^ r445;
  wire _741 = _739 ^ _740;
  wire _742 = _738 ^ _741;
  wire _743 = r456 ^ r553;
  wire _744 = r581 ^ r652;
  wire _745 = _743 ^ _744;
  wire _746 = r742 ^ r779;
  wire _747 = r833 ^ r909;
  wire _748 = _746 ^ _747;
  wire _749 = _745 ^ _748;
  wire _750 = _742 ^ _749;
  wire _751 = r969 ^ r1005;
  wire _752 = r1109 ^ r1118;
  wire _753 = _751 ^ _752;
  wire _754 = r1182 ^ r1257;
  wire _755 = r1325 ^ r1367;
  wire _756 = _754 ^ _755;
  wire _757 = _753 ^ _756;
  wire _758 = r1389 ^ r1423;
  wire _759 = r1444 ^ r1476;
  wire _760 = _758 ^ _759;
  wire _761 = r1630 ^ r1754;
  wire _762 = r1802 ^ r1813;
  wire _763 = _761 ^ _762;
  wire _764 = _760 ^ _763;
  wire _765 = _757 ^ _764;
  wire _766 = _750 ^ _765;
  wire _767 = _735 | _766;
  wire _768 = _704 | _767;
  wire _769 = _641 | _768;
  wire _770 = r30 ^ r72;
  wire _771 = r118 ^ r203;
  wire _772 = _770 ^ _771;
  wire _773 = r273 ^ r288;
  wire _774 = r335 ^ r444;
  wire _775 = _773 ^ _774;
  wire _776 = _772 ^ _775;
  wire _777 = r455 ^ r552;
  wire _778 = r580 ^ r651;
  wire _779 = _777 ^ _778;
  wire _780 = r670 ^ r741;
  wire _781 = r778 ^ r832;
  wire _782 = _780 ^ _781;
  wire _783 = _779 ^ _782;
  wire _784 = _776 ^ _783;
  wire _785 = r908 ^ r968;
  wire _786 = r1004 ^ r1117;
  wire _787 = _785 ^ _786;
  wire _788 = r1181 ^ r1324;
  wire _789 = r1366 ^ r1388;
  wire _790 = _788 ^ _789;
  wire _791 = _787 ^ _790;
  wire _792 = r1422 ^ r1443;
  wire _793 = r1506 ^ r1667;
  wire _794 = _792 ^ _793;
  wire _795 = r1695 ^ r1760;
  wire _796 = r1784 ^ r1814;
  wire _797 = _795 ^ _796;
  wire _798 = _794 ^ _797;
  wire _799 = _791 ^ _798;
  wire _800 = _784 ^ _799;
  wire _801 = r29 ^ r71;
  wire _802 = r117 ^ r202;
  wire _803 = _801 ^ _802;
  wire _804 = r287 ^ r443;
  wire _805 = r454 ^ r551;
  wire _806 = _804 ^ _805;
  wire _807 = _803 ^ _806;
  wire _808 = r579 ^ r650;
  wire _809 = r669 ^ r740;
  wire _810 = _808 ^ _809;
  wire _811 = r831 ^ r907;
  wire _812 = r967 ^ r1107;
  wire _813 = _811 ^ _812;
  wire _814 = _810 ^ _813;
  wire _815 = _807 ^ _814;
  wire _816 = r1116 ^ r1180;
  wire _817 = r1256 ^ r1323;
  wire _818 = _816 ^ _817;
  wire _819 = r1365 ^ r1387;
  wire _820 = r1466 ^ r1504;
  wire _821 = _819 ^ _820;
  wire _822 = _818 ^ _821;
  wire _823 = r1629 ^ r1759;
  wire _824 = r1766 ^ r1800;
  wire _825 = _823 ^ _824;
  wire _826 = r1841 ^ r1862;
  wire _827 = r1875 ^ r1877;
  wire _828 = _826 ^ _827;
  wire _829 = _825 ^ _828;
  wire _830 = _822 ^ _829;
  wire _831 = _815 ^ _830;
  wire _832 = _800 | _831;
  wire _833 = r28 ^ r70;
  wire _834 = r116 ^ r201;
  wire _835 = _833 ^ _834;
  wire _836 = r272 ^ r286;
  wire _837 = r334 ^ r442;
  wire _838 = _836 ^ _837;
  wire _839 = _835 ^ _838;
  wire _840 = r453 ^ r550;
  wire _841 = r578 ^ r649;
  wire _842 = _840 ^ _841;
  wire _843 = r721 ^ r739;
  wire _844 = r829 ^ r886;
  wire _845 = _843 ^ _844;
  wire _846 = _842 ^ _845;
  wire _847 = _839 ^ _846;
  wire _848 = r906 ^ r966;
  wire _849 = r1058 ^ r1106;
  wire _850 = _848 ^ _849;
  wire _851 = r1115 ^ r1179;
  wire _852 = r1255 ^ r1322;
  wire _853 = _851 ^ _852;
  wire _854 = _850 ^ _853;
  wire _855 = r1364 ^ r1386;
  wire _856 = r1421 ^ r1465;
  wire _857 = _855 ^ _856;
  wire _858 = r1558 ^ r1666;
  wire _859 = r1694 ^ r1731;
  wire _860 = _858 ^ _859;
  wire _861 = _857 ^ _860;
  wire _862 = _854 ^ _861;
  wire _863 = _847 ^ _862;
  wire _864 = r27 ^ r69;
  wire _865 = r115 ^ r200;
  wire _866 = _864 ^ _865;
  wire _867 = r285 ^ r441;
  wire _868 = r452 ^ r549;
  wire _869 = _867 ^ _868;
  wire _870 = _866 ^ _869;
  wire _871 = r648 ^ r720;
  wire _872 = r738 ^ r828;
  wire _873 = _871 ^ _872;
  wire _874 = r885 ^ r905;
  wire _875 = r965 ^ r1057;
  wire _876 = _874 ^ _875;
  wire _877 = _873 ^ _876;
  wire _878 = _870 ^ _877;
  wire _879 = r1105 ^ r1178;
  wire _880 = r1321 ^ r1385;
  wire _881 = _879 ^ _880;
  wire _882 = r1420 ^ r1464;
  wire _883 = r1557 ^ r1665;
  wire _884 = _882 ^ _883;
  wire _885 = _881 ^ _884;
  wire _886 = r1769 ^ r1780;
  wire _887 = r1828 ^ r1839;
  wire _888 = _886 ^ _887;
  wire _889 = r1848 ^ r1869;
  wire _890 = r1933 ^ r1935;
  wire _891 = _889 ^ _890;
  wire _892 = _888 ^ _891;
  wire _893 = _885 ^ _892;
  wire _894 = _878 ^ _893;
  wire _895 = _863 | _894;
  wire _896 = _832 | _895;
  wire _897 = r26 ^ r68;
  wire _898 = r114 ^ r199;
  wire _899 = _897 ^ _898;
  wire _900 = r271 ^ r333;
  wire _901 = r440 ^ r451;
  wire _902 = _900 ^ _901;
  wire _903 = _899 ^ _902;
  wire _904 = r548 ^ r577;
  wire _905 = r647 ^ r719;
  wire _906 = _904 ^ _905;
  wire _907 = r737 ^ r827;
  wire _908 = r884 ^ r904;
  wire _909 = _907 ^ _908;
  wire _910 = _906 ^ _909;
  wire _911 = _903 ^ _910;
  wire _912 = r964 ^ r1056;
  wire _913 = r1104 ^ r1114;
  wire _914 = _912 ^ _913;
  wire _915 = r1177 ^ r1254;
  wire _916 = r1320 ^ r1363;
  wire _917 = _915 ^ _916;
  wire _918 = _914 ^ _917;
  wire _919 = r1384 ^ r1419;
  wire _920 = r1463 ^ r1556;
  wire _921 = _919 ^ _920;
  wire _922 = r1628 ^ r1664;
  wire _923 = r1693 ^ r1732;
  wire _924 = _922 ^ _923;
  wire _925 = _921 ^ _924;
  wire _926 = _918 ^ _925;
  wire _927 = _911 ^ _926;
  wire _928 = r25 ^ r67;
  wire _929 = r113 ^ r270;
  wire _930 = _928 ^ _929;
  wire _931 = r450 ^ r547;
  wire _932 = r576 ^ r646;
  wire _933 = _931 ^ _932;
  wire _934 = _930 ^ _933;
  wire _935 = r883 ^ r903;
  wire _936 = r1055 ^ r1103;
  wire _937 = _935 ^ _936;
  wire _938 = r1253 ^ r1319;
  wire _939 = r1362 ^ r1418;
  wire _940 = _938 ^ _939;
  wire _941 = _937 ^ _940;
  wire _942 = _934 ^ _941;
  wire _943 = r1462 ^ r1555;
  wire _944 = r1627 ^ r1758;
  wire _945 = _943 ^ _944;
  wire _946 = r1781 ^ r1803;
  wire _947 = r1894 ^ r1898;
  wire _948 = _946 ^ _947;
  wire _949 = _945 ^ _948;
  wire _950 = r1913 ^ r1922;
  wire _951 = r1955 ^ r1960;
  wire _952 = _950 ^ _951;
  wire _953 = r1980 ^ r1985;
  wire _954 = r1988 ^ r1990;
  wire _955 = _953 ^ _954;
  wire _956 = _952 ^ _955;
  wire _957 = _949 ^ _956;
  wire _958 = _942 ^ _957;
  wire _959 = _927 | _958;
  wire _960 = r24 ^ r66;
  wire _961 = r112 ^ r198;
  wire _962 = _960 ^ _961;
  wire _963 = r269 ^ r284;
  wire _964 = r390 ^ r439;
  wire _965 = _963 ^ _964;
  wire _966 = _962 ^ _965;
  wire _967 = r449 ^ r546;
  wire _968 = r575 ^ r645;
  wire _969 = _967 ^ _968;
  wire _970 = r718 ^ r736;
  wire _971 = r882 ^ r902;
  wire _972 = _970 ^ _971;
  wire _973 = _969 ^ _972;
  wire _974 = _966 ^ _973;
  wire _975 = r963 ^ r1054;
  wire _976 = r1102 ^ r1176;
  wire _977 = _975 ^ _976;
  wire _978 = r1252 ^ r1318;
  wire _979 = r1334 ^ r1361;
  wire _980 = _978 ^ _979;
  wire _981 = _977 ^ _980;
  wire _982 = r1417 ^ r1461;
  wire _983 = r1513 ^ r1663;
  wire _984 = _982 ^ _983;
  wire _985 = r1692 ^ r1771;
  wire _986 = r1806 ^ r1815;
  wire _987 = _985 ^ _986;
  wire _988 = _984 ^ _987;
  wire _989 = _981 ^ _988;
  wire _990 = _974 ^ _989;
  wire _991 = r23 ^ r65;
  wire _992 = r197 ^ r283;
  wire _993 = _991 ^ _992;
  wire _994 = r389 ^ r438;
  wire _995 = r448 ^ r545;
  wire _996 = _994 ^ _995;
  wire _997 = _993 ^ _996;
  wire _998 = r574 ^ r644;
  wire _999 = r717 ^ r735;
  wire _1000 = _998 ^ _999;
  wire _1001 = r826 ^ r881;
  wire _1002 = r901 ^ r962;
  wire _1003 = _1001 ^ _1002;
  wire _1004 = _1000 ^ _1003;
  wire _1005 = _997 ^ _1004;
  wire _1006 = r1053 ^ r1101;
  wire _1007 = r1175 ^ r1251;
  wire _1008 = _1006 ^ _1007;
  wire _1009 = r1317 ^ r1333;
  wire _1010 = r1360 ^ r1416;
  wire _1011 = _1009 ^ _1010;
  wire _1012 = _1008 ^ _1011;
  wire _1013 = r1460 ^ r1554;
  wire _1014 = r1626 ^ r1782;
  wire _1015 = _1013 ^ _1014;
  wire _1016 = r1790 ^ r1921;
  wire _1017 = r1952 ^ r1962;
  wire _1018 = _1016 ^ _1017;
  wire _1019 = _1015 ^ _1018;
  wire _1020 = _1012 ^ _1019;
  wire _1021 = _1005 ^ _1020;
  wire _1022 = _990 | _1021;
  wire _1023 = _959 | _1022;
  wire _1024 = _896 | _1023;
  wire _1025 = _769 | _1024;
  wire _1026 = _514 | _1025;
  wire _1027 = r22 ^ r64;
  wire _1028 = r111 ^ r268;
  wire _1029 = _1027 ^ _1028;
  wire _1030 = r388 ^ r504;
  wire _1031 = r544 ^ r573;
  wire _1032 = _1030 ^ _1031;
  wire _1033 = _1029 ^ _1032;
  wire _1034 = r643 ^ r734;
  wire _1035 = r825 ^ r880;
  wire _1036 = _1034 ^ _1035;
  wire _1037 = r900 ^ r961;
  wire _1038 = r1052 ^ r1250;
  wire _1039 = _1037 ^ _1038;
  wire _1040 = _1036 ^ _1039;
  wire _1041 = _1033 ^ _1040;
  wire _1042 = r1316 ^ r1359;
  wire _1043 = r1459 ^ r1662;
  wire _1044 = _1042 ^ _1043;
  wire _1045 = r1691 ^ r1742;
  wire _1046 = r1826 ^ r1831;
  wire _1047 = _1045 ^ _1046;
  wire _1048 = _1044 ^ _1047;
  wire _1049 = r1943 ^ r1958;
  wire _1050 = r1959 ^ r1973;
  wire _1051 = _1049 ^ _1050;
  wire _1052 = r1999 ^ r2008;
  wire _1053 = r2027 ^ r2029;
  wire _1054 = _1052 ^ _1053;
  wire _1055 = _1051 ^ _1054;
  wire _1056 = _1048 ^ _1055;
  wire _1057 = _1041 ^ _1056;
  wire _1058 = r21 ^ r63;
  wire _1059 = r169 ^ r196;
  wire _1060 = _1058 ^ _1059;
  wire _1061 = r267 ^ r282;
  wire _1062 = r387 ^ r437;
  wire _1063 = _1061 ^ _1062;
  wire _1064 = _1060 ^ _1063;
  wire _1065 = r503 ^ r543;
  wire _1066 = r572 ^ r642;
  wire _1067 = _1065 ^ _1066;
  wire _1068 = r716 ^ r733;
  wire _1069 = r824 ^ r879;
  wire _1070 = _1068 ^ _1069;
  wire _1071 = _1067 ^ _1070;
  wire _1072 = _1064 ^ _1071;
  wire _1073 = r899 ^ r960;
  wire _1074 = r1051 ^ r1100;
  wire _1075 = _1073 ^ _1074;
  wire _1076 = r1174 ^ r1249;
  wire _1077 = r1315 ^ r1332;
  wire _1078 = _1076 ^ _1077;
  wire _1079 = _1075 ^ _1078;
  wire _1080 = r1358 ^ r1415;
  wire _1081 = r1458 ^ r1512;
  wire _1082 = _1080 ^ _1081;
  wire _1083 = r1574 ^ r1625;
  wire _1084 = r1690 ^ r1733;
  wire _1085 = _1083 ^ _1084;
  wire _1086 = _1082 ^ _1085;
  wire _1087 = _1079 ^ _1086;
  wire _1088 = _1072 ^ _1087;
  wire _1089 = _1057 | _1088;
  wire _1090 = r20 ^ r62;
  wire _1091 = r168 ^ r195;
  wire _1092 = _1090 ^ _1091;
  wire _1093 = r266 ^ r281;
  wire _1094 = r386 ^ r436;
  wire _1095 = _1093 ^ _1094;
  wire _1096 = _1092 ^ _1095;
  wire _1097 = r502 ^ r542;
  wire _1098 = r571 ^ r641;
  wire _1099 = _1097 ^ _1098;
  wire _1100 = r715 ^ r732;
  wire _1101 = r823 ^ r878;
  wire _1102 = _1100 ^ _1101;
  wire _1103 = _1099 ^ _1102;
  wire _1104 = _1096 ^ _1103;
  wire _1105 = r898 ^ r959;
  wire _1106 = r1050 ^ r1099;
  wire _1107 = _1105 ^ _1106;
  wire _1108 = r1173 ^ r1248;
  wire _1109 = r1314 ^ r1331;
  wire _1110 = _1108 ^ _1109;
  wire _1111 = _1107 ^ _1110;
  wire _1112 = r1414 ^ r1511;
  wire _1113 = r1573 ^ r1606;
  wire _1114 = _1112 ^ _1113;
  wire _1115 = r1624 ^ r1661;
  wire _1116 = r1822 ^ r1878;
  wire _1117 = _1115 ^ _1116;
  wire _1118 = _1114 ^ _1117;
  wire _1119 = _1111 ^ _1118;
  wire _1120 = _1104 ^ _1119;
  wire _1121 = r19 ^ r61;
  wire _1122 = r167 ^ r194;
  wire _1123 = _1121 ^ _1122;
  wire _1124 = r265 ^ r280;
  wire _1125 = r385 ^ r435;
  wire _1126 = _1124 ^ _1125;
  wire _1127 = _1123 ^ _1126;
  wire _1128 = r501 ^ r541;
  wire _1129 = r570 ^ r640;
  wire _1130 = _1128 ^ _1129;
  wire _1131 = r714 ^ r731;
  wire _1132 = r822 ^ r877;
  wire _1133 = _1131 ^ _1132;
  wire _1134 = _1130 ^ _1133;
  wire _1135 = _1127 ^ _1134;
  wire _1136 = r897 ^ r958;
  wire _1137 = r1049 ^ r1098;
  wire _1138 = _1136 ^ _1137;
  wire _1139 = r1172 ^ r1247;
  wire _1140 = r1313 ^ r1330;
  wire _1141 = _1139 ^ _1140;
  wire _1142 = _1138 ^ _1141;
  wire _1143 = r1357 ^ r1413;
  wire _1144 = r1510 ^ r1605;
  wire _1145 = _1143 ^ _1144;
  wire _1146 = r1623 ^ r1660;
  wire _1147 = r1689 ^ r1734;
  wire _1148 = _1146 ^ _1147;
  wire _1149 = _1145 ^ _1148;
  wire _1150 = _1142 ^ _1149;
  wire _1151 = _1135 ^ _1150;
  wire _1152 = _1120 | _1151;
  wire _1153 = _1089 | _1152;
  wire _1154 = r18 ^ r60;
  wire _1155 = r166 ^ r264;
  wire _1156 = _1154 ^ _1155;
  wire _1157 = r384 ^ r434;
  wire _1158 = r500 ^ r540;
  wire _1159 = _1157 ^ _1158;
  wire _1160 = _1156 ^ _1159;
  wire _1161 = r639 ^ r821;
  wire _1162 = r896 ^ r957;
  wire _1163 = _1161 ^ _1162;
  wire _1164 = r1048 ^ r1171;
  wire _1165 = r1246 ^ r1329;
  wire _1166 = _1164 ^ _1165;
  wire _1167 = _1163 ^ _1166;
  wire _1168 = _1160 ^ _1167;
  wire _1169 = r1356 ^ r1412;
  wire _1170 = r1604 ^ r1622;
  wire _1171 = _1169 ^ _1170;
  wire _1172 = r1659 ^ r1743;
  wire _1173 = r1873 ^ r1888;
  wire _1174 = _1172 ^ _1173;
  wire _1175 = _1171 ^ _1174;
  wire _1176 = r1947 ^ r1950;
  wire _1177 = r1969 ^ r1976;
  wire _1178 = _1176 ^ _1177;
  wire _1179 = r1995 ^ r2002;
  wire _1180 = r2022 ^ r2030;
  wire _1181 = _1179 ^ _1180;
  wire _1182 = _1178 ^ _1181;
  wire _1183 = _1175 ^ _1182;
  wire _1184 = _1168 ^ _1183;
  wire _1185 = r17 ^ r59;
  wire _1186 = r165 ^ r193;
  wire _1187 = _1185 ^ _1186;
  wire _1188 = r263 ^ r331;
  wire _1189 = r383 ^ r433;
  wire _1190 = _1188 ^ _1189;
  wire _1191 = _1187 ^ _1190;
  wire _1192 = r499 ^ r539;
  wire _1193 = r569 ^ r638;
  wire _1194 = _1192 ^ _1193;
  wire _1195 = r713 ^ r730;
  wire _1196 = r820 ^ r876;
  wire _1197 = _1195 ^ _1196;
  wire _1198 = _1194 ^ _1197;
  wire _1199 = _1191 ^ _1198;
  wire _1200 = r895 ^ r956;
  wire _1201 = r1047 ^ r1097;
  wire _1202 = _1200 ^ _1201;
  wire _1203 = r1163 ^ r1170;
  wire _1204 = r1245 ^ r1282;
  wire _1205 = _1203 ^ _1204;
  wire _1206 = _1202 ^ _1205;
  wire _1207 = r1312 ^ r1355;
  wire _1208 = r1572 ^ r1603;
  wire _1209 = _1207 ^ _1208;
  wire _1210 = r1621 ^ r1658;
  wire _1211 = r1688 ^ r1735;
  wire _1212 = _1210 ^ _1211;
  wire _1213 = _1209 ^ _1212;
  wire _1214 = _1206 ^ _1213;
  wire _1215 = _1199 ^ _1214;
  wire _1216 = _1184 | _1215;
  wire _1217 = r16 ^ r58;
  wire _1218 = r164 ^ r192;
  wire _1219 = _1217 ^ _1218;
  wire _1220 = r262 ^ r330;
  wire _1221 = r382 ^ r432;
  wire _1222 = _1220 ^ _1221;
  wire _1223 = _1219 ^ _1222;
  wire _1224 = r498 ^ r538;
  wire _1225 = r568 ^ r637;
  wire _1226 = _1224 ^ _1225;
  wire _1227 = r712 ^ r729;
  wire _1228 = r875 ^ r894;
  wire _1229 = _1227 ^ _1228;
  wire _1230 = _1226 ^ _1229;
  wire _1231 = _1223 ^ _1230;
  wire _1232 = r955 ^ r1046;
  wire _1233 = r1096 ^ r1162;
  wire _1234 = _1232 ^ _1233;
  wire _1235 = r1244 ^ r1281;
  wire _1236 = r1311 ^ r1411;
  wire _1237 = _1235 ^ _1236;
  wire _1238 = _1234 ^ _1237;
  wire _1239 = r1518 ^ r1571;
  wire _1240 = r1620 ^ r1767;
  wire _1241 = _1239 ^ _1240;
  wire _1242 = r1881 ^ r1897;
  wire _1243 = r1909 ^ r1915;
  wire _1244 = _1242 ^ _1243;
  wire _1245 = _1241 ^ _1244;
  wire _1246 = _1238 ^ _1245;
  wire _1247 = _1231 ^ _1246;
  wire _1248 = r15 ^ r57;
  wire _1249 = r163 ^ r191;
  wire _1250 = _1248 ^ _1249;
  wire _1251 = r261 ^ r329;
  wire _1252 = r381 ^ r431;
  wire _1253 = _1251 ^ _1252;
  wire _1254 = _1250 ^ _1253;
  wire _1255 = r497 ^ r537;
  wire _1256 = r567 ^ r636;
  wire _1257 = _1255 ^ _1256;
  wire _1258 = r711 ^ r728;
  wire _1259 = r819 ^ r874;
  wire _1260 = _1258 ^ _1259;
  wire _1261 = _1257 ^ _1260;
  wire _1262 = _1254 ^ _1261;
  wire _1263 = r893 ^ r954;
  wire _1264 = r1045 ^ r1095;
  wire _1265 = _1263 ^ _1264;
  wire _1266 = r1161 ^ r1243;
  wire _1267 = r1280 ^ r1310;
  wire _1268 = _1266 ^ _1267;
  wire _1269 = _1265 ^ _1268;
  wire _1270 = r1354 ^ r1410;
  wire _1271 = r1517 ^ r1570;
  wire _1272 = _1270 ^ _1271;
  wire _1273 = r1602 ^ r1619;
  wire _1274 = r1657 ^ r1736;
  wire _1275 = _1273 ^ _1274;
  wire _1276 = _1272 ^ _1275;
  wire _1277 = _1269 ^ _1276;
  wire _1278 = _1262 ^ _1277;
  wire _1279 = _1247 | _1278;
  wire _1280 = _1216 | _1279;
  wire _1281 = _1153 | _1280;
  wire _1282 = r14 ^ r56;
  wire _1283 = r162 ^ r260;
  wire _1284 = _1282 ^ _1283;
  wire _1285 = r380 ^ r430;
  wire _1286 = r496 ^ r536;
  wire _1287 = _1285 ^ _1286;
  wire _1288 = _1284 ^ _1287;
  wire _1289 = r566 ^ r635;
  wire _1290 = r727 ^ r818;
  wire _1291 = _1289 ^ _1290;
  wire _1292 = r873 ^ r892;
  wire _1293 = r953 ^ r1044;
  wire _1294 = _1292 ^ _1293;
  wire _1295 = _1291 ^ _1294;
  wire _1296 = _1288 ^ _1295;
  wire _1297 = r1160 ^ r1242;
  wire _1298 = r1279 ^ r1353;
  wire _1299 = _1297 ^ _1298;
  wire _1300 = r1409 ^ r1569;
  wire _1301 = r1601 ^ r1618;
  wire _1302 = _1300 ^ _1301;
  wire _1303 = _1299 ^ _1302;
  wire _1304 = r1656 ^ r1717;
  wire _1305 = r1856 ^ r1912;
  wire _1306 = _1304 ^ _1305;
  wire _1307 = r1974 ^ r1984;
  wire _1308 = r1991 ^ r1992;
  wire _1309 = _1307 ^ _1308;
  wire _1310 = _1306 ^ _1309;
  wire _1311 = _1303 ^ _1310;
  wire _1312 = _1296 ^ _1311;
  wire _1313 = r13 ^ r55;
  wire _1314 = r161 ^ r190;
  wire _1315 = _1313 ^ _1314;
  wire _1316 = r259 ^ r328;
  wire _1317 = r379 ^ r429;
  wire _1318 = _1316 ^ _1317;
  wire _1319 = _1315 ^ _1318;
  wire _1320 = r495 ^ r535;
  wire _1321 = r565 ^ r634;
  wire _1322 = _1320 ^ _1321;
  wire _1323 = r710 ^ r726;
  wire _1324 = r817 ^ r872;
  wire _1325 = _1323 ^ _1324;
  wire _1326 = _1322 ^ _1325;
  wire _1327 = _1319 ^ _1326;
  wire _1328 = r891 ^ r952;
  wire _1329 = r1043 ^ r1094;
  wire _1330 = _1328 ^ _1329;
  wire _1331 = r1159 ^ r1278;
  wire _1332 = r1309 ^ r1352;
  wire _1333 = _1331 ^ _1332;
  wire _1334 = _1330 ^ _1333;
  wire _1335 = r1408 ^ r1568;
  wire _1336 = r1600 ^ r1617;
  wire _1337 = _1335 ^ _1336;
  wire _1338 = r1716 ^ r1748;
  wire _1339 = r1755 ^ r1816;
  wire _1340 = _1338 ^ _1339;
  wire _1341 = _1337 ^ _1340;
  wire _1342 = _1334 ^ _1341;
  wire _1343 = _1327 ^ _1342;
  wire _1344 = _1312 | _1343;
  wire _1345 = r12 ^ r54;
  wire _1346 = r160 ^ r189;
  wire _1347 = _1345 ^ _1346;
  wire _1348 = r258 ^ r327;
  wire _1349 = r378 ^ r428;
  wire _1350 = _1348 ^ _1349;
  wire _1351 = _1347 ^ _1350;
  wire _1352 = r494 ^ r534;
  wire _1353 = r564 ^ r633;
  wire _1354 = _1352 ^ _1353;
  wire _1355 = r709 ^ r725;
  wire _1356 = r816 ^ r871;
  wire _1357 = _1355 ^ _1356;
  wire _1358 = _1354 ^ _1357;
  wire _1359 = _1351 ^ _1358;
  wire _1360 = r890 ^ r951;
  wire _1361 = r1042 ^ r1093;
  wire _1362 = _1360 ^ _1361;
  wire _1363 = r1158 ^ r1241;
  wire _1364 = r1308 ^ r1351;
  wire _1365 = _1363 ^ _1364;
  wire _1366 = _1362 ^ _1365;
  wire _1367 = r1407 ^ r1516;
  wire _1368 = r1553 ^ r1567;
  wire _1369 = _1367 ^ _1368;
  wire _1370 = r1616 ^ r1655;
  wire _1371 = r1715 ^ r1737;
  wire _1372 = _1370 ^ _1371;
  wire _1373 = _1369 ^ _1372;
  wire _1374 = _1366 ^ _1373;
  wire _1375 = _1359 ^ _1374;
  wire _1376 = r109 ^ r159;
  wire _1377 = r188 ^ r257;
  wire _1378 = _1376 ^ _1377;
  wire _1379 = r326 ^ r377;
  wire _1380 = r427 ^ r493;
  wire _1381 = _1379 ^ _1380;
  wire _1382 = _1378 ^ _1381;
  wire _1383 = r533 ^ r563;
  wire _1384 = r632 ^ r708;
  wire _1385 = _1383 ^ _1384;
  wire _1386 = r815 ^ r870;
  wire _1387 = r889 ^ r950;
  wire _1388 = _1386 ^ _1387;
  wire _1389 = _1385 ^ _1388;
  wire _1390 = _1382 ^ _1389;
  wire _1391 = r1041 ^ r1092;
  wire _1392 = r1157 ^ r1277;
  wire _1393 = _1391 ^ _1392;
  wire _1394 = r1307 ^ r1350;
  wire _1395 = r1406 ^ r1515;
  wire _1396 = _1394 ^ _1395;
  wire _1397 = _1393 ^ _1396;
  wire _1398 = r1566 ^ r1599;
  wire _1399 = r1615 ^ r1654;
  wire _1400 = _1398 ^ _1399;
  wire _1401 = r1749 ^ r1762;
  wire _1402 = r1889 ^ r1906;
  wire _1403 = _1401 ^ _1402;
  wire _1404 = _1400 ^ _1403;
  wire _1405 = _1397 ^ _1404;
  wire _1406 = _1390 ^ _1405;
  wire _1407 = _1375 | _1406;
  wire _1408 = _1344 | _1407;
  wire _1409 = r11 ^ r108;
  wire _1410 = r158 ^ r187;
  wire _1411 = _1409 ^ _1410;
  wire _1412 = r256 ^ r325;
  wire _1413 = r376 ^ r426;
  wire _1414 = _1412 ^ _1413;
  wire _1415 = _1411 ^ _1414;
  wire _1416 = r492 ^ r532;
  wire _1417 = r562 ^ r631;
  wire _1418 = _1416 ^ _1417;
  wire _1419 = r707 ^ r724;
  wire _1420 = r814 ^ r869;
  wire _1421 = _1419 ^ _1420;
  wire _1422 = _1418 ^ _1421;
  wire _1423 = _1415 ^ _1422;
  wire _1424 = r888 ^ r949;
  wire _1425 = r1040 ^ r1091;
  wire _1426 = _1424 ^ _1425;
  wire _1427 = r1156 ^ r1217;
  wire _1428 = r1240 ^ r1276;
  wire _1429 = _1427 ^ _1428;
  wire _1430 = _1426 ^ _1429;
  wire _1431 = r1306 ^ r1349;
  wire _1432 = r1405 ^ r1565;
  wire _1433 = _1431 ^ _1432;
  wire _1434 = r1598 ^ r1614;
  wire _1435 = r1714 ^ r1738;
  wire _1436 = _1434 ^ _1435;
  wire _1437 = _1433 ^ _1436;
  wire _1438 = _1430 ^ _1437;
  wire _1439 = _1423 ^ _1438;
  wire _1440 = r10 ^ r107;
  wire _1441 = r157 ^ r186;
  wire _1442 = _1440 ^ _1441;
  wire _1443 = r255 ^ r324;
  wire _1444 = r375 ^ r425;
  wire _1445 = _1443 ^ _1444;
  wire _1446 = _1442 ^ _1445;
  wire _1447 = r491 ^ r531;
  wire _1448 = r561 ^ r630;
  wire _1449 = _1447 ^ _1448;
  wire _1450 = r706 ^ r723;
  wire _1451 = r813 ^ r868;
  wire _1452 = _1450 ^ _1451;
  wire _1453 = _1449 ^ _1452;
  wire _1454 = _1446 ^ _1453;
  wire _1455 = r943 ^ r948;
  wire _1456 = r1039 ^ r1090;
  wire _1457 = _1455 ^ _1456;
  wire _1458 = r1155 ^ r1216;
  wire _1459 = r1224 ^ r1305;
  wire _1460 = _1458 ^ _1459;
  wire _1461 = _1457 ^ _1460;
  wire _1462 = r1348 ^ r1404;
  wire _1463 = r1564 ^ r1597;
  wire _1464 = _1462 ^ _1463;
  wire _1465 = r1653 ^ r1713;
  wire _1466 = r1756 ^ r1817;
  wire _1467 = _1465 ^ _1466;
  wire _1468 = _1464 ^ _1467;
  wire _1469 = _1461 ^ _1468;
  wire _1470 = _1454 ^ _1469;
  wire _1471 = _1439 | _1470;
  wire _1472 = r9 ^ r106;
  wire _1473 = r156 ^ r185;
  wire _1474 = _1472 ^ _1473;
  wire _1475 = r254 ^ r323;
  wire _1476 = r374 ^ r424;
  wire _1477 = _1475 ^ _1476;
  wire _1478 = _1474 ^ _1477;
  wire _1479 = r490 ^ r530;
  wire _1480 = r615 ^ r705;
  wire _1481 = _1479 ^ _1480;
  wire _1482 = r776 ^ r812;
  wire _1483 = r867 ^ r947;
  wire _1484 = _1482 ^ _1483;
  wire _1485 = _1481 ^ _1484;
  wire _1486 = _1478 ^ _1485;
  wire _1487 = r1038 ^ r1154;
  wire _1488 = r1215 ^ r1223;
  wire _1489 = _1487 ^ _1488;
  wire _1490 = r1239 ^ r1304;
  wire _1491 = r1347 ^ r1403;
  wire _1492 = _1490 ^ _1491;
  wire _1493 = _1489 ^ _1492;
  wire _1494 = r1563 ^ r1596;
  wire _1495 = r1613 ^ r1791;
  wire _1496 = _1494 ^ _1495;
  wire _1497 = r1825 ^ r1832;
  wire _1498 = r1861 ^ r1879;
  wire _1499 = _1497 ^ _1498;
  wire _1500 = _1496 ^ _1499;
  wire _1501 = _1493 ^ _1500;
  wire _1502 = _1486 ^ _1501;
  wire _1503 = r8 ^ r155;
  wire _1504 = r253 ^ r373;
  wire _1505 = _1503 ^ _1504;
  wire _1506 = r489 ^ r529;
  wire _1507 = r614 ^ r629;
  wire _1508 = _1506 ^ _1507;
  wire _1509 = _1505 ^ _1508;
  wire _1510 = r811 ^ r942;
  wire _1511 = r946 ^ r1037;
  wire _1512 = _1510 ^ _1511;
  wire _1513 = r1222 ^ r1238;
  wire _1514 = r1346 ^ r1402;
  wire _1515 = _1513 ^ _1514;
  wire _1516 = _1512 ^ _1515;
  wire _1517 = _1509 ^ _1516;
  wire _1518 = r1612 ^ r1652;
  wire _1519 = r1741 ^ r1746;
  wire _1520 = _1518 ^ _1519;
  wire _1521 = r1893 ^ r1896;
  wire _1522 = r1899 ^ r1923;
  wire _1523 = _1521 ^ _1522;
  wire _1524 = _1520 ^ _1523;
  wire _1525 = r1956 ^ r1968;
  wire _1526 = r2001 ^ r2020;
  wire _1527 = _1525 ^ _1526;
  wire _1528 = r2021 ^ r2033;
  wire _1529 = r2044 ^ r2045;
  wire _1530 = _1528 ^ _1529;
  wire _1531 = _1527 ^ _1530;
  wire _1532 = _1524 ^ _1531;
  wire _1533 = _1517 ^ _1532;
  wire _1534 = _1502 | _1533;
  wire _1535 = _1471 | _1534;
  wire _1536 = _1408 | _1535;
  wire _1537 = _1281 | _1536;
  wire _1538 = r7 ^ r154;
  wire _1539 = r322 ^ r372;
  wire _1540 = _1538 ^ _1539;
  wire _1541 = r423 ^ r488;
  wire _1542 = r528 ^ r613;
  wire _1543 = _1541 ^ _1542;
  wire _1544 = _1540 ^ _1543;
  wire _1545 = r704 ^ r775;
  wire _1546 = r810 ^ r941;
  wire _1547 = _1545 ^ _1546;
  wire _1548 = r945 ^ r1036;
  wire _1549 = r1089 ^ r1153;
  wire _1550 = _1548 ^ _1549;
  wire _1551 = _1547 ^ _1550;
  wire _1552 = _1544 ^ _1551;
  wire _1553 = r1221 ^ r1237;
  wire _1554 = r1345 ^ r1401;
  wire _1555 = _1553 ^ _1554;
  wire _1556 = r1562 ^ r1595;
  wire _1557 = r1763 ^ r1796;
  wire _1558 = _1556 ^ _1557;
  wire _1559 = _1555 ^ _1558;
  wire _1560 = r1823 ^ r1887;
  wire _1561 = r1911 ^ r1938;
  wire _1562 = _1560 ^ _1561;
  wire _1563 = r1954 ^ r1979;
  wire _1564 = r2004 ^ r2005;
  wire _1565 = _1563 ^ _1564;
  wire _1566 = _1562 ^ _1565;
  wire _1567 = _1559 ^ _1566;
  wire _1568 = _1552 ^ _1567;
  wire _1569 = r6 ^ r105;
  wire _1570 = r153 ^ r184;
  wire _1571 = _1569 ^ _1570;
  wire _1572 = r252 ^ r321;
  wire _1573 = r371 ^ r422;
  wire _1574 = _1572 ^ _1573;
  wire _1575 = _1571 ^ _1574;
  wire _1576 = r487 ^ r527;
  wire _1577 = r612 ^ r628;
  wire _1578 = _1576 ^ _1577;
  wire _1579 = r703 ^ r774;
  wire _1580 = r809 ^ r866;
  wire _1581 = _1579 ^ _1580;
  wire _1582 = _1578 ^ _1581;
  wire _1583 = _1575 ^ _1582;
  wire _1584 = r940 ^ r944;
  wire _1585 = r1035 ^ r1088;
  wire _1586 = _1584 ^ _1585;
  wire _1587 = r1152 ^ r1214;
  wire _1588 = r1220 ^ r1236;
  wire _1589 = _1587 ^ _1588;
  wire _1590 = _1586 ^ _1589;
  wire _1591 = r1303 ^ r1344;
  wire _1592 = r1400 ^ r1561;
  wire _1593 = _1591 ^ _1592;
  wire _1594 = r1594 ^ r1611;
  wire _1595 = r1651 ^ r1739;
  wire _1596 = _1594 ^ _1595;
  wire _1597 = _1593 ^ _1596;
  wire _1598 = _1590 ^ _1597;
  wire _1599 = _1583 ^ _1598;
  wire _1600 = _1568 | _1599;
  wire _1601 = r5 ^ r104;
  wire _1602 = r152 ^ r183;
  wire _1603 = _1601 ^ _1602;
  wire _1604 = r251 ^ r320;
  wire _1605 = r370 ^ r421;
  wire _1606 = _1604 ^ _1605;
  wire _1607 = _1603 ^ _1606;
  wire _1608 = r486 ^ r526;
  wire _1609 = r611 ^ r627;
  wire _1610 = _1608 ^ _1609;
  wire _1611 = r702 ^ r773;
  wire _1612 = r808 ^ r865;
  wire _1613 = _1611 ^ _1612;
  wire _1614 = _1610 ^ _1613;
  wire _1615 = _1607 ^ _1614;
  wire _1616 = r939 ^ r1002;
  wire _1617 = r1034 ^ r1151;
  wire _1618 = _1616 ^ _1617;
  wire _1619 = r1213 ^ r1219;
  wire _1620 = r1235 ^ r1302;
  wire _1621 = _1619 ^ _1620;
  wire _1622 = _1618 ^ _1621;
  wire _1623 = r1343 ^ r1399;
  wire _1624 = r1560 ^ r1593;
  wire _1625 = _1623 ^ _1624;
  wire _1626 = r1610 ^ r1712;
  wire _1627 = r1777 ^ r1818;
  wire _1628 = _1626 ^ _1627;
  wire _1629 = _1625 ^ _1628;
  wire _1630 = _1622 ^ _1629;
  wire _1631 = _1615 ^ _1630;
  wire _1632 = r4 ^ r103;
  wire _1633 = r182 ^ r250;
  wire _1634 = _1632 ^ _1633;
  wire _1635 = r319 ^ r369;
  wire _1636 = r420 ^ r485;
  wire _1637 = _1635 ^ _1636;
  wire _1638 = _1634 ^ _1637;
  wire _1639 = r525 ^ r610;
  wire _1640 = r626 ^ r701;
  wire _1641 = _1639 ^ _1640;
  wire _1642 = r807 ^ r938;
  wire _1643 = r1001 ^ r1087;
  wire _1644 = _1642 ^ _1643;
  wire _1645 = _1641 ^ _1644;
  wire _1646 = _1638 ^ _1645;
  wire _1647 = r1150 ^ r1218;
  wire _1648 = r1342 ^ r1398;
  wire _1649 = _1647 ^ _1648;
  wire _1650 = r1457 ^ r1592;
  wire _1651 = r1609 ^ r1834;
  wire _1652 = _1650 ^ _1651;
  wire _1653 = _1649 ^ _1652;
  wire _1654 = r1835 ^ r1864;
  wire _1655 = r1866 ^ r1868;
  wire _1656 = _1654 ^ _1655;
  wire _1657 = r1926 ^ r1939;
  wire _1658 = r1998 ^ r2000;
  wire _1659 = _1657 ^ _1658;
  wire _1660 = _1656 ^ _1659;
  wire _1661 = _1653 ^ _1660;
  wire _1662 = _1646 ^ _1661;
  wire _1663 = _1631 | _1662;
  wire _1664 = _1600 | _1663;
  wire _1665 = r102 ^ r151;
  wire _1666 = r181 ^ r318;
  wire _1667 = _1665 ^ _1666;
  wire _1668 = r368 ^ r419;
  wire _1669 = r524 ^ r609;
  wire _1670 = _1668 ^ _1669;
  wire _1671 = _1667 ^ _1670;
  wire _1672 = r625 ^ r700;
  wire _1673 = r772 ^ r806;
  wire _1674 = _1672 ^ _1673;
  wire _1675 = r864 ^ r937;
  wire _1676 = r1000 ^ r1033;
  wire _1677 = _1675 ^ _1676;
  wire _1678 = _1674 ^ _1677;
  wire _1679 = _1671 ^ _1678;
  wire _1680 = r1086 ^ r1149;
  wire _1681 = r1169 ^ r1212;
  wire _1682 = _1680 ^ _1681;
  wire _1683 = r1234 ^ r1301;
  wire _1684 = r1341 ^ r1397;
  wire _1685 = _1683 ^ _1684;
  wire _1686 = _1682 ^ _1685;
  wire _1687 = r1559 ^ r1711;
  wire _1688 = r1872 ^ r1908;
  wire _1689 = _1687 ^ _1688;
  wire _1690 = r1916 ^ r1945;
  wire _1691 = r2024 ^ r2026;
  wire _1692 = _1690 ^ _1691;
  wire _1693 = _1689 ^ _1692;
  wire _1694 = _1686 ^ _1693;
  wire _1695 = _1679 ^ _1694;
  wire _1696 = r3 ^ r150;
  wire _1697 = r180 ^ r249;
  wire _1698 = _1696 ^ _1697;
  wire _1699 = r317 ^ r367;
  wire _1700 = r418 ^ r484;
  wire _1701 = _1699 ^ _1700;
  wire _1702 = _1698 ^ _1701;
  wire _1703 = r608 ^ r699;
  wire _1704 = r771 ^ r863;
  wire _1705 = _1703 ^ _1704;
  wire _1706 = r936 ^ r1032;
  wire _1707 = r1085 ^ r1148;
  wire _1708 = _1706 ^ _1707;
  wire _1709 = _1705 ^ _1708;
  wire _1710 = _1702 ^ _1709;
  wire _1711 = r1168 ^ r1211;
  wire _1712 = r1233 ^ r1340;
  wire _1713 = _1711 ^ _1712;
  wire _1714 = r1396 ^ r1456;
  wire _1715 = r1650 ^ r1776;
  wire _1716 = _1714 ^ _1715;
  wire _1717 = _1713 ^ _1716;
  wire _1718 = r1836 ^ r1905;
  wire _1719 = r1917 ^ r1930;
  wire _1720 = _1718 ^ _1719;
  wire _1721 = r2025 ^ r2031;
  wire _1722 = r2046 ^ r2047;
  wire _1723 = _1721 ^ _1722;
  wire _1724 = _1720 ^ _1723;
  wire _1725 = _1717 ^ _1724;
  wire _1726 = _1710 ^ _1725;
  wire _1727 = _1695 | _1726;
  wire _1728 = r2 ^ r101;
  wire _1729 = r149 ^ r179;
  wire _1730 = _1728 ^ _1729;
  wire _1731 = r316 ^ r366;
  wire _1732 = r417 ^ r523;
  wire _1733 = _1731 ^ _1732;
  wire _1734 = _1730 ^ _1733;
  wire _1735 = r698 ^ r770;
  wire _1736 = r805 ^ r862;
  wire _1737 = _1735 ^ _1736;
  wire _1738 = r935 ^ r999;
  wire _1739 = r1031 ^ r1084;
  wire _1740 = _1738 ^ _1739;
  wire _1741 = _1737 ^ _1740;
  wire _1742 = _1734 ^ _1741;
  wire _1743 = r1147 ^ r1210;
  wire _1744 = r1232 ^ r1300;
  wire _1745 = _1743 ^ _1744;
  wire _1746 = r1339 ^ r1475;
  wire _1747 = r1608 ^ r1649;
  wire _1748 = _1746 ^ _1747;
  wire _1749 = _1745 ^ _1748;
  wire _1750 = r1752 ^ r1785;
  wire _1751 = r1797 ^ r1840;
  wire _1752 = _1750 ^ _1751;
  wire _1753 = r1847 ^ r1890;
  wire _1754 = r1931 ^ r1936;
  wire _1755 = _1753 ^ _1754;
  wire _1756 = _1752 ^ _1755;
  wire _1757 = _1749 ^ _1756;
  wire _1758 = _1742 ^ _1757;
  wire _1759 = r1 ^ r100;
  wire _1760 = r148 ^ r178;
  wire _1761 = _1759 ^ _1760;
  wire _1762 = r248 ^ r315;
  wire _1763 = r365 ^ r416;
  wire _1764 = _1762 ^ _1763;
  wire _1765 = _1761 ^ _1764;
  wire _1766 = r483 ^ r522;
  wire _1767 = r607 ^ r624;
  wire _1768 = _1766 ^ _1767;
  wire _1769 = r697 ^ r769;
  wire _1770 = r804 ^ r861;
  wire _1771 = _1769 ^ _1770;
  wire _1772 = _1768 ^ _1771;
  wire _1773 = _1765 ^ _1772;
  wire _1774 = r934 ^ r998;
  wire _1775 = r1030 ^ r1083;
  wire _1776 = _1774 ^ _1775;
  wire _1777 = r1146 ^ r1167;
  wire _1778 = r1209 ^ r1231;
  wire _1779 = _1777 ^ _1778;
  wire _1780 = _1776 ^ _1779;
  wire _1781 = r1299 ^ r1338;
  wire _1782 = r1395 ^ r1474;
  wire _1783 = _1781 ^ _1782;
  wire _1784 = r1494 ^ r1591;
  wire _1785 = r1710 ^ r1740;
  wire _1786 = _1784 ^ _1785;
  wire _1787 = _1783 ^ _1786;
  wire _1788 = _1780 ^ _1787;
  wire _1789 = _1773 ^ _1788;
  wire _1790 = _1758 | _1789;
  wire _1791 = _1727 | _1790;
  wire _1792 = _1664 | _1791;
  wire _1793 = r0 ^ r99;
  wire _1794 = r147 ^ r177;
  wire _1795 = _1793 ^ _1794;
  wire _1796 = r247 ^ r314;
  wire _1797 = r364 ^ r415;
  wire _1798 = _1796 ^ _1797;
  wire _1799 = _1795 ^ _1798;
  wire _1800 = r482 ^ r521;
  wire _1801 = r606 ^ r623;
  wire _1802 = _1800 ^ _1801;
  wire _1803 = r696 ^ r803;
  wire _1804 = r860 ^ r933;
  wire _1805 = _1803 ^ _1804;
  wire _1806 = _1802 ^ _1805;
  wire _1807 = _1799 ^ _1806;
  wire _1808 = r997 ^ r1029;
  wire _1809 = r1082 ^ r1145;
  wire _1810 = _1808 ^ _1809;
  wire _1811 = r1166 ^ r1208;
  wire _1812 = r1230 ^ r1298;
  wire _1813 = _1811 ^ _1812;
  wire _1814 = _1810 ^ _1813;
  wire _1815 = r1394 ^ r1473;
  wire _1816 = r1493 ^ r1495;
  wire _1817 = _1815 ^ _1816;
  wire _1818 = r1709 ^ r1745;
  wire _1819 = r1789 ^ r1819;
  wire _1820 = _1818 ^ _1819;
  wire _1821 = _1817 ^ _1820;
  wire _1822 = _1814 ^ _1821;
  wire _1823 = _1807 ^ _1822;
  wire _1824 = r98 ^ r146;
  wire _1825 = r176 ^ r246;
  wire _1826 = _1824 ^ _1825;
  wire _1827 = r313 ^ r363;
  wire _1828 = r414 ^ r481;
  wire _1829 = _1827 ^ _1828;
  wire _1830 = _1826 ^ _1829;
  wire _1831 = r520 ^ r605;
  wire _1832 = r622 ^ r695;
  wire _1833 = _1831 ^ _1832;
  wire _1834 = r768 ^ r802;
  wire _1835 = r859 ^ r932;
  wire _1836 = _1834 ^ _1835;
  wire _1837 = _1833 ^ _1836;
  wire _1838 = _1830 ^ _1837;
  wire _1839 = r996 ^ r1081;
  wire _1840 = r1144 ^ r1165;
  wire _1841 = _1839 ^ _1840;
  wire _1842 = r1207 ^ r1229;
  wire _1843 = r1297 ^ r1337;
  wire _1844 = _1842 ^ _1843;
  wire _1845 = _1841 ^ _1844;
  wire _1846 = r1472 ^ r1485;
  wire _1847 = r1590 ^ r1686;
  wire _1848 = _1846 ^ _1847;
  wire _1849 = r1723 ^ r1798;
  wire _1850 = r1804 ^ r1820;
  wire _1851 = _1849 ^ _1850;
  wire _1852 = _1848 ^ _1851;
  wire _1853 = _1845 ^ _1852;
  wire _1854 = _1838 ^ _1853;
  wire _1855 = _1823 | _1854;
  wire _1856 = r97 ^ r145;
  wire _1857 = r175 ^ r312;
  wire _1858 = _1856 ^ _1857;
  wire _1859 = r362 ^ r413;
  wire _1860 = r480 ^ r519;
  wire _1861 = _1859 ^ _1860;
  wire _1862 = _1858 ^ _1861;
  wire _1863 = r604 ^ r621;
  wire _1864 = r694 ^ r767;
  wire _1865 = _1863 ^ _1864;
  wire _1866 = r801 ^ r858;
  wire _1867 = r931 ^ r995;
  wire _1868 = _1866 ^ _1867;
  wire _1869 = _1865 ^ _1868;
  wire _1870 = _1862 ^ _1869;
  wire _1871 = r1028 ^ r1080;
  wire _1872 = r1143 ^ r1164;
  wire _1873 = _1871 ^ _1872;
  wire _1874 = r1206 ^ r1228;
  wire _1875 = r1336 ^ r1393;
  wire _1876 = _1874 ^ _1875;
  wire _1877 = _1873 ^ _1876;
  wire _1878 = r1471 ^ r1589;
  wire _1879 = r1685 ^ r1838;
  wire _1880 = _1878 ^ _1879;
  wire _1881 = r1851 ^ r1870;
  wire _1882 = r1928 ^ r1929;
  wire _1883 = _1881 ^ _1882;
  wire _1884 = _1880 ^ _1883;
  wire _1885 = _1877 ^ _1884;
  wire _1886 = _1870 ^ _1885;
  wire _1887 = r144 ^ r174;
  wire _1888 = r245 ^ r311;
  wire _1889 = _1887 ^ _1888;
  wire _1890 = r361 ^ r412;
  wire _1891 = r479 ^ r603;
  wire _1892 = _1890 ^ _1891;
  wire _1893 = _1889 ^ _1892;
  wire _1894 = r693 ^ r766;
  wire _1895 = r857 ^ r994;
  wire _1896 = _1894 ^ _1895;
  wire _1897 = r1027 ^ r1113;
  wire _1898 = r1142 ^ r1205;
  wire _1899 = _1897 ^ _1898;
  wire _1900 = _1896 ^ _1899;
  wire _1901 = _1893 ^ _1900;
  wire _1902 = r1227 ^ r1296;
  wire _1903 = r1470 ^ r1484;
  wire _1904 = _1902 ^ _1903;
  wire _1905 = r1722 ^ r1751;
  wire _1906 = r1757 ^ r1774;
  wire _1907 = _1905 ^ _1906;
  wire _1908 = _1904 ^ _1907;
  wire _1909 = r1794 ^ r1874;
  wire _1910 = r1920 ^ r1927;
  wire _1911 = _1909 ^ _1910;
  wire _1912 = r1983 ^ r2012;
  wire _1913 = r2015 ^ r2017;
  wire _1914 = _1912 ^ _1913;
  wire _1915 = _1911 ^ _1914;
  wire _1916 = _1908 ^ _1915;
  wire _1917 = _1901 ^ _1916;
  wire _1918 = _1886 | _1917;
  wire _1919 = _1855 | _1918;
  wire _1920 = r96 ^ r143;
  wire _1921 = r173 ^ r244;
  wire _1922 = _1920 ^ _1921;
  wire _1923 = r310 ^ r360;
  wire _1924 = r411 ^ r478;
  wire _1925 = _1923 ^ _1924;
  wire _1926 = _1922 ^ _1925;
  wire _1927 = r518 ^ r692;
  wire _1928 = r765 ^ r800;
  wire _1929 = _1927 ^ _1928;
  wire _1930 = r993 ^ r1026;
  wire _1931 = r1112 ^ r1141;
  wire _1932 = _1930 ^ _1931;
  wire _1933 = _1929 ^ _1932;
  wire _1934 = _1926 ^ _1933;
  wire _1935 = r1204 ^ r1226;
  wire _1936 = r1295 ^ r1469;
  wire _1937 = _1935 ^ _1936;
  wire _1938 = r1492 ^ r1588;
  wire _1939 = r1684 ^ r1721;
  wire _1940 = _1938 ^ _1939;
  wire _1941 = _1937 ^ _1940;
  wire _1942 = r1744 ^ r1768;
  wire _1943 = r1846 ^ r1853;
  wire _1944 = _1942 ^ _1943;
  wire _1945 = r1871 ^ r1883;
  wire _1946 = r1966 ^ r1972;
  wire _1947 = _1945 ^ _1946;
  wire _1948 = _1944 ^ _1947;
  wire _1949 = _1941 ^ _1948;
  wire _1950 = _1934 ^ _1949;
  wire _1951 = r95 ^ r142;
  wire _1952 = r172 ^ r243;
  wire _1953 = _1951 ^ _1952;
  wire _1954 = r309 ^ r359;
  wire _1955 = r410 ^ r477;
  wire _1956 = _1954 ^ _1955;
  wire _1957 = _1953 ^ _1956;
  wire _1958 = r517 ^ r602;
  wire _1959 = r620 ^ r691;
  wire _1960 = _1958 ^ _1959;
  wire _1961 = r764 ^ r856;
  wire _1962 = r930 ^ r992;
  wire _1963 = _1961 ^ _1962;
  wire _1964 = _1960 ^ _1963;
  wire _1965 = _1957 ^ _1964;
  wire _1966 = r1025 ^ r1079;
  wire _1967 = r1110 ^ r1140;
  wire _1968 = _1966 ^ _1967;
  wire _1969 = r1203 ^ r1225;
  wire _1970 = r1294 ^ r1335;
  wire _1971 = _1969 ^ _1970;
  wire _1972 = _1968 ^ _1971;
  wire _1973 = r1392 ^ r1468;
  wire _1974 = r1491 ^ r1683;
  wire _1975 = _1973 ^ _1974;
  wire _1976 = r1719 ^ r1799;
  wire _1977 = r1805 ^ r1821;
  wire _1978 = _1976 ^ _1977;
  wire _1979 = _1975 ^ _1978;
  wire _1980 = _1972 ^ _1979;
  wire _1981 = _1965 ^ _1980;
  wire _1982 = _1950 | _1981;
  wire _1983 = r94 ^ r141;
  wire _1984 = r171 ^ r242;
  wire _1985 = _1983 ^ _1984;
  wire _1986 = r308 ^ r358;
  wire _1987 = r409 ^ r619;
  wire _1988 = _1986 ^ _1987;
  wire _1989 = _1985 ^ _1988;
  wire _1990 = r690 ^ r799;
  wire _1991 = r855 ^ r929;
  wire _1992 = _1990 ^ _1991;
  wire _1993 = r1078 ^ r1108;
  wire _1994 = r1139 ^ r1202;
  wire _1995 = _1993 ^ _1994;
  wire _1996 = _1992 ^ _1995;
  wire _1997 = _1989 ^ _1996;
  wire _1998 = r1293 ^ r1391;
  wire _1999 = r1467 ^ r1490;
  wire _2000 = _1998 ^ _1999;
  wire _2001 = r1524 ^ r1587;
  wire _2002 = r1682 ^ r1720;
  wire _2003 = _2001 ^ _2002;
  wire _2004 = _2000 ^ _2003;
  wire _2005 = r1775 ^ r1779;
  wire _2006 = r1827 ^ r1863;
  wire _2007 = _2005 ^ _2006;
  wire _2008 = r1880 ^ r2010;
  wire _2009 = r2016 ^ r2018;
  wire _2010 = _2008 ^ _2009;
  wire _2011 = _2007 ^ _2010;
  wire _2012 = _2004 ^ _2011;
  wire _2013 = _1997 ^ _2012;
  wire _2014 = r52 ^ r93;
  wire _2015 = r140 ^ r357;
  wire _2016 = _2014 ^ _2015;
  wire _2017 = r516 ^ r601;
  wire _2018 = r618 ^ r763;
  wire _2019 = _2017 ^ _2018;
  wire _2020 = _2016 ^ _2019;
  wire _2021 = r798 ^ r928;
  wire _2022 = r991 ^ r1024;
  wire _2023 = _2021 ^ _2022;
  wire _2024 = r1060 ^ r1201;
  wire _2025 = r1489 ^ r1523;
  wire _2026 = _2024 ^ _2025;
  wire _2027 = _2023 ^ _2026;
  wire _2028 = _2020 ^ _2027;
  wire _2029 = r1551 ^ r1586;
  wire _2030 = r1708 ^ r1761;
  wire _2031 = _2029 ^ _2030;
  wire _2032 = r1783 ^ r1855;
  wire _2033 = r1865 ^ r1949;
  wire _2034 = _2032 ^ _2033;
  wire _2035 = _2031 ^ _2034;
  wire _2036 = r1963 ^ r1967;
  wire _2037 = r1970 ^ r1975;
  wire _2038 = _2036 ^ _2037;
  wire _2039 = r2011 ^ r2039;
  wire _2040 = r2040 ^ r2043;
  wire _2041 = _2039 ^ _2040;
  wire _2042 = _2038 ^ _2041;
  wire _2043 = _2035 ^ _2042;
  wire _2044 = _2028 ^ _2043;
  wire _2045 = _2013 | _2044;
  wire _2046 = _1982 | _2045;
  wire _2047 = _1919 | _2046;
  wire _2048 = _1792 | _2047;
  wire _2049 = _1537 | _2048;
  wire _2050 = _1026 | _2049;
  wire _2051 = r53 ^ r109;
  wire _2052 = r130 ^ r245;
  wire _2053 = _2051 ^ _2052;
  wire _2054 = r299 ^ r342;
  wire _2055 = r442 ^ r458;
  wire _2056 = _2054 ^ _2055;
  wire _2057 = _2053 ^ _2056;
  wire _2058 = r535 ^ r580;
  wire _2059 = r641 ^ r763;
  wire _2060 = _2058 ^ _2059;
  wire _2061 = r796 ^ r859;
  wire _2062 = r894 ^ r944;
  wire _2063 = _2061 ^ _2062;
  wire _2064 = _2060 ^ _2063;
  wire _2065 = _2057 ^ _2064;
  wire _2066 = r1038 ^ r1074;
  wire _2067 = r1158 ^ r1171;
  wire _2068 = _2066 ^ _2067;
  wire _2069 = r1245 ^ r1287;
  wire _2070 = r1346 ^ r1416;
  wire _2071 = _2069 ^ _2070;
  wire _2072 = _2068 ^ _2071;
  wire _2073 = r1574 ^ r1582;
  wire _2074 = r1664 ^ r1740;
  wire _2075 = _2073 ^ _2074;
  wire _2076 = r1902 ^ r1960;
  wire _2077 = r1992 ^ r1994;
  wire _2078 = _2076 ^ _2077;
  wire _2079 = _2075 ^ _2078;
  wire _2080 = _2072 ^ _2079;
  wire _2081 = _2065 ^ _2080;
  wire _2082 = r51 ^ r74;
  wire _2083 = r141 ^ r189;
  wire _2084 = _2082 ^ _2083;
  wire _2085 = r286 ^ r386;
  wire _2086 = r399 ^ r478;
  wire _2087 = _2085 ^ _2086;
  wire _2088 = _2084 ^ _2087;
  wire _2089 = r521 ^ r587;
  wire _2090 = r655 ^ r707;
  wire _2091 = _2089 ^ _2090;
  wire _2092 = r757 ^ r787;
  wire _2093 = r943 ^ r982;
  wire _2094 = _2092 ^ _2093;
  wire _2095 = _2091 ^ _2094;
  wire _2096 = _2088 ^ _2095;
  wire _2097 = r1015 ^ r1100;
  wire _2098 = r1190 ^ r1231;
  wire _2099 = _2097 ^ _2098;
  wire _2100 = r1360 ^ r1402;
  wire _2101 = r1466 ^ r1557;
  wire _2102 = _2100 ^ _2101;
  wire _2103 = _2099 ^ _2102;
  wire _2104 = r1621 ^ r1669;
  wire _2105 = r1718 ^ r1787;
  wire _2106 = _2104 ^ _2105;
  wire _2107 = r1851 ^ r1855;
  wire _2108 = r1978 ^ r1980;
  wire _2109 = _2107 ^ _2108;
  wire _2110 = _2106 ^ _2109;
  wire _2111 = _2103 ^ _2110;
  wire _2112 = _2096 ^ _2111;
  wire _2113 = _2081 | _2112;
  wire _2114 = r50 ^ r66;
  wire _2115 = r155 ^ r244;
  wire _2116 = _2114 ^ _2115;
  wire _2117 = r404 ^ r480;
  wire _2118 = r531 ^ r609;
  wire _2119 = _2117 ^ _2118;
  wire _2120 = _2116 ^ _2119;
  wire _2121 = r666 ^ r701;
  wire _2122 = r751 ^ r871;
  wire _2123 = _2121 ^ _2122;
  wire _2124 = r933 ^ r973;
  wire _2125 = r1045 ^ r1065;
  wire _2126 = _2124 ^ _2125;
  wire _2127 = _2123 ^ _2126;
  wire _2128 = _2120 ^ _2127;
  wire _2129 = r1144 ^ r1174;
  wire _2130 = r1265 ^ r1322;
  wire _2131 = _2129 ^ _2130;
  wire _2132 = r1391 ^ r1606;
  wire _2133 = r1675 ^ r1705;
  wire _2134 = _2132 ^ _2133;
  wire _2135 = _2131 ^ _2134;
  wire _2136 = r1854 ^ r1860;
  wire _2137 = r1875 ^ r1930;
  wire _2138 = _2136 ^ _2137;
  wire _2139 = r1940 ^ r1995;
  wire _2140 = r2011 ^ r2019;
  wire _2141 = _2139 ^ _2140;
  wire _2142 = _2138 ^ _2141;
  wire _2143 = _2135 ^ _2142;
  wire _2144 = _2128 ^ _2143;
  wire _2145 = r97 ^ r275;
  wire _2146 = r322 ^ r365;
  wire _2147 = _2145 ^ _2146;
  wire _2148 = r393 ^ r449;
  wire _2149 = r524 ^ r561;
  wire _2150 = _2148 ^ _2149;
  wire _2151 = _2147 ^ _2150;
  wire _2152 = r638 ^ r734;
  wire _2153 = r874 ^ r960;
  wire _2154 = _2152 ^ _2153;
  wire _2155 = r1003 ^ r1042;
  wire _2156 = r1069 ^ r1154;
  wire _2157 = _2155 ^ _2156;
  wire _2158 = _2154 ^ _2157;
  wire _2159 = _2151 ^ _2158;
  wire _2160 = r1248 ^ r1313;
  wire _2161 = r1353 ^ r1405;
  wire _2162 = _2160 ^ _2161;
  wire _2163 = r1483 ^ r1500;
  wire _2164 = r1561 ^ r1702;
  wire _2165 = _2163 ^ _2164;
  wire _2166 = _2162 ^ _2165;
  wire _2167 = r1811 ^ r1812;
  wire _2168 = r1833 ^ r1849;
  wire _2169 = _2167 ^ _2168;
  wire _2170 = r1900 ^ r1926;
  wire _2171 = r2014 ^ r2020;
  wire _2172 = _2170 ^ _2171;
  wire _2173 = _2169 ^ _2172;
  wire _2174 = _2166 ^ _2173;
  wire _2175 = _2159 ^ _2174;
  wire _2176 = _2144 | _2175;
  wire _2177 = _2113 | _2176;
  wire _2178 = r49 ^ r112;
  wire _2179 = r210 ^ r256;
  wire _2180 = _2178 ^ _2179;
  wire _2181 = r318 ^ r381;
  wire _2182 = r417 ^ r485;
  wire _2183 = _2181 ^ _2182;
  wire _2184 = _2180 ^ _2183;
  wire _2185 = r528 ^ r601;
  wire _2186 = r627 ^ r694;
  wire _2187 = _2185 ^ _2186;
  wire _2188 = r741 ^ r791;
  wire _2189 = r861 ^ r897;
  wire _2190 = _2188 ^ _2189;
  wire _2191 = _2187 ^ _2190;
  wire _2192 = _2184 ^ _2191;
  wire _2193 = r979 ^ r1148;
  wire _2194 = r1195 ^ r1260;
  wire _2195 = _2193 ^ _2194;
  wire _2196 = r1350 ^ r1424;
  wire _2197 = r1442 ^ r1485;
  wire _2198 = _2196 ^ _2197;
  wire _2199 = _2195 ^ _2198;
  wire _2200 = r1504 ^ r1509;
  wire _2201 = r1529 ^ r1556;
  wire _2202 = _2200 ^ _2201;
  wire _2203 = r1578 ^ r1676;
  wire _2204 = r1690 ^ r1741;
  wire _2205 = _2203 ^ _2204;
  wire _2206 = _2202 ^ _2205;
  wire _2207 = _2199 ^ _2206;
  wire _2208 = _2192 ^ _2207;
  wire _2209 = r48 ^ r101;
  wire _2210 = r135 ^ r215;
  wire _2211 = _2209 ^ _2210;
  wire _2212 = r259 ^ r283;
  wire _2213 = r351 ^ r498;
  wire _2214 = _2212 ^ _2213;
  wire _2215 = _2211 ^ _2214;
  wire _2216 = r602 ^ r674;
  wire _2217 = r785 ^ r836;
  wire _2218 = _2216 ^ _2217;
  wire _2219 = r910 ^ r951;
  wire _2220 = r1051 ^ r1152;
  wire _2221 = _2219 ^ _2220;
  wire _2222 = _2218 ^ _2221;
  wire _2223 = _2215 ^ _2222;
  wire _2224 = r1272 ^ r1282;
  wire _2225 = r1364 ^ r1517;
  wire _2226 = _2224 ^ _2225;
  wire _2227 = r1540 ^ r1563;
  wire _2228 = r1607 ^ r1759;
  wire _2229 = _2227 ^ _2228;
  wire _2230 = _2226 ^ _2229;
  wire _2231 = r1773 ^ r1779;
  wire _2232 = r1839 ^ r1948;
  wire _2233 = _2231 ^ _2232;
  wire _2234 = r1951 ^ r1982;
  wire _2235 = r2015 ^ r2021;
  wire _2236 = _2234 ^ _2235;
  wire _2237 = _2233 ^ _2236;
  wire _2238 = _2230 ^ _2237;
  wire _2239 = _2223 ^ _2238;
  wire _2240 = _2208 | _2239;
  wire _2241 = r47 ^ r104;
  wire _2242 = r136 ^ r206;
  wire _2243 = _2241 ^ _2242;
  wire _2244 = r246 ^ r301;
  wire _2245 = r389 ^ r407;
  wire _2246 = _2244 ^ _2245;
  wire _2247 = _2243 ^ _2246;
  wire _2248 = r450 ^ r556;
  wire _2249 = r572 ^ r629;
  wire _2250 = _2248 ^ _2249;
  wire _2251 = r713 ^ r762;
  wire _2252 = r822 ^ r857;
  wire _2253 = _2251 ^ _2252;
  wire _2254 = _2250 ^ _2253;
  wire _2255 = _2247 ^ _2254;
  wire _2256 = r921 ^ r948;
  wire _2257 = r1025 ^ r1063;
  wire _2258 = _2256 ^ _2257;
  wire _2259 = r1141 ^ r1212;
  wire _2260 = r1242 ^ r1388;
  wire _2261 = _2259 ^ _2260;
  wire _2262 = _2258 ^ _2261;
  wire _2263 = r1448 ^ r1495;
  wire _2264 = r1532 ^ r1577;
  wire _2265 = _2263 ^ _2264;
  wire _2266 = r1614 ^ r1708;
  wire _2267 = r1786 ^ r1822;
  wire _2268 = _2266 ^ _2267;
  wire _2269 = _2265 ^ _2268;
  wire _2270 = _2262 ^ _2269;
  wire _2271 = _2255 ^ _2270;
  wire _2272 = r46 ^ r95;
  wire _2273 = r176 ^ r276;
  wire _2274 = _2272 ^ _2273;
  wire _2275 = r302 ^ r353;
  wire _2276 = r479 ^ r538;
  wire _2277 = _2275 ^ _2276;
  wire _2278 = _2274 ^ _2277;
  wire _2279 = r650 ^ r739;
  wire _2280 = r828 ^ r883;
  wire _2281 = _2279 ^ _2280;
  wire _2282 = r891 ^ r964;
  wire _2283 = r1034 ^ r1121;
  wire _2284 = _2282 ^ _2283;
  wire _2285 = _2281 ^ _2284;
  wire _2286 = _2278 ^ _2285;
  wire _2287 = r1198 ^ r1233;
  wire _2288 = r1284 ^ r1431;
  wire _2289 = _2287 ^ _2288;
  wire _2290 = r1452 ^ r1481;
  wire _2291 = r1541 ^ r1651;
  wire _2292 = _2290 ^ _2291;
  wire _2293 = _2289 ^ _2292;
  wire _2294 = r1707 ^ r1813;
  wire _2295 = r1847 ^ r1937;
  wire _2296 = _2294 ^ _2295;
  wire _2297 = r1952 ^ r2018;
  wire _2298 = r2030 ^ r2039;
  wire _2299 = _2297 ^ _2298;
  wire _2300 = _2296 ^ _2299;
  wire _2301 = _2293 ^ _2300;
  wire _2302 = _2286 ^ _2301;
  wire _2303 = _2271 | _2302;
  wire _2304 = _2240 | _2303;
  wire _2305 = _2177 | _2304;
  wire _2306 = r45 ^ r75;
  wire _2307 = r162 ^ r183;
  wire _2308 = _2306 ^ _2307;
  wire _2309 = r243 ^ r367;
  wire _2310 = r435 ^ r493;
  wire _2311 = _2309 ^ _2310;
  wire _2312 = _2308 ^ _2311;
  wire _2313 = r552 ^ r565;
  wire _2314 = r657 ^ r680;
  wire _2315 = _2313 ^ _2314;
  wire _2316 = r775 ^ r867;
  wire _2317 = r935 ^ r957;
  wire _2318 = _2316 ^ _2317;
  wire _2319 = _2315 ^ _2318;
  wire _2320 = _2312 ^ _2319;
  wire _2321 = r1104 ^ r1161;
  wire _2322 = r1214 ^ r1275;
  wire _2323 = _2321 ^ _2322;
  wire _2324 = r1342 ^ r1423;
  wire _2325 = r1527 ^ r1603;
  wire _2326 = _2324 ^ _2325;
  wire _2327 = _2323 ^ _2326;
  wire _2328 = r1629 ^ r1679;
  wire _2329 = r1724 ^ r1820;
  wire _2330 = _2328 ^ _2329;
  wire _2331 = r1848 ^ r1986;
  wire _2332 = r2003 ^ r2008;
  wire _2333 = _2331 ^ _2332;
  wire _2334 = _2330 ^ _2333;
  wire _2335 = _2327 ^ _2334;
  wire _2336 = _2320 ^ _2335;
  wire _2337 = r44 ^ r56;
  wire _2338 = r121 ^ r219;
  wire _2339 = _2337 ^ _2338;
  wire _2340 = r328 ^ r363;
  wire _2341 = r415 ^ r507;
  wire _2342 = _2340 ^ _2341;
  wire _2343 = _2339 ^ _2342;
  wire _2344 = r573 ^ r708;
  wire _2345 = r723 ^ r795;
  wire _2346 = _2344 ^ _2345;
  wire _2347 = r838 ^ r923;
  wire _2348 = r990 ^ r1032;
  wire _2349 = _2347 ^ _2348;
  wire _2350 = _2346 ^ _2349;
  wire _2351 = _2343 ^ _2350;
  wire _2352 = r1075 ^ r1116;
  wire _2353 = r1178 ^ r1235;
  wire _2354 = _2352 ^ _2353;
  wire _2355 = r1311 ^ r1336;
  wire _2356 = r1432 ^ r1451;
  wire _2357 = _2355 ^ _2356;
  wire _2358 = _2354 ^ _2357;
  wire _2359 = r1462 ^ r1619;
  wire _2360 = r1739 ^ r1837;
  wire _2361 = _2359 ^ _2360;
  wire _2362 = r1857 ^ r1914;
  wire _2363 = r1920 ^ r1921;
  wire _2364 = _2362 ^ _2363;
  wire _2365 = _2361 ^ _2364;
  wire _2366 = _2358 ^ _2365;
  wire _2367 = _2351 ^ _2366;
  wire _2368 = _2336 | _2367;
  wire _2369 = r43 ^ r70;
  wire _2370 = r125 ^ r221;
  wire _2371 = _2369 ^ _2370;
  wire _2372 = r290 ^ r384;
  wire _2373 = r427 ^ r501;
  wire _2374 = _2372 ^ _2373;
  wire _2375 = _2371 ^ _2374;
  wire _2376 = r532 ^ r658;
  wire _2377 = r696 ^ r764;
  wire _2378 = _2376 ^ _2377;
  wire _2379 = r885 ^ r938;
  wire _2380 = r1023 ^ r1073;
  wire _2381 = _2379 ^ _2380;
  wire _2382 = _2378 ^ _2381;
  wire _2383 = _2375 ^ _2382;
  wire _2384 = r1127 ^ r1187;
  wire _2385 = r1254 ^ r1318;
  wire _2386 = _2384 ^ _2385;
  wire _2387 = r1339 ^ r1387;
  wire _2388 = r1397 ^ r1446;
  wire _2389 = _2387 ^ _2388;
  wire _2390 = _2386 ^ _2389;
  wire _2391 = r1583 ^ r1634;
  wire _2392 = r1658 ^ r1758;
  wire _2393 = _2391 ^ _2392;
  wire _2394 = r1791 ^ r1796;
  wire _2395 = r1836 ^ r1880;
  wire _2396 = _2394 ^ _2395;
  wire _2397 = _2393 ^ _2396;
  wire _2398 = _2390 ^ _2397;
  wire _2399 = _2383 ^ _2398;
  wire _2400 = r42 ^ r81;
  wire _2401 = r170 ^ r192;
  wire _2402 = _2400 ^ _2401;
  wire _2403 = r278 ^ r294;
  wire _2404 = r347 ^ r436;
  wire _2405 = _2403 ^ _2404;
  wire _2406 = _2402 ^ _2405;
  wire _2407 = r468 ^ r520;
  wire _2408 = r615 ^ r649;
  wire _2409 = _2407 ^ _2408;
  wire _2410 = r682 ^ r740;
  wire _2411 = r807 ^ r872;
  wire _2412 = _2410 ^ _2411;
  wire _2413 = _2409 ^ _2412;
  wire _2414 = _2406 ^ _2413;
  wire _2415 = r903 ^ r993;
  wire _2416 = r1004 ^ r1102;
  wire _2417 = _2415 ^ _2416;
  wire _2418 = r1155 ^ r1183;
  wire _2419 = r1262 ^ r1279;
  wire _2420 = _2418 ^ _2419;
  wire _2421 = _2417 ^ _2420;
  wire _2422 = r1288 ^ r1468;
  wire _2423 = r1534 ^ r1545;
  wire _2424 = _2422 ^ _2423;
  wire _2425 = r1581 ^ r1685;
  wire _2426 = r1775 ^ r1823;
  wire _2427 = _2425 ^ _2426;
  wire _2428 = _2424 ^ _2427;
  wire _2429 = _2421 ^ _2428;
  wire _2430 = _2414 ^ _2429;
  wire _2431 = _2399 | _2430;
  wire _2432 = _2368 | _2431;
  wire _2433 = r41 ^ r106;
  wire _2434 = r124 ^ r174;
  wire _2435 = _2433 ^ _2434;
  wire _2436 = r270 ^ r332;
  wire _2437 = r348 ^ r408;
  wire _2438 = _2436 ^ _2437;
  wire _2439 = _2435 ^ _2438;
  wire _2440 = r481 ^ r509;
  wire _2441 = r588 ^ r619;
  wire _2442 = _2440 ^ _2441;
  wire _2443 = r699 ^ r761;
  wire _2444 = r810 ^ r835;
  wire _2445 = _2443 ^ _2444;
  wire _2446 = _2442 ^ _2445;
  wire _2447 = _2439 ^ _2446;
  wire _2448 = r912 ^ r997;
  wire _2449 = r1041 ^ r1086;
  wire _2450 = _2448 ^ _2449;
  wire _2451 = r1143 ^ r1188;
  wire _2452 = r1257 ^ r1286;
  wire _2453 = _2451 ^ _2452;
  wire _2454 = _2450 ^ _2453;
  wire _2455 = r1365 ^ r1460;
  wire _2456 = r1475 ^ r1547;
  wire _2457 = _2455 ^ _2456;
  wire _2458 = r1609 ^ r1653;
  wire _2459 = r1694 ^ r1742;
  wire _2460 = _2458 ^ _2459;
  wire _2461 = _2457 ^ _2460;
  wire _2462 = _2454 ^ _2461;
  wire _2463 = _2447 ^ _2462;
  wire _2464 = r119 ^ r185;
  wire _2465 = r257 ^ r293;
  wire _2466 = _2464 ^ _2465;
  wire _2467 = r383 ^ r423;
  wire _2468 = r477 ^ r523;
  wire _2469 = _2467 ^ _2468;
  wire _2470 = _2466 ^ _2469;
  wire _2471 = r568 ^ r624;
  wire _2472 = r717 ^ r722;
  wire _2473 = _2471 ^ _2472;
  wire _2474 = r731 ^ r797;
  wire _2475 = r865 ^ r908;
  wire _2476 = _2474 ^ _2475;
  wire _2477 = _2473 ^ _2476;
  wire _2478 = _2470 ^ _2477;
  wire _2479 = r987 ^ r1055;
  wire _2480 = r1088 ^ r1177;
  wire _2481 = _2479 ^ _2480;
  wire _2482 = r1263 ^ r1316;
  wire _2483 = r1349 ^ r1409;
  wire _2484 = _2482 ^ _2483;
  wire _2485 = _2481 ^ _2484;
  wire _2486 = r1435 ^ r1624;
  wire _2487 = r1659 ^ r1810;
  wire _2488 = _2486 ^ _2487;
  wire _2489 = r1845 ^ r2013;
  wire _2490 = r2017 ^ r2031;
  wire _2491 = _2489 ^ _2490;
  wire _2492 = _2488 ^ _2491;
  wire _2493 = _2485 ^ _2492;
  wire _2494 = _2478 ^ _2493;
  wire _2495 = _2463 | _2494;
  wire _2496 = r40 ^ r84;
  wire _2497 = r159 ^ r193;
  wire _2498 = _2496 ^ _2497;
  wire _2499 = r274 ^ r288;
  wire _2500 = r374 ^ r391;
  wire _2501 = _2499 ^ _2500;
  wire _2502 = _2498 ^ _2501;
  wire _2503 = r395 ^ r496;
  wire _2504 = r544 ^ r590;
  wire _2505 = _2503 ^ _2504;
  wire _2506 = r662 ^ r672;
  wire _2507 = r772 ^ r827;
  wire _2508 = _2506 ^ _2507;
  wire _2509 = _2505 ^ _2508;
  wire _2510 = _2502 ^ _2509;
  wire _2511 = r863 ^ r913;
  wire _2512 = r965 ^ r1009;
  wire _2513 = _2511 ^ _2512;
  wire _2514 = r1076 ^ r1146;
  wire _2515 = r1200 ^ r1253;
  wire _2516 = _2514 ^ _2515;
  wire _2517 = _2513 ^ _2516;
  wire _2518 = r1300 ^ r1361;
  wire _2519 = r1392 ^ r1437;
  wire _2520 = _2518 ^ _2519;
  wire _2521 = r1593 ^ r1616;
  wire _2522 = r1680 ^ r1743;
  wire _2523 = _2521 ^ _2522;
  wire _2524 = _2520 ^ _2523;
  wire _2525 = _2517 ^ _2524;
  wire _2526 = _2510 ^ _2525;
  wire _2527 = r39 ^ r99;
  wire _2528 = r167 ^ r220;
  wire _2529 = _2527 ^ _2528;
  wire _2530 = r325 ^ r430;
  wire _2531 = r463 ^ r721;
  wire _2532 = _2530 ^ _2531;
  wire _2533 = _2529 ^ _2532;
  wire _2534 = r742 ^ r794;
  wire _2535 = r902 ^ r947;
  wire _2536 = _2534 ^ _2535;
  wire _2537 = r1035 ^ r1103;
  wire _2538 = r1207 ^ r1331;
  wire _2539 = _2537 ^ _2538;
  wire _2540 = _2536 ^ _2539;
  wire _2541 = _2533 ^ _2540;
  wire _2542 = r1371 ^ r1401;
  wire _2543 = r1512 ^ r1521;
  wire _2544 = _2542 ^ _2543;
  wire _2545 = r1567 ^ r1727;
  wire _2546 = r1769 ^ r1776;
  wire _2547 = _2545 ^ _2546;
  wire _2548 = _2544 ^ _2547;
  wire _2549 = r1777 ^ r1801;
  wire _2550 = r1866 ^ r1883;
  wire _2551 = _2549 ^ _2550;
  wire _2552 = r1891 ^ r1950;
  wire _2553 = r2026 ^ r2032;
  wire _2554 = _2552 ^ _2553;
  wire _2555 = _2551 ^ _2554;
  wire _2556 = _2548 ^ _2555;
  wire _2557 = _2541 ^ _2556;
  wire _2558 = _2526 | _2557;
  wire _2559 = _2495 | _2558;
  wire _2560 = _2432 | _2559;
  wire _2561 = _2305 | _2560;
  wire _2562 = r38 ^ r62;
  wire _2563 = r131 ^ r182;
  wire _2564 = _2562 ^ _2563;
  wire _2565 = r248 ^ r337;
  wire _2566 = r397 ^ r549;
  wire _2567 = _2565 ^ _2566;
  wire _2568 = _2564 ^ _2567;
  wire _2569 = r600 ^ r632;
  wire _2570 = r673 ^ r733;
  wire _2571 = _2569 ^ _2570;
  wire _2572 = r869 ^ r926;
  wire _2573 = r961 ^ r1072;
  wire _2574 = _2572 ^ _2573;
  wire _2575 = _2571 ^ _2574;
  wire _2576 = _2568 ^ _2575;
  wire _2577 = r1118 ^ r1166;
  wire _2578 = r1192 ^ r1228;
  wire _2579 = _2577 ^ _2578;
  wire _2580 = r1289 ^ r1343;
  wire _2581 = r1410 ^ r1461;
  wire _2582 = _2580 ^ _2581;
  wire _2583 = _2579 ^ _2582;
  wire _2584 = r1484 ^ r1695;
  wire _2585 = r1730 ^ r1915;
  wire _2586 = _2584 ^ _2585;
  wire _2587 = r1961 ^ r1967;
  wire _2588 = r2010 ^ r2022;
  wire _2589 = _2587 ^ _2588;
  wire _2590 = _2586 ^ _2589;
  wire _2591 = _2583 ^ _2590;
  wire _2592 = _2576 ^ _2591;
  wire _2593 = r37 ^ r72;
  wire _2594 = r129 ^ r262;
  wire _2595 = _2593 ^ _2594;
  wire _2596 = r409 ^ r495;
  wire _2597 = r554 ^ r563;
  wire _2598 = _2596 ^ _2597;
  wire _2599 = _2595 ^ _2598;
  wire _2600 = r617 ^ r804;
  wire _2601 = r846 ^ r972;
  wire _2602 = _2600 ^ _2601;
  wire _2603 = r1012 ^ r1095;
  wire _2604 = r1114 ^ r1168;
  wire _2605 = _2603 ^ _2604;
  wire _2606 = _2602 ^ _2605;
  wire _2607 = _2599 ^ _2606;
  wire _2608 = r1267 ^ r1317;
  wire _2609 = r1496 ^ r1546;
  wire _2610 = _2608 ^ _2609;
  wire _2611 = r1560 ^ r1580;
  wire _2612 = r1647 ^ r1655;
  wire _2613 = _2611 ^ _2612;
  wire _2614 = _2610 ^ _2613;
  wire _2615 = r1867 ^ r1874;
  wire _2616 = r1878 ^ r1949;
  wire _2617 = _2615 ^ _2616;
  wire _2618 = r1956 ^ r1957;
  wire _2619 = r1971 ^ r1973;
  wire _2620 = _2618 ^ _2619;
  wire _2621 = _2617 ^ _2620;
  wire _2622 = _2614 ^ _2621;
  wire _2623 = _2607 ^ _2622;
  wire _2624 = _2592 | _2623;
  wire _2625 = r36 ^ r67;
  wire _2626 = r165 ^ r188;
  wire _2627 = _2625 ^ _2626;
  wire _2628 = r254 ^ r298;
  wire _2629 = r336 ^ r486;
  wire _2630 = _2628 ^ _2629;
  wire _2631 = _2627 ^ _2630;
  wire _2632 = r543 ^ r584;
  wire _2633 = r626 ^ r685;
  wire _2634 = _2632 ^ _2633;
  wire _2635 = r738 ^ r777;
  wire _2636 = r829 ^ r856;
  wire _2637 = _2635 ^ _2636;
  wire _2638 = _2634 ^ _2637;
  wire _2639 = _2631 ^ _2638;
  wire _2640 = r916 ^ r1000;
  wire _2641 = r1027 ^ r1082;
  wire _2642 = _2640 ^ _2641;
  wire _2643 = r1119 ^ r1216;
  wire _2644 = r1269 ^ r1374;
  wire _2645 = _2643 ^ _2644;
  wire _2646 = _2642 ^ _2645;
  wire _2647 = r1396 ^ r1490;
  wire _2648 = r1568 ^ r1601;
  wire _2649 = _2647 ^ _2648;
  wire _2650 = r1670 ^ r1763;
  wire _2651 = r1788 ^ r1824;
  wire _2652 = _2650 ^ _2651;
  wire _2653 = _2649 ^ _2652;
  wire _2654 = _2646 ^ _2653;
  wire _2655 = _2639 ^ _2654;
  wire _2656 = r35 ^ r73;
  wire _2657 = r144 ^ r208;
  wire _2658 = _2656 ^ _2657;
  wire _2659 = r232 ^ r330;
  wire _2660 = r425 ^ r448;
  wire _2661 = _2659 ^ _2660;
  wire _2662 = _2658 ^ _2661;
  wire _2663 = r511 ^ r585;
  wire _2664 = r633 ^ r691;
  wire _2665 = _2663 ^ _2664;
  wire _2666 = r821 ^ r850;
  wire _2667 = r918 ^ r989;
  wire _2668 = _2666 ^ _2667;
  wire _2669 = _2665 ^ _2668;
  wire _2670 = _2662 ^ _2669;
  wire _2671 = r1047 ^ r1105;
  wire _2672 = r1239 ^ r1309;
  wire _2673 = _2671 ^ _2672;
  wire _2674 = r1332 ^ r1425;
  wire _2675 = r1436 ^ r1511;
  wire _2676 = _2674 ^ _2675;
  wire _2677 = _2673 ^ _2676;
  wire _2678 = r1590 ^ r1641;
  wire _2679 = r1681 ^ r1693;
  wire _2680 = _2678 ^ _2679;
  wire _2681 = r1819 ^ r1871;
  wire _2682 = r1919 ^ r1922;
  wire _2683 = _2681 ^ _2682;
  wire _2684 = _2680 ^ _2683;
  wire _2685 = _2677 ^ _2684;
  wire _2686 = _2670 ^ _2685;
  wire _2687 = _2655 | _2686;
  wire _2688 = _2624 | _2687;
  wire _2689 = r34 ^ r61;
  wire _2690 = r147 ^ r222;
  wire _2691 = _2689 ^ _2690;
  wire _2692 = r310 ^ r371;
  wire _2693 = r392 ^ r453;
  wire _2694 = _2692 ^ _2693;
  wire _2695 = _2691 ^ _2694;
  wire _2696 = r562 ^ r663;
  wire _2697 = r676 ^ r766;
  wire _2698 = _2696 ^ _2697;
  wire _2699 = r808 ^ r854;
  wire _2700 = r942 ^ r975;
  wire _2701 = _2699 ^ _2700;
  wire _2702 = _2698 ^ _2701;
  wire _2703 = _2695 ^ _2702;
  wire _2704 = r1057 ^ r1097;
  wire _2705 = r1132 ^ r1211;
  wire _2706 = _2704 ^ _2705;
  wire _2707 = r1404 ^ r1455;
  wire _2708 = r1463 ^ r1474;
  wire _2709 = _2707 ^ _2708;
  wire _2710 = _2706 ^ _2709;
  wire _2711 = r1625 ^ r1678;
  wire _2712 = r1761 ^ r1804;
  wire _2713 = _2711 ^ _2712;
  wire _2714 = r1863 ^ r1870;
  wire _2715 = r1897 ^ r1907;
  wire _2716 = _2714 ^ _2715;
  wire _2717 = _2713 ^ _2716;
  wire _2718 = _2710 ^ _2717;
  wire _2719 = _2703 ^ _2718;
  wire _2720 = r33 ^ r132;
  wire _2721 = r218 ^ r235;
  wire _2722 = _2720 ^ _2721;
  wire _2723 = r313 ^ r379;
  wire _2724 = r505 ^ r558;
  wire _2725 = _2723 ^ _2724;
  wire _2726 = _2722 ^ _2725;
  wire _2727 = r608 ^ r623;
  wire _2728 = r677 ^ r725;
  wire _2729 = _2727 ^ _2728;
  wire _2730 = r843 ^ r924;
  wire _2731 = r1052 ^ r1087;
  wire _2732 = _2730 ^ _2731;
  wire _2733 = _2729 ^ _2732;
  wire _2734 = _2726 ^ _2733;
  wire _2735 = r1217 ^ r1232;
  wire _2736 = r1277 ^ r1319;
  wire _2737 = _2735 ^ _2736;
  wire _2738 = r1363 ^ r1389;
  wire _2739 = r1652 ^ r1768;
  wire _2740 = _2738 ^ _2739;
  wire _2741 = _2737 ^ _2740;
  wire _2742 = r1770 ^ r1772;
  wire _2743 = r1815 ^ r1872;
  wire _2744 = _2742 ^ _2743;
  wire _2745 = r1909 ^ r2016;
  wire _2746 = r2038 ^ r2043;
  wire _2747 = _2745 ^ _2746;
  wire _2748 = _2744 ^ _2747;
  wire _2749 = _2741 ^ _2748;
  wire _2750 = _2734 ^ _2749;
  wire _2751 = _2719 | _2750;
  wire _2752 = r32 ^ r166;
  wire _2753 = r239 ^ r343;
  wire _2754 = _2752 ^ _2753;
  wire _2755 = r424 ^ r452;
  wire _2756 = r559 ^ r571;
  wire _2757 = _2755 ^ _2756;
  wire _2758 = _2754 ^ _2757;
  wire _2759 = r651 ^ r703;
  wire _2760 = r773 ^ r877;
  wire _2761 = _2759 ^ _2760;
  wire _2762 = r934 ^ r953;
  wire _2763 = r1058 ^ r1101;
  wire _2764 = _2762 ^ _2763;
  wire _2765 = _2761 ^ _2764;
  wire _2766 = _2758 ^ _2765;
  wire _2767 = r1112 ^ r1122;
  wire _2768 = r1310 ^ r1358;
  wire _2769 = _2767 ^ _2768;
  wire _2770 = r1620 ^ r1756;
  wire _2771 = r1762 ^ r1802;
  wire _2772 = _2770 ^ _2771;
  wire _2773 = _2769 ^ _2772;
  wire _2774 = r1916 ^ r1944;
  wire _2775 = r1946 ^ r1954;
  wire _2776 = _2774 ^ _2775;
  wire _2777 = r1983 ^ r1993;
  wire _2778 = r1996 ^ r2001;
  wire _2779 = _2777 ^ _2778;
  wire _2780 = _2776 ^ _2779;
  wire _2781 = _2773 ^ _2780;
  wire _2782 = _2766 ^ _2781;
  wire _2783 = r31 ^ r77;
  wire _2784 = r128 ^ r203;
  wire _2785 = _2783 ^ _2784;
  wire _2786 = r229 ^ r331;
  wire _2787 = r341 ^ r416;
  wire _2788 = _2786 ^ _2787;
  wire _2789 = _2785 ^ _2788;
  wire _2790 = r503 ^ r526;
  wire _2791 = r576 ^ r683;
  wire _2792 = _2790 ^ _2791;
  wire _2793 = r799 ^ r862;
  wire _2794 = r963 ^ r1046;
  wire _2795 = _2793 ^ _2794;
  wire _2796 = _2792 ^ _2795;
  wire _2797 = _2789 ^ _2796;
  wire _2798 = r1124 ^ r1206;
  wire _2799 = r1268 ^ r1426;
  wire _2800 = _2798 ^ _2799;
  wire _2801 = r1459 ^ r1544;
  wire _2802 = r1554 ^ r1731;
  wire _2803 = _2801 ^ _2802;
  wire _2804 = _2800 ^ _2803;
  wire _2805 = r1765 ^ r1832;
  wire _2806 = r1842 ^ r1853;
  wire _2807 = _2805 ^ _2806;
  wire _2808 = r1869 ^ r1917;
  wire _2809 = r2000 ^ r2005;
  wire _2810 = _2808 ^ _2809;
  wire _2811 = _2807 ^ _2810;
  wire _2812 = _2804 ^ _2811;
  wire _2813 = _2797 ^ _2812;
  wire _2814 = _2782 | _2813;
  wire _2815 = _2751 | _2814;
  wire _2816 = _2688 | _2815;
  wire _2817 = r30 ^ r79;
  wire _2818 = r156 ^ r204;
  wire _2819 = _2817 ^ _2818;
  wire _2820 = r263 ^ r297;
  wire _2821 = r377 ^ r434;
  wire _2822 = _2820 ^ _2821;
  wire _2823 = _2819 ^ _2822;
  wire _2824 = r484 ^ r616;
  wire _2825 = r695 ^ r759;
  wire _2826 = _2824 ^ _2825;
  wire _2827 = r813 ^ r873;
  wire _2828 = r917 ^ r958;
  wire _2829 = _2827 ^ _2828;
  wire _2830 = _2826 ^ _2829;
  wire _2831 = _2823 ^ _2830;
  wire _2832 = r1014 ^ r1150;
  wire _2833 = r1179 ^ r1227;
  wire _2834 = _2832 ^ _2833;
  wire _2835 = r1278 ^ r1315;
  wire _2836 = r1354 ^ r1399;
  wire _2837 = _2835 ^ _2836;
  wire _2838 = _2834 ^ _2837;
  wire _2839 = r1438 ^ r1700;
  wire _2840 = r1799 ^ r1903;
  wire _2841 = _2839 ^ _2840;
  wire _2842 = r1911 ^ r1929;
  wire _2843 = r2037 ^ r2040;
  wire _2844 = _2842 ^ _2843;
  wire _2845 = _2841 ^ _2844;
  wire _2846 = _2838 ^ _2845;
  wire _2847 = _2831 ^ _2846;
  wire _2848 = r29 ^ r102;
  wire _2849 = r140 ^ r184;
  wire _2850 = _2848 ^ _2849;
  wire _2851 = r247 ^ r355;
  wire _2852 = r438 ^ r491;
  wire _2853 = _2851 ^ _2852;
  wire _2854 = _2850 ^ _2853;
  wire _2855 = r519 ^ r575;
  wire _2856 = r664 ^ r704;
  wire _2857 = _2855 ^ _2856;
  wire _2858 = r752 ^ r884;
  wire _2859 = r1130 ^ r1167;
  wire _2860 = _2858 ^ _2859;
  wire _2861 = _2857 ^ _2860;
  wire _2862 = _2854 ^ _2861;
  wire _2863 = r1213 ^ r1293;
  wire _2864 = r1377 ^ r1421;
  wire _2865 = _2863 ^ _2864;
  wire _2866 = r1585 ^ r1643;
  wire _2867 = r1686 ^ r1725;
  wire _2868 = _2866 ^ _2867;
  wire _2869 = _2865 ^ _2868;
  wire _2870 = r1861 ^ r1892;
  wire _2871 = r1894 ^ r1918;
  wire _2872 = _2870 ^ _2871;
  wire _2873 = r1935 ^ r1972;
  wire _2874 = r2025 ^ r2033;
  wire _2875 = _2873 ^ _2874;
  wire _2876 = _2872 ^ _2875;
  wire _2877 = _2869 ^ _2876;
  wire _2878 = _2862 ^ _2877;
  wire _2879 = _2847 | _2878;
  wire _2880 = r28 ^ r85;
  wire _2881 = r168 ^ r175;
  wire _2882 = _2880 ^ _2881;
  wire _2883 = r258 ^ r307;
  wire _2884 = r358 ^ r447;
  wire _2885 = _2883 ^ _2884;
  wire _2886 = _2882 ^ _2885;
  wire _2887 = r459 ^ r527;
  wire _2888 = r661 ^ r756;
  wire _2889 = _2887 ^ _2888;
  wire _2890 = r783 ^ r904;
  wire _2891 = r952 ^ r1084;
  wire _2892 = _2890 ^ _2891;
  wire _2893 = _2889 ^ _2892;
  wire _2894 = _2886 ^ _2893;
  wire _2895 = r1142 ^ r1181;
  wire _2896 = r1291 ^ r1330;
  wire _2897 = _2895 ^ _2896;
  wire _2898 = r1383 ^ r1559;
  wire _2899 = r1630 ^ r1703;
  wire _2900 = _2898 ^ _2899;
  wire _2901 = _2897 ^ _2900;
  wire _2902 = r1834 ^ r1841;
  wire _2903 = r1846 ^ r1881;
  wire _2904 = _2902 ^ _2903;
  wire _2905 = r1882 ^ r1888;
  wire _2906 = r1923 ^ r1925;
  wire _2907 = _2905 ^ _2906;
  wire _2908 = _2904 ^ _2907;
  wire _2909 = _2901 ^ _2908;
  wire _2910 = _2894 ^ _2909;
  wire _2911 = r27 ^ r96;
  wire _2912 = r158 ^ r191;
  wire _2913 = _2911 ^ _2912;
  wire _2914 = r269 ^ r280;
  wire _2915 = r344 ^ r457;
  wire _2916 = _2914 ^ _2915;
  wire _2917 = _2913 ^ _2916;
  wire _2918 = r606 ^ r690;
  wire _2919 = r746 ^ r792;
  wire _2920 = _2918 ^ _2919;
  wire _2921 = r845 ^ r937;
  wire _2922 = r978 ^ r1007;
  wire _2923 = _2921 ^ _2922;
  wire _2924 = _2920 ^ _2923;
  wire _2925 = _2917 ^ _2924;
  wire _2926 = r1059 ^ r1151;
  wire _2927 = r1193 ^ r1256;
  wire _2928 = _2926 ^ _2927;
  wire _2929 = r1367 ^ r1384;
  wire _2930 = r1398 ^ r1591;
  wire _2931 = _2929 ^ _2930;
  wire _2932 = _2928 ^ _2931;
  wire _2933 = r1645 ^ r1733;
  wire _2934 = r1792 ^ r1905;
  wire _2935 = _2933 ^ _2934;
  wire _2936 = r1979 ^ r1999;
  wire _2937 = r2028 ^ r2034;
  wire _2938 = _2936 ^ _2937;
  wire _2939 = _2935 ^ _2938;
  wire _2940 = _2932 ^ _2939;
  wire _2941 = _2925 ^ _2940;
  wire _2942 = _2910 | _2941;
  wire _2943 = _2879 | _2942;
  wire _2944 = r26 ^ r103;
  wire _2945 = r145 ^ r195;
  wire _2946 = _2944 ^ _2945;
  wire _2947 = r242 ^ r324;
  wire _2948 = r378 ^ r432;
  wire _2949 = _2947 ^ _2948;
  wire _2950 = _2946 ^ _2949;
  wire _2951 = r489 ^ r516;
  wire _2952 = r613 ^ r646;
  wire _2953 = _2951 ^ _2952;
  wire _2954 = r718 ^ r726;
  wire _2955 = r786 ^ r831;
  wire _2956 = _2954 ^ _2955;
  wire _2957 = _2953 ^ _2956;
  wire _2958 = _2950 ^ _2957;
  wire _2959 = r887 ^ r906;
  wire _2960 = r984 ^ r1030;
  wire _2961 = _2959 ^ _2960;
  wire _2962 = r1070 ^ r1123;
  wire _2963 = r1191 ^ r1270;
  wire _2964 = _2962 ^ _2963;
  wire _2965 = _2961 ^ _2964;
  wire _2966 = r1298 ^ r1369;
  wire _2967 = r1385 ^ r1478;
  wire _2968 = _2966 ^ _2967;
  wire _2969 = r1613 ^ r1687;
  wire _2970 = r1697 ^ r1744;
  wire _2971 = _2969 ^ _2970;
  wire _2972 = _2968 ^ _2971;
  wire _2973 = _2965 ^ _2972;
  wire _2974 = _2958 ^ _2973;
  wire _2975 = r25 ^ r78;
  wire _2976 = r164 ^ r224;
  wire _2977 = _2975 ^ _2976;
  wire _2978 = r231 ^ r311;
  wire _2979 = r340 ^ r413;
  wire _2980 = _2978 ^ _2979;
  wire _2981 = _2977 ^ _2980;
  wire _2982 = r471 ^ r545;
  wire _2983 = r581 ^ r647;
  wire _2984 = _2982 ^ _2983;
  wire _2985 = r698 ^ r765;
  wire _2986 = r790 ^ r848;
  wire _2987 = _2985 ^ _2986;
  wire _2988 = _2984 ^ _2987;
  wire _2989 = _2981 ^ _2988;
  wire _2990 = r919 ^ r967;
  wire _2991 = r1013 ^ r1064;
  wire _2992 = _2990 ^ _2991;
  wire _2993 = r1138 ^ r1209;
  wire _2994 = r1219 ^ r1266;
  wire _2995 = _2993 ^ _2994;
  wire _2996 = _2992 ^ _2995;
  wire _2997 = r1327 ^ r1408;
  wire _2998 = r1456 ^ r1579;
  wire _2999 = _2997 ^ _2998;
  wire _3000 = r1622 ^ r1661;
  wire _3001 = r1715 ^ r1745;
  wire _3002 = _3000 ^ _3001;
  wire _3003 = _2999 ^ _3002;
  wire _3004 = _2996 ^ _3003;
  wire _3005 = _2989 ^ _3004;
  wire _3006 = _2974 | _3005;
  wire _3007 = r24 ^ r92;
  wire _3008 = r194 ^ r329;
  wire _3009 = _3007 ^ _3008;
  wire _3010 = r368 ^ r421;
  wire _3011 = r474 ^ r522;
  wire _3012 = _3010 ^ _3011;
  wire _3013 = _3009 ^ _3012;
  wire _3014 = r579 ^ r719;
  wire _3015 = r776 ^ r780;
  wire _3016 = _3014 ^ _3015;
  wire _3017 = r915 ^ r969;
  wire _3018 = r1024 ^ r1068;
  wire _3019 = _3017 ^ _3018;
  wire _3020 = _3016 ^ _3019;
  wire _3021 = _3013 ^ _3020;
  wire _3022 = r1164 ^ r1175;
  wire _3023 = r1230 ^ r1375;
  wire _3024 = _3022 ^ _3023;
  wire _3025 = r1412 ^ r1467;
  wire _3026 = r1482 ^ r1617;
  wire _3027 = _3025 ^ _3026;
  wire _3028 = _3024 ^ _3027;
  wire _3029 = r1656 ^ r1805;
  wire _3030 = r1887 ^ r1895;
  wire _3031 = _3029 ^ _3030;
  wire _3032 = r1901 ^ r1933;
  wire _3033 = r1936 ^ r1943;
  wire _3034 = _3032 ^ _3033;
  wire _3035 = _3031 ^ _3034;
  wire _3036 = _3028 ^ _3035;
  wire _3037 = _3021 ^ _3036;
  wire _3038 = r23 ^ r63;
  wire _3039 = r134 ^ r190;
  wire _3040 = _3038 ^ _3039;
  wire _3041 = r234 ^ r303;
  wire _3042 = r352 ^ r443;
  wire _3043 = _3041 ^ _3042;
  wire _3044 = _3040 ^ _3043;
  wire _3045 = r460 ^ r547;
  wire _3046 = r611 ^ r618;
  wire _3047 = _3045 ^ _3046;
  wire _3048 = r678 ^ r732;
  wire _3049 = r814 ^ r875;
  wire _3050 = _3048 ^ _3049;
  wire _3051 = _3047 ^ _3050;
  wire _3052 = _3044 ^ _3051;
  wire _3053 = r932 ^ r995;
  wire _3054 = r1031 ^ r1145;
  wire _3055 = _3053 ^ _3054;
  wire _3056 = r1176 ^ r1250;
  wire _3057 = r1444 ^ r1487;
  wire _3058 = _3056 ^ _3057;
  wire _3059 = _3055 ^ _3058;
  wire _3060 = r1507 ^ r1528;
  wire _3061 = r1535 ^ r1552;
  wire _3062 = _3060 ^ _3061;
  wire _3063 = r1566 ^ r1623;
  wire _3064 = r1684 ^ r1746;
  wire _3065 = _3063 ^ _3064;
  wire _3066 = _3062 ^ _3065;
  wire _3067 = _3059 ^ _3066;
  wire _3068 = _3052 ^ _3067;
  wire _3069 = _3037 | _3068;
  wire _3070 = _3006 | _3069;
  wire _3071 = _2943 | _3070;
  wire _3072 = _2816 | _3071;
  wire _3073 = _2561 | _3072;
  wire _3074 = r22 ^ r98;
  wire _3075 = r150 ^ r172;
  wire _3076 = _3074 ^ _3075;
  wire _3077 = r251 ^ r380;
  wire _3078 = r441 ^ r490;
  wire _3079 = _3077 ^ _3078;
  wire _3080 = _3076 ^ _3079;
  wire _3081 = r560 ^ r592;
  wire _3082 = r631 ^ r675;
  wire _3083 = _3081 ^ _3082;
  wire _3084 = r760 ^ r798;
  wire _3085 = r870 ^ r899;
  wire _3086 = _3084 ^ _3085;
  wire _3087 = _3083 ^ _3086;
  wire _3088 = _3080 ^ _3087;
  wire _3089 = r976 ^ r1006;
  wire _3090 = r1090 ^ r1208;
  wire _3091 = _3089 ^ _3090;
  wire _3092 = r1251 ^ r1283;
  wire _3093 = r1338 ^ r1453;
  wire _3094 = _3092 ^ _3093;
  wire _3095 = _3091 ^ _3094;
  wire _3096 = r1476 ^ r1513;
  wire _3097 = r1571 ^ r1612;
  wire _3098 = _3096 ^ _3097;
  wire _3099 = r1689 ^ r1735;
  wire _3100 = r1886 ^ r1908;
  wire _3101 = _3099 ^ _3100;
  wire _3102 = _3098 ^ _3101;
  wire _3103 = _3095 ^ _3102;
  wire _3104 = _3088 ^ _3103;
  wire _3105 = r21 ^ r65;
  wire _3106 = r142 ^ r180;
  wire _3107 = _3105 ^ _3106;
  wire _3108 = r260 ^ r316;
  wire _3109 = r370 ^ r419;
  wire _3110 = _3108 ^ _3109;
  wire _3111 = _3107 ^ _3110;
  wire _3112 = r456 ^ r557;
  wire _3113 = r595 ^ r636;
  wire _3114 = _3112 ^ _3113;
  wire _3115 = r693 ^ r748;
  wire _3116 = r809 ^ r876;
  wire _3117 = _3115 ^ _3116;
  wire _3118 = _3114 ^ _3117;
  wire _3119 = _3111 ^ _3118;
  wire _3120 = r900 ^ r988;
  wire _3121 = r1020 ^ r1077;
  wire _3122 = _3120 ^ _3121;
  wire _3123 = r1125 ^ r1199;
  wire _3124 = r1229 ^ r1324;
  wire _3125 = _3123 ^ _3124;
  wire _3126 = _3122 ^ _3125;
  wire _3127 = r1368 ^ r1406;
  wire _3128 = r1447 ^ r1575;
  wire _3129 = _3127 ^ _3128;
  wire _3130 = r1596 ^ r1633;
  wire _3131 = r1665 ^ r1747;
  wire _3132 = _3130 ^ _3131;
  wire _3133 = _3129 ^ _3132;
  wire _3134 = _3126 ^ _3133;
  wire _3135 = _3119 ^ _3134;
  wire _3136 = _3104 | _3135;
  wire _3137 = r20 ^ r116;
  wire _3138 = r199 ^ r255;
  wire _3139 = _3137 ^ _3138;
  wire _3140 = r308 ^ r356;
  wire _3141 = r400 ^ r482;
  wire _3142 = _3140 ^ _3141;
  wire _3143 = _3139 ^ _3142;
  wire _3144 = r518 ^ r582;
  wire _3145 = r668 ^ r714;
  wire _3146 = _3144 ^ _3145;
  wire _3147 = r735 ^ r820;
  wire _3148 = r866 ^ r931;
  wire _3149 = _3147 ^ _3148;
  wire _3150 = _3146 ^ _3149;
  wire _3151 = _3143 ^ _3150;
  wire _3152 = r996 ^ r1048;
  wire _3153 = r1215 ^ r1382;
  wire _3154 = _3152 ^ _3153;
  wire _3155 = r1450 ^ r1520;
  wire _3156 = r1551 ^ r1570;
  wire _3157 = _3155 ^ _3156;
  wire _3158 = _3154 ^ _3157;
  wire _3159 = r1584 ^ r1638;
  wire _3160 = r1699 ^ r1781;
  wire _3161 = _3159 ^ _3160;
  wire _3162 = r1818 ^ r1968;
  wire _3163 = r2036 ^ r2041;
  wire _3164 = _3162 ^ _3163;
  wire _3165 = _3161 ^ _3164;
  wire _3166 = _3158 ^ _3165;
  wire _3167 = _3151 ^ _3166;
  wire _3168 = r19 ^ r76;
  wire _3169 = r126 ^ r198;
  wire _3170 = _3168 ^ _3169;
  wire _3171 = r261 ^ r285;
  wire _3172 = r376 ^ r402;
  wire _3173 = _3171 ^ _3172;
  wire _3174 = _3170 ^ _3173;
  wire _3175 = r467 ^ r540;
  wire _3176 = r612 ^ r635;
  wire _3177 = _3175 ^ _3176;
  wire _3178 = r715 ^ r750;
  wire _3179 = r793 ^ r834;
  wire _3180 = _3178 ^ _3179;
  wire _3181 = _3177 ^ _3180;
  wire _3182 = _3174 ^ _3181;
  wire _3183 = r925 ^ r968;
  wire _3184 = r1026 ^ r1096;
  wire _3185 = _3183 ^ _3184;
  wire _3186 = r1140 ^ r1238;
  wire _3187 = r1290 ^ r1355;
  wire _3188 = _3186 ^ _3187;
  wire _3189 = _3185 ^ _3188;
  wire _3190 = r1395 ^ r1558;
  wire _3191 = r1564 ^ r1592;
  wire _3192 = _3190 ^ _3191;
  wire _3193 = r1626 ^ r1649;
  wire _3194 = r1691 ^ r1748;
  wire _3195 = _3193 ^ _3194;
  wire _3196 = _3192 ^ _3195;
  wire _3197 = _3189 ^ _3196;
  wire _3198 = _3182 ^ _3197;
  wire _3199 = _3167 | _3198;
  wire _3200 = _3136 | _3199;
  wire _3201 = r18 ^ r94;
  wire _3202 = r120 ^ r178;
  wire _3203 = _3201 ^ _3202;
  wire _3204 = r250 ^ r295;
  wire _3205 = r349 ^ r444;
  wire _3206 = _3204 ^ _3205;
  wire _3207 = _3203 ^ _3206;
  wire _3208 = r492 ^ r541;
  wire _3209 = r578 ^ r692;
  wire _3210 = _3208 ^ _3209;
  wire _3211 = r770 ^ r782;
  wire _3212 = r840 ^ r941;
  wire _3213 = _3211 ^ _3212;
  wire _3214 = _3210 ^ _3213;
  wire _3215 = _3207 ^ _3214;
  wire _3216 = r983 ^ r1050;
  wire _3217 = r1071 ^ r1163;
  wire _3218 = _3216 ^ _3217;
  wire _3219 = r1220 ^ r1241;
  wire _3220 = r1301 ^ r1335;
  wire _3221 = _3219 ^ _3220;
  wire _3222 = _3218 ^ _3221;
  wire _3223 = r1417 ^ r1441;
  wire _3224 = r1519 ^ r1602;
  wire _3225 = _3223 ^ _3224;
  wire _3226 = r1627 ^ r1671;
  wire _3227 = r1778 ^ r1825;
  wire _3228 = _3226 ^ _3227;
  wire _3229 = _3225 ^ _3228;
  wire _3230 = _3222 ^ _3229;
  wire _3231 = _3215 ^ _3230;
  wire _3232 = r17 ^ r58;
  wire _3233 = r123 ^ r211;
  wire _3234 = _3232 ^ _3233;
  wire _3235 = r273 ^ r289;
  wire _3236 = r346 ^ r420;
  wire _3237 = _3235 ^ _3236;
  wire _3238 = _3234 ^ _3237;
  wire _3239 = r517 ^ r603;
  wire _3240 = r684 ^ r724;
  wire _3241 = _3239 ^ _3240;
  wire _3242 = r823 ^ r830;
  wire _3243 = r879 ^ r889;
  wire _3244 = _3242 ^ _3243;
  wire _3245 = _3241 ^ _3244;
  wire _3246 = _3238 ^ _3245;
  wire _3247 = r954 ^ r1357;
  wire _3248 = r1472 ^ r1488;
  wire _3249 = _3247 ^ _3248;
  wire _3250 = r1508 ^ r1516;
  wire _3251 = r1525 ^ r1674;
  wire _3252 = _3250 ^ _3251;
  wire _3253 = _3249 ^ _3252;
  wire _3254 = r1710 ^ r1831;
  wire _3255 = r1840 ^ r1850;
  wire _3256 = _3254 ^ _3255;
  wire _3257 = r1884 ^ r1912;
  wire _3258 = r1997 ^ r2002;
  wire _3259 = _3257 ^ _3258;
  wire _3260 = _3256 ^ _3259;
  wire _3261 = _3253 ^ _3260;
  wire _3262 = _3246 ^ _3261;
  wire _3263 = _3231 | _3262;
  wire _3264 = r16 ^ r59;
  wire _3265 = r113 ^ r214;
  wire _3266 = _3264 ^ _3265;
  wire _3267 = r226 ^ r361;
  wire _3268 = r440 ^ r472;
  wire _3269 = _3267 ^ _3268;
  wire _3270 = _3266 ^ _3269;
  wire _3271 = r510 ^ r589;
  wire _3272 = r621 ^ r702;
  wire _3273 = _3271 ^ _3272;
  wire _3274 = r774 ^ r881;
  wire _3275 = r991 ^ r1005;
  wire _3276 = _3274 ^ _3275;
  wire _3277 = _3273 ^ _3276;
  wire _3278 = _3270 ^ _3277;
  wire _3279 = r1098 ^ r1139;
  wire _3280 = r1285 ^ r1477;
  wire _3281 = _3279 ^ _3280;
  wire _3282 = r1502 ^ r1631;
  wire _3283 = r1666 ^ r1713;
  wire _3284 = _3282 ^ _3283;
  wire _3285 = _3281 ^ _3284;
  wire _3286 = r1798 ^ r1844;
  wire _3287 = r1890 ^ r1906;
  wire _3288 = _3286 ^ _3287;
  wire _3289 = r1989 ^ r2004;
  wire _3290 = r2023 ^ r2027;
  wire _3291 = _3289 ^ _3290;
  wire _3292 = _3288 ^ _3291;
  wire _3293 = _3285 ^ _3292;
  wire _3294 = _3278 ^ _3293;
  wire _3295 = r15 ^ r93;
  wire _3296 = r151 ^ r200;
  wire _3297 = _3295 ^ _3296;
  wire _3298 = r265 ^ r284;
  wire _3299 = r354 ^ r410;
  wire _3300 = _3298 ^ _3299;
  wire _3301 = _3297 ^ _3300;
  wire _3302 = r488 ^ r525;
  wire _3303 = r614 ^ r642;
  wire _3304 = _3302 ^ _3303;
  wire _3305 = r706 ^ r802;
  wire _3306 = r852 ^ r888;
  wire _3307 = _3305 ^ _3306;
  wire _3308 = _3304 ^ _3307;
  wire _3309 = _3301 ^ _3308;
  wire _3310 = r956 ^ r1022;
  wire _3311 = r1062 ^ r1131;
  wire _3312 = _3310 ^ _3311;
  wire _3313 = r1197 ^ r1236;
  wire _3314 = r1326 ^ r1366;
  wire _3315 = _3313 ^ _3314;
  wire _3316 = _3312 ^ _3315;
  wire _3317 = r1538 ^ r1553;
  wire _3318 = r1573 ^ r1604;
  wire _3319 = _3317 ^ _3318;
  wire _3320 = r1642 ^ r1650;
  wire _3321 = r1712 ^ r1749;
  wire _3322 = _3320 ^ _3321;
  wire _3323 = _3319 ^ _3322;
  wire _3324 = _3316 ^ _3323;
  wire _3325 = _3309 ^ _3324;
  wire _3326 = _3294 | _3325;
  wire _3327 = _3263 | _3326;
  wire _3328 = _3200 | _3327;
  wire _3329 = r14 ^ r86;
  wire _3330 = r133 ^ r179;
  wire _3331 = _3329 ^ _3330;
  wire _3332 = r267 ^ r317;
  wire _3333 = r388 ^ r396;
  wire _3334 = _3332 ^ _3333;
  wire _3335 = _3331 ^ _3334;
  wire _3336 = r464 ^ r530;
  wire _3337 = r605 ^ r640;
  wire _3338 = _3336 ^ _3337;
  wire _3339 = r769 ^ r811;
  wire _3340 = r832 ^ r939;
  wire _3341 = _3339 ^ _3340;
  wire _3342 = _3338 ^ _3341;
  wire _3343 = _3335 ^ _3342;
  wire _3344 = r970 ^ r1043;
  wire _3345 = r1080 ^ r1149;
  wire _3346 = _3344 ^ _3345;
  wire _3347 = r1204 ^ r1274;
  wire _3348 = r1312 ^ r1454;
  wire _3349 = _3347 ^ _3348;
  wire _3350 = _3346 ^ _3349;
  wire _3351 = r1470 ^ r1480;
  wire _3352 = r1489 ^ r1498;
  wire _3353 = _3351 ^ _3352;
  wire _3354 = r1533 ^ r1663;
  wire _3355 = r1714 ^ r1750;
  wire _3356 = _3354 ^ _3355;
  wire _3357 = _3353 ^ _3356;
  wire _3358 = _3350 ^ _3357;
  wire _3359 = _3343 ^ _3358;
  wire _3360 = r13 ^ r146;
  wire _3361 = r197 ^ r237;
  wire _3362 = _3360 ^ _3361;
  wire _3363 = r300 ^ r338;
  wire _3364 = r422 ^ r462;
  wire _3365 = _3363 ^ _3364;
  wire _3366 = _3362 ^ _3365;
  wire _3367 = r593 ^ r705;
  wire _3368 = r737 ^ r806;
  wire _3369 = _3367 ^ _3368;
  wire _3370 = r844 ^ r922;
  wire _3371 = r966 ^ r1044;
  wire _3372 = _3370 ^ _3371;
  wire _3373 = _3369 ^ _3372;
  wire _3374 = _3366 ^ _3373;
  wire _3375 = r1089 ^ r1172;
  wire _3376 = r1225 ^ r1351;
  wire _3377 = _3375 ^ _3376;
  wire _3378 = r1418 ^ r1428;
  wire _3379 = r1443 ^ r1497;
  wire _3380 = _3378 ^ _3379;
  wire _3381 = _3377 ^ _3380;
  wire _3382 = r1526 ^ r1709;
  wire _3383 = r1783 ^ r1806;
  wire _3384 = _3382 ^ _3383;
  wire _3385 = r1966 ^ r2012;
  wire _3386 = r2044 ^ r2046;
  wire _3387 = _3385 ^ _3386;
  wire _3388 = _3384 ^ _3387;
  wire _3389 = _3381 ^ _3388;
  wire _3390 = _3374 ^ _3389;
  wire _3391 = _3359 | _3390;
  wire _3392 = r12 ^ r157;
  wire _3393 = r223 ^ r272;
  wire _3394 = _3392 ^ _3393;
  wire _3395 = r312 ^ r333;
  wire _3396 = r412 ^ r529;
  wire _3397 = _3395 ^ _3396;
  wire _3398 = _3394 ^ _3397;
  wire _3399 = r610 ^ r700;
  wire _3400 = r744 ^ r812;
  wire _3401 = _3399 ^ _3400;
  wire _3402 = r853 ^ r929;
  wire _3403 = r986 ^ r1021;
  wire _3404 = _3402 ^ _3403;
  wire _3405 = _3401 ^ _3404;
  wire _3406 = _3398 ^ _3405;
  wire _3407 = r1085 ^ r1170;
  wire _3408 = r1246 ^ r1280;
  wire _3409 = _3407 ^ _3408;
  wire _3410 = r1295 ^ r1352;
  wire _3411 = r1394 ^ r1514;
  wire _3412 = _3410 ^ _3411;
  wire _3413 = _3409 ^ _3412;
  wire _3414 = r1594 ^ r1637;
  wire _3415 = r1803 ^ r1807;
  wire _3416 = _3414 ^ _3415;
  wire _3417 = r1885 ^ r1938;
  wire _3418 = r1953 ^ r1963;
  wire _3419 = _3417 ^ _3418;
  wire _3420 = _3416 ^ _3419;
  wire _3421 = _3413 ^ _3420;
  wire _3422 = _3406 ^ _3421;
  wire _3423 = r110 ^ r127;
  wire _3424 = r207 ^ r230;
  wire _3425 = _3423 ^ _3424;
  wire _3426 = r323 ^ r335;
  wire _3427 = r469 ^ r586;
  wire _3428 = _3426 ^ _3427;
  wire _3429 = _3425 ^ _3428;
  wire _3430 = r656 ^ r681;
  wire _3431 = r728 ^ r801;
  wire _3432 = _3430 ^ _3431;
  wire _3433 = r880 ^ r895;
  wire _3434 = r949 ^ r1153;
  wire _3435 = _3433 ^ _3434;
  wire _3436 = _3432 ^ _3435;
  wire _3437 = _3429 ^ _3436;
  wire _3438 = r1202 ^ r1244;
  wire _3439 = r1302 ^ r1333;
  wire _3440 = _3438 ^ _3439;
  wire _3441 = r1415 ^ r1445;
  wire _3442 = r1729 ^ r1793;
  wire _3443 = _3441 ^ _3442;
  wire _3444 = _3440 ^ _3443;
  wire _3445 = r1797 ^ r1817;
  wire _3446 = r1835 ^ r1889;
  wire _3447 = _3445 ^ _3446;
  wire _3448 = r1977 ^ r1981;
  wire _3449 = r2045 ^ r2047;
  wire _3450 = _3448 ^ _3449;
  wire _3451 = _3447 ^ _3450;
  wire _3452 = _3444 ^ _3451;
  wire _3453 = _3437 ^ _3452;
  wire _3454 = _3422 | _3453;
  wire _3455 = _3391 | _3454;
  wire _3456 = r11 ^ r105;
  wire _3457 = r115 ^ r181;
  wire _3458 = _3456 ^ _3457;
  wire _3459 = r238 ^ r296;
  wire _3460 = r385 ^ r418;
  wire _3461 = _3459 ^ _3460;
  wire _3462 = _3458 ^ _3461;
  wire _3463 = r500 ^ r508;
  wire _3464 = r583 ^ r643;
  wire _3465 = _3463 ^ _3464;
  wire _3466 = r689 ^ r730;
  wire _3467 = r826 ^ r839;
  wire _3468 = _3466 ^ _3467;
  wire _3469 = _3465 ^ _3468;
  wire _3470 = _3462 ^ _3469;
  wire _3471 = r893 ^ r950;
  wire _3472 = r1029 ^ r1108;
  wire _3473 = _3471 ^ _3472;
  wire _3474 = r1147 ^ r1184;
  wire _3475 = r1299 ^ r1376;
  wire _3476 = _3474 ^ _3475;
  wire _3477 = _3473 ^ _3476;
  wire _3478 = r1471 ^ r1523;
  wire _3479 = r1548 ^ r1595;
  wire _3480 = _3478 ^ _3479;
  wire _3481 = r1644 ^ r1683;
  wire _3482 = r1717 ^ r1751;
  wire _3483 = _3481 ^ _3482;
  wire _3484 = _3480 ^ _3483;
  wire _3485 = _3477 ^ _3484;
  wire _3486 = _3470 ^ _3485;
  wire _3487 = r10 ^ r100;
  wire _3488 = r160 ^ r171;
  wire _3489 = _3487 ^ _3488;
  wire _3490 = r266 ^ r362;
  wire _3491 = r454 ^ r598;
  wire _3492 = _3490 ^ _3491;
  wire _3493 = _3489 ^ _3492;
  wire _3494 = r711 ^ r754;
  wire _3495 = r778 ^ r927;
  wire _3496 = _3494 ^ _3495;
  wire _3497 = r985 ^ r1129;
  wire _3498 = r1169 ^ r1186;
  wire _3499 = _3497 ^ _3498;
  wire _3500 = _3496 ^ _3499;
  wire _3501 = _3493 ^ _3500;
  wire _3502 = r1258 ^ r1303;
  wire _3503 = r1337 ^ r1588;
  wire _3504 = _3502 ^ _3503;
  wire _3505 = r1615 ^ r1672;
  wire _3506 = r1732 ^ r1734;
  wire _3507 = _3505 ^ _3506;
  wire _3508 = _3504 ^ _3507;
  wire _3509 = r1767 ^ r1858;
  wire _3510 = r1893 ^ r1927;
  wire _3511 = _3509 ^ _3510;
  wire _3512 = r1939 ^ r2007;
  wire _3513 = r2029 ^ r2042;
  wire _3514 = _3512 ^ _3513;
  wire _3515 = _3511 ^ _3514;
  wire _3516 = _3508 ^ _3515;
  wire _3517 = _3501 ^ _3516;
  wire _3518 = _3486 | _3517;
  wire _3519 = r9 ^ r83;
  wire _3520 = r118 ^ r212;
  wire _3521 = _3519 ^ _3520;
  wire _3522 = r225 ^ r326;
  wire _3523 = r345 ^ r446;
  wire _3524 = _3522 ^ _3523;
  wire _3525 = _3521 ^ _3524;
  wire _3526 = r504 ^ r536;
  wire _3527 = r591 ^ r639;
  wire _3528 = _3526 ^ _3527;
  wire _3529 = r710 ^ r736;
  wire _3530 = r816 ^ r847;
  wire _3531 = _3529 ^ _3530;
  wire _3532 = _3528 ^ _3531;
  wire _3533 = _3525 ^ _3532;
  wire _3534 = r909 ^ r977;
  wire _3535 = r1107 ^ r1136;
  wire _3536 = _3534 ^ _3535;
  wire _3537 = r1165 ^ r1173;
  wire _3538 = r1261 ^ r1294;
  wire _3539 = _3537 ^ _3538;
  wire _3540 = _3536 ^ _3539;
  wire _3541 = r1341 ^ r1439;
  wire _3542 = r1458 ^ r1494;
  wire _3543 = _3541 ^ _3542;
  wire _3544 = r1505 ^ r1628;
  wire _3545 = r1704 ^ r1752;
  wire _3546 = _3544 ^ _3545;
  wire _3547 = _3543 ^ _3546;
  wire _3548 = _3540 ^ _3547;
  wire _3549 = _3533 ^ _3548;
  wire _3550 = r8 ^ r90;
  wire _3551 = r138 ^ r177;
  wire _3552 = _3550 ^ _3551;
  wire _3553 = r252 ^ r287;
  wire _3554 = r357 ^ r405;
  wire _3555 = _3553 ^ _3554;
  wire _3556 = _3552 ^ _3555;
  wire _3557 = r451 ^ r534;
  wire _3558 = r567 ^ r665;
  wire _3559 = _3557 ^ _3558;
  wire _3560 = r687 ^ r747;
  wire _3561 = r818 ^ r868;
  wire _3562 = _3560 ^ _3561;
  wire _3563 = _3559 ^ _3562;
  wire _3564 = _3556 ^ _3563;
  wire _3565 = r911 ^ r994;
  wire _3566 = r1033 ^ r1092;
  wire _3567 = _3565 ^ _3566;
  wire _3568 = r1159 ^ r1203;
  wire _3569 = r1218 ^ r1247;
  wire _3570 = _3568 ^ _3569;
  wire _3571 = _3567 ^ _3570;
  wire _3572 = r1314 ^ r1390;
  wire _3573 = r1465 ^ r1536;
  wire _3574 = _3572 ^ _3573;
  wire _3575 = r1550 ^ r1668;
  wire _3576 = r1782 ^ r1826;
  wire _3577 = _3575 ^ _3576;
  wire _3578 = _3574 ^ _3577;
  wire _3579 = _3571 ^ _3578;
  wire _3580 = _3564 ^ _3579;
  wire _3581 = _3549 | _3580;
  wire _3582 = _3518 | _3581;
  wire _3583 = _3455 | _3582;
  wire _3584 = _3328 | _3583;
  wire _3585 = r7 ^ r54;
  wire _3586 = r148 ^ r205;
  wire _3587 = _3585 ^ _3586;
  wire _3588 = r233 ^ r305;
  wire _3589 = r369 ^ r398;
  wire _3590 = _3588 ^ _3589;
  wire _3591 = _3587 ^ _3590;
  wire _3592 = r497 ^ r513;
  wire _3593 = r577 ^ r652;
  wire _3594 = _3592 ^ _3593;
  wire _3595 = r669 ^ r755;
  wire _3596 = r788 ^ r882;
  wire _3597 = _3595 ^ _3596;
  wire _3598 = _3594 ^ _3597;
  wire _3599 = _3591 ^ _3598;
  wire _3600 = r896 ^ r999;
  wire _3601 = r1028 ^ r1060;
  wire _3602 = _3600 ^ _3601;
  wire _3603 = r1094 ^ r1157;
  wire _3604 = r1321 ^ r1340;
  wire _3605 = _3603 ^ _3604;
  wire _3606 = _3602 ^ _3605;
  wire _3607 = r1473 ^ r1518;
  wire _3608 = r1524 ^ r1598;
  wire _3609 = _3607 ^ _3608;
  wire _3610 = r1640 ^ r1667;
  wire _3611 = r1698 ^ r1753;
  wire _3612 = _3610 ^ _3611;
  wire _3613 = _3609 ^ _3612;
  wire _3614 = _3606 ^ _3613;
  wire _3615 = _3599 ^ _3614;
  wire _3616 = r6 ^ r108;
  wire _3617 = r143 ^ r202;
  wire _3618 = _3616 ^ _3617;
  wire _3619 = r253 ^ r314;
  wire _3620 = r339 ^ r429;
  wire _3621 = _3619 ^ _3620;
  wire _3622 = _3618 ^ _3621;
  wire _3623 = r550 ^ r570;
  wire _3624 = r622 ^ r671;
  wire _3625 = _3623 ^ _3624;
  wire _3626 = r729 ^ r824;
  wire _3627 = r878 ^ r928;
  wire _3628 = _3626 ^ _3627;
  wire _3629 = _3625 ^ _3628;
  wire _3630 = _3622 ^ _3629;
  wire _3631 = r1011 ^ r1066;
  wire _3632 = r1134 ^ r1194;
  wire _3633 = _3631 ^ _3632;
  wire _3634 = r1243 ^ r1305;
  wire _3635 = r1329 ^ r1393;
  wire _3636 = _3634 ^ _3635;
  wire _3637 = _3633 ^ _3636;
  wire _3638 = r1440 ^ r1503;
  wire _3639 = r1610 ^ r1677;
  wire _3640 = _3638 ^ _3639;
  wire _3641 = r1728 ^ r1737;
  wire _3642 = r1794 ^ r1827;
  wire _3643 = _3641 ^ _3642;
  wire _3644 = _3640 ^ _3643;
  wire _3645 = _3637 ^ _3644;
  wire _3646 = _3630 ^ _3645;
  wire _3647 = _3615 | _3646;
  wire _3648 = r5 ^ r88;
  wire _3649 = r149 ^ r216;
  wire _3650 = _3648 ^ _3649;
  wire _3651 = r268 ^ r309;
  wire _3652 = r387 ^ r439;
  wire _3653 = _3651 ^ _3652;
  wire _3654 = _3650 ^ _3653;
  wire _3655 = r461 ^ r553;
  wire _3656 = r574 ^ r667;
  wire _3657 = _3655 ^ _3656;
  wire _3658 = r712 ^ r743;
  wire _3659 = r781 ^ r842;
  wire _3660 = _3658 ^ _3659;
  wire _3661 = _3657 ^ _3660;
  wire _3662 = _3654 ^ _3661;
  wire _3663 = r892 ^ r998;
  wire _3664 = r1018 ^ r1099;
  wire _3665 = _3663 ^ _3664;
  wire _3666 = r1180 ^ r1271;
  wire _3667 = r1307 ^ r1373;
  wire _3668 = _3666 ^ _3667;
  wire _3669 = _3665 ^ _3668;
  wire _3670 = r1422 ^ r1429;
  wire _3671 = r1486 ^ r1555;
  wire _3672 = _3670 ^ _3671;
  wire _3673 = r1611 ^ r1736;
  wire _3674 = r1809 ^ r1828;
  wire _3675 = _3673 ^ _3674;
  wire _3676 = _3672 ^ _3675;
  wire _3677 = _3669 ^ _3676;
  wire _3678 = _3662 ^ _3677;
  wire _3679 = r4 ^ r68;
  wire _3680 = r137 ^ r209;
  wire _3681 = _3679 ^ _3680;
  wire _3682 = r264 ^ r315;
  wire _3683 = r372 ^ r433;
  wire _3684 = _3682 ^ _3683;
  wire _3685 = _3681 ^ _3684;
  wire _3686 = r473 ^ r537;
  wire _3687 = r564 ^ r654;
  wire _3688 = _3686 ^ _3687;
  wire _3689 = r688 ^ r771;
  wire _3690 = r789 ^ r864;
  wire _3691 = _3689 ^ _3690;
  wire _3692 = _3688 ^ _3691;
  wire _3693 = _3685 ^ _3692;
  wire _3694 = r920 ^ r992;
  wire _3695 = r1039 ^ r1111;
  wire _3696 = _3694 ^ _3695;
  wire _3697 = r1117 ^ r1205;
  wire _3698 = r1222 ^ r1255;
  wire _3699 = _3697 ^ _3698;
  wire _3700 = _3696 ^ _3699;
  wire _3701 = r1380 ^ r1420;
  wire _3702 = r1469 ^ r1530;
  wire _3703 = _3701 ^ _3702;
  wire _3704 = r1605 ^ r1639;
  wire _3705 = r1654 ^ r1754;
  wire _3706 = _3704 ^ _3705;
  wire _3707 = _3703 ^ _3706;
  wire _3708 = _3700 ^ _3707;
  wire _3709 = _3693 ^ _3708;
  wire _3710 = _3678 | _3709;
  wire _3711 = _3647 | _3710;
  wire _3712 = r71 ^ r163;
  wire _3713 = r187 ^ r228;
  wire _3714 = _3712 ^ _3713;
  wire _3715 = r304 ^ r390;
  wire _3716 = r437 ^ r483;
  wire _3717 = _3715 ^ _3716;
  wire _3718 = _3714 ^ _3717;
  wire _3719 = r514 ^ r599;
  wire _3720 = r620 ^ r709;
  wire _3721 = _3719 ^ _3720;
  wire _3722 = r749 ^ r817;
  wire _3723 = r905 ^ r974;
  wire _3724 = _3722 ^ _3723;
  wire _3725 = _3721 ^ _3724;
  wire _3726 = _3718 ^ _3725;
  wire _3727 = r1037 ^ r1067;
  wire _3728 = r1160 ^ r1196;
  wire _3729 = _3727 ^ _3728;
  wire _3730 = r1224 ^ r1226;
  wire _3731 = r1347 ^ r1386;
  wire _3732 = _3730 ^ _3731;
  wire _3733 = _3729 ^ _3732;
  wire _3734 = r1542 ^ r1632;
  wire _3735 = r1662 ^ r1785;
  wire _3736 = _3734 ^ _3735;
  wire _3737 = r1947 ^ r1998;
  wire _3738 = r2024 ^ r2035;
  wire _3739 = _3737 ^ _3738;
  wire _3740 = _3736 ^ _3739;
  wire _3741 = _3733 ^ _3740;
  wire _3742 = _3726 ^ _3741;
  wire _3743 = r3 ^ r55;
  wire _3744 = r111 ^ r196;
  wire _3745 = _3743 ^ _3744;
  wire _3746 = r426 ^ r455;
  wire _3747 = r533 ^ r648;
  wire _3748 = _3746 ^ _3747;
  wire _3749 = _3745 ^ _3748;
  wire _3750 = r679 ^ r841;
  wire _3751 = r930 ^ r981;
  wire _3752 = _3750 ^ _3751;
  wire _3753 = r1016 ^ r1093;
  wire _3754 = r1135 ^ r1185;
  wire _3755 = _3753 ^ _3754;
  wire _3756 = _3752 ^ _3755;
  wire _3757 = _3749 ^ _3756;
  wire _3758 = r1273 ^ r1325;
  wire _3759 = r1345 ^ r1449;
  wire _3760 = _3758 ^ _3759;
  wire _3761 = r1537 ^ r1576;
  wire _3762 = r1657 ^ r1701;
  wire _3763 = _3761 ^ _3762;
  wire _3764 = _3760 ^ _3763;
  wire _3765 = r1808 ^ r1864;
  wire _3766 = r1877 ^ r1913;
  wire _3767 = _3765 ^ _3766;
  wire _3768 = r1931 ^ r1934;
  wire _3769 = r1965 ^ r1974;
  wire _3770 = _3768 ^ _3769;
  wire _3771 = _3767 ^ _3770;
  wire _3772 = _3764 ^ _3771;
  wire _3773 = _3757 ^ _3772;
  wire _3774 = _3742 | _3773;
  wire _3775 = r2 ^ r89;
  wire _3776 = r152 ^ r249;
  wire _3777 = _3775 ^ _3776;
  wire _3778 = r282 ^ r359;
  wire _3779 = r406 ^ r499;
  wire _3780 = _3778 ^ _3779;
  wire _3781 = _3777 ^ _3780;
  wire _3782 = r506 ^ r594;
  wire _3783 = r645 ^ r803;
  wire _3784 = _3782 ^ _3783;
  wire _3785 = r833 ^ r945;
  wire _3786 = r1053 ^ r1106;
  wire _3787 = _3785 ^ _3786;
  wire _3788 = _3784 ^ _3787;
  wire _3789 = _3781 ^ _3788;
  wire _3790 = r1156 ^ r1201;
  wire _3791 = r1259 ^ r1281;
  wire _3792 = _3790 ^ _3791;
  wire _3793 = r1378 ^ r1403;
  wire _3794 = r1433 ^ r1492;
  wire _3795 = _3793 ^ _3794;
  wire _3796 = _3792 ^ _3795;
  wire _3797 = r1531 ^ r1599;
  wire _3798 = r1660 ^ r1711;
  wire _3799 = _3797 ^ _3798;
  wire _3800 = r1873 ^ r1924;
  wire _3801 = r1984 ^ r1985;
  wire _3802 = _3800 ^ _3801;
  wire _3803 = _3799 ^ _3802;
  wire _3804 = _3796 ^ _3803;
  wire _3805 = _3789 ^ _3804;
  wire _3806 = r1 ^ r107;
  wire _3807 = r154 ^ r227;
  wire _3808 = _3806 ^ _3807;
  wire _3809 = r319 ^ r445;
  wire _3810 = r546 ^ r604;
  wire _3811 = _3809 ^ _3810;
  wire _3812 = _3808 ^ _3811;
  wire _3813 = r659 ^ r727;
  wire _3814 = r784 ^ r851;
  wire _3815 = _3813 ^ _3814;
  wire _3816 = r1002 ^ r1056;
  wire _3817 = r1081 ^ r1126;
  wire _3818 = _3816 ^ _3817;
  wire _3819 = _3815 ^ _3818;
  wire _3820 = _3812 ^ _3819;
  wire _3821 = r1306 ^ r1359;
  wire _3822 = r1413 ^ r1427;
  wire _3823 = _3821 ^ _3822;
  wire _3824 = r1464 ^ r1522;
  wire _3825 = r1648 ^ r1688;
  wire _3826 = _3824 ^ _3825;
  wire _3827 = _3823 ^ _3826;
  wire _3828 = r1800 ^ r1879;
  wire _3829 = r1941 ^ r1942;
  wire _3830 = _3828 ^ _3829;
  wire _3831 = r1945 ^ r1955;
  wire _3832 = r1969 ^ r1975;
  wire _3833 = _3831 ^ _3832;
  wire _3834 = _3830 ^ _3833;
  wire _3835 = _3827 ^ _3834;
  wire _3836 = _3820 ^ _3835;
  wire _3837 = _3805 | _3836;
  wire _3838 = _3774 | _3837;
  wire _3839 = _3711 | _3838;
  wire _3840 = r0 ^ r80;
  wire _3841 = r321 ^ r360;
  wire _3842 = _3840 ^ _3841;
  wire _3843 = r401 ^ r502;
  wire _3844 = r515 ^ r653;
  wire _3845 = _3843 ^ _3844;
  wire _3846 = _3842 ^ _3845;
  wire _3847 = r745 ^ r805;
  wire _3848 = r855 ^ r980;
  wire _3849 = _3847 ^ _3848;
  wire _3850 = r1040 ^ r1061;
  wire _3851 = r1252 ^ r1320;
  wire _3852 = _3850 ^ _3851;
  wire _3853 = _3849 ^ _3852;
  wire _3854 = _3846 ^ _3853;
  wire _3855 = r1362 ^ r1407;
  wire _3856 = r1491 ^ r1562;
  wire _3857 = _3855 ^ _3856;
  wire _3858 = r1589 ^ r1716;
  wire _3859 = r1726 ^ r1780;
  wire _3860 = _3858 ^ _3859;
  wire _3861 = _3857 ^ _3860;
  wire _3862 = r1790 ^ r1852;
  wire _3863 = r1862 ^ r1899;
  wire _3864 = _3862 ^ _3863;
  wire _3865 = r1904 ^ r1958;
  wire _3866 = r2006 ^ r2009;
  wire _3867 = _3865 ^ _3866;
  wire _3868 = _3864 ^ _3867;
  wire _3869 = _3861 ^ _3868;
  wire _3870 = _3854 ^ _3869;
  wire _3871 = r64 ^ r161;
  wire _3872 = r217 ^ r236;
  wire _3873 = _3871 ^ _3872;
  wire _3874 = r291 ^ r350;
  wire _3875 = r411 ^ r466;
  wire _3876 = _3874 ^ _3875;
  wire _3877 = _3873 ^ _3876;
  wire _3878 = r566 ^ r628;
  wire _3879 = r670 ^ r767;
  wire _3880 = _3878 ^ _3879;
  wire _3881 = r819 ^ r901;
  wire _3882 = r959 ^ r1017;
  wire _3883 = _3881 ^ _3882;
  wire _3884 = _3880 ^ _3883;
  wire _3885 = _3877 ^ _3884;
  wire _3886 = r1083 ^ r1137;
  wire _3887 = r1189 ^ r1223;
  wire _3888 = _3886 ^ _3887;
  wire _3889 = r1249 ^ r1296;
  wire _3890 = r1348 ^ r1411;
  wire _3891 = _3889 ^ _3890;
  wire _3892 = _3888 ^ _3891;
  wire _3893 = r1479 ^ r1501;
  wire _3894 = r1572 ^ r1646;
  wire _3895 = _3893 ^ _3894;
  wire _3896 = r1696 ^ r1723;
  wire _3897 = r1766 ^ r1829;
  wire _3898 = _3896 ^ _3897;
  wire _3899 = _3895 ^ _3898;
  wire _3900 = _3892 ^ _3899;
  wire _3901 = _3885 ^ _3900;
  wire _3902 = _3870 | _3901;
  wire _3903 = r91 ^ r114;
  wire _3904 = r201 ^ r241;
  wire _3905 = _3903 ^ _3904;
  wire _3906 = r327 ^ r375;
  wire _3907 = r475 ^ r551;
  wire _3908 = _3906 ^ _3907;
  wire _3909 = _3905 ^ _3908;
  wire _3910 = r607 ^ r637;
  wire _3911 = r686 ^ r768;
  wire _3912 = _3910 ^ _3911;
  wire _3913 = r815 ^ r898;
  wire _3914 = r962 ^ r1036;
  wire _3915 = _3913 ^ _3914;
  wire _3916 = _3912 ^ _3915;
  wire _3917 = _3909 ^ _3916;
  wire _3918 = r1128 ^ r1182;
  wire _3919 = r1264 ^ r1328;
  wire _3920 = _3918 ^ _3919;
  wire _3921 = r1379 ^ r1400;
  wire _3922 = r1565 ^ r1673;
  wire _3923 = _3921 ^ _3922;
  wire _3924 = _3920 ^ _3923;
  wire _3925 = r1760 ^ r1771;
  wire _3926 = r1774 ^ r1789;
  wire _3927 = _3925 ^ _3926;
  wire _3928 = r1865 ^ r1928;
  wire _3929 = r1990 ^ r1991;
  wire _3930 = _3928 ^ _3929;
  wire _3931 = _3927 ^ _3930;
  wire _3932 = _3924 ^ _3931;
  wire _3933 = _3917 ^ _3932;
  wire _3934 = r82 ^ r122;
  wire _3935 = r213 ^ r279;
  wire _3936 = _3934 ^ _3935;
  wire _3937 = r382 ^ r428;
  wire _3938 = r470 ^ r512;
  wire _3939 = _3937 ^ _3938;
  wire _3940 = _3936 ^ _3939;
  wire _3941 = r569 ^ r630;
  wire _3942 = r716 ^ r849;
  wire _3943 = _3941 ^ _3942;
  wire _3944 = r914 ^ r946;
  wire _3945 = r1008 ^ r1091;
  wire _3946 = _3944 ^ _3945;
  wire _3947 = _3943 ^ _3946;
  wire _3948 = _3940 ^ _3947;
  wire _3949 = r1110 ^ r1115;
  wire _3950 = r1297 ^ r1344;
  wire _3951 = _3949 ^ _3950;
  wire _3952 = r1543 ^ r1569;
  wire _3953 = r1600 ^ r1636;
  wire _3954 = _3952 ^ _3953;
  wire _3955 = _3951 ^ _3954;
  wire _3956 = r1682 ^ r1722;
  wire _3957 = r1814 ^ r1838;
  wire _3958 = _3956 ^ _3957;
  wire _3959 = r1868 ^ r1876;
  wire _3960 = r1987 ^ r1988;
  wire _3961 = _3959 ^ _3960;
  wire _3962 = _3958 ^ _3961;
  wire _3963 = _3955 ^ _3962;
  wire _3964 = _3948 ^ _3963;
  wire _3965 = _3933 | _3964;
  wire _3966 = _3902 | _3965;
  wire _3967 = r69 ^ r153;
  wire _3968 = r240 ^ r292;
  wire _3969 = _3967 ^ _3968;
  wire _3970 = r364 ^ r414;
  wire _3971 = r476 ^ r542;
  wire _3972 = _3970 ^ _3971;
  wire _3973 = _3969 ^ _3972;
  wire _3974 = r634 ^ r886;
  wire _3975 = r907 ^ r1049;
  wire _3976 = _3974 ^ _3975;
  wire _3977 = r1109 ^ r1133;
  wire _3978 = r1234 ^ r1308;
  wire _3979 = _3977 ^ _3978;
  wire _3980 = _3976 ^ _3979;
  wire _3981 = _3973 ^ _3980;
  wire _3982 = r1370 ^ r1419;
  wire _3983 = r1457 ^ r1597;
  wire _3984 = _3982 ^ _3983;
  wire _3985 = r1608 ^ r1721;
  wire _3986 = r1795 ^ r1821;
  wire _3987 = _3985 ^ _3986;
  wire _3988 = _3984 ^ _3987;
  wire _3989 = r1843 ^ r1856;
  wire _3990 = r1898 ^ r1910;
  wire _3991 = _3989 ^ _3990;
  wire _3992 = r1932 ^ r1962;
  wire _3993 = r1970 ^ r1976;
  wire _3994 = _3992 ^ _3993;
  wire _3995 = _3991 ^ _3994;
  wire _3996 = _3988 ^ _3995;
  wire _3997 = _3981 ^ _3996;
  wire _3998 = r87 ^ r169;
  wire _3999 = r320 ^ r366;
  wire _4000 = _3998 ^ _3999;
  wire _4001 = r431 ^ r465;
  wire _4002 = r539 ^ r596;
  wire _4003 = _4001 ^ _4002;
  wire _4004 = _4000 ^ _4003;
  wire _4005 = r625 ^ r753;
  wire _4006 = r800 ^ r837;
  wire _4007 = _4005 ^ _4006;
  wire _4008 = r936 ^ r1001;
  wire _4009 = r1019 ^ r1078;
  wire _4010 = _4008 ^ _4009;
  wire _4011 = _4007 ^ _4010;
  wire _4012 = _4004 ^ _4011;
  wire _4013 = r1113 ^ r1304;
  wire _4014 = r1356 ^ r1434;
  wire _4015 = _4013 ^ _4014;
  wire _4016 = r1493 ^ r1510;
  wire _4017 = r1539 ^ r1692;
  wire _4018 = _4016 ^ _4017;
  wire _4019 = _4015 ^ _4018;
  wire _4020 = r1719 ^ r1738;
  wire _4021 = r1784 ^ r1816;
  wire _4022 = _4020 ^ _4021;
  wire _4023 = r1859 ^ r1896;
  wire _4024 = r1959 ^ r1964;
  wire _4025 = _4023 ^ _4024;
  wire _4026 = _4022 ^ _4025;
  wire _4027 = _4019 ^ _4026;
  wire _4028 = _4012 ^ _4027;
  wire _4029 = _3997 | _4028;
  wire _4030 = r60 ^ r139;
  wire _4031 = r186 ^ r271;
  wire _4032 = _4030 ^ _4031;
  wire _4033 = r281 ^ r334;
  wire _4034 = r394 ^ r487;
  wire _4035 = _4033 ^ _4034;
  wire _4036 = _4032 ^ _4035;
  wire _4037 = r555 ^ r660;
  wire _4038 = r720 ^ r758;
  wire _4039 = _4037 ^ _4038;
  wire _4040 = r779 ^ r860;
  wire _4041 = r890 ^ r971;
  wire _4042 = _4040 ^ _4041;
  wire _4043 = _4039 ^ _4042;
  wire _4044 = _4036 ^ _4043;
  wire _4045 = r1010 ^ r1079;
  wire _4046 = r1162 ^ r1237;
  wire _4047 = _4045 ^ _4046;
  wire _4048 = r1276 ^ r1323;
  wire _4049 = r1334 ^ r1381;
  wire _4050 = _4048 ^ _4049;
  wire _4051 = _4047 ^ _4050;
  wire _4052 = r1515 ^ r1549;
  wire _4053 = r1586 ^ r1635;
  wire _4054 = _4052 ^ _4053;
  wire _4055 = r1720 ^ r1757;
  wire _4056 = r1764 ^ r1830;
  wire _4057 = _4055 ^ _4056;
  wire _4058 = _4054 ^ _4057;
  wire _4059 = _4051 ^ _4058;
  wire _4060 = _4044 ^ _4059;
  wire _4061 = r52 ^ r57;
  wire _4062 = r117 ^ r173;
  wire _4063 = _4061 ^ _4062;
  wire _4064 = r277 ^ r306;
  wire _4065 = r373 ^ r403;
  wire _4066 = _4064 ^ _4065;
  wire _4067 = _4063 ^ _4066;
  wire _4068 = r494 ^ r548;
  wire _4069 = r597 ^ r644;
  wire _4070 = _4068 ^ _4069;
  wire _4071 = r697 ^ r825;
  wire _4072 = r858 ^ r940;
  wire _4073 = _4071 ^ _4072;
  wire _4074 = _4070 ^ _4073;
  wire _4075 = _4067 ^ _4074;
  wire _4076 = r955 ^ r1054;
  wire _4077 = r1120 ^ r1210;
  wire _4078 = _4076 ^ _4077;
  wire _4079 = r1221 ^ r1240;
  wire _4080 = r1292 ^ r1372;
  wire _4081 = _4079 ^ _4080;
  wire _4082 = _4078 ^ _4081;
  wire _4083 = r1414 ^ r1430;
  wire _4084 = r1499 ^ r1506;
  wire _4085 = _4083 ^ _4084;
  wire _4086 = r1587 ^ r1618;
  wire _4087 = r1706 ^ r1755;
  wire _4088 = _4086 ^ _4087;
  wire _4089 = _4085 ^ _4088;
  wire _4090 = _4082 ^ _4089;
  wire _4091 = _4075 ^ _4090;
  wire _4092 = _4060 | _4091;
  wire _4093 = _4029 | _4092;
  wire _4094 = _3966 | _4093;
  wire _4095 = _3839 | _4094;
  wire _4096 = _3584 | _4095;
  wire _4097 = _3073 | _4096;
  wire _4098 = _2050 | _4097;
  wire _4099 = r53 ^ r108;
  wire _4100 = r129 ^ r198;
  wire _4101 = _4099 ^ _4100;
  wire _4102 = r244 ^ r298;
  wire _4103 = r341 ^ r391;
  wire _4104 = _4102 ^ _4103;
  wire _4105 = _4101 ^ _4104;
  wire _4106 = r441 ^ r457;
  wire _4107 = r534 ^ r579;
  wire _4108 = _4106 ^ _4107;
  wire _4109 = r640 ^ r710;
  wire _4110 = r762 ^ r795;
  wire _4111 = _4109 ^ _4110;
  wire _4112 = _4108 ^ _4111;
  wire _4113 = _4105 ^ _4112;
  wire _4114 = r858 ^ r893;
  wire _4115 = r1002 ^ r1037;
  wire _4116 = _4114 ^ _4115;
  wire _4117 = r1073 ^ r1157;
  wire _4118 = r1170 ^ r1244;
  wire _4119 = _4117 ^ _4118;
  wire _4120 = _4116 ^ _4119;
  wire _4121 = r1286 ^ r1345;
  wire _4122 = r1493 ^ r1573;
  wire _4123 = _4121 ^ _4122;
  wire _4124 = r1581 ^ r1707;
  wire _4125 = r1781 ^ r1831;
  wire _4126 = _4124 ^ _4125;
  wire _4127 = _4123 ^ _4126;
  wire _4128 = _4120 ^ _4127;
  wire _4129 = _4113 ^ _4128;
  wire _4130 = r51 ^ r56;
  wire _4131 = r116 ^ r172;
  wire _4132 = _4130 ^ _4131;
  wire _4133 = r276 ^ r305;
  wire _4134 = r372 ^ r402;
  wire _4135 = _4133 ^ _4134;
  wire _4136 = _4132 ^ _4135;
  wire _4137 = r493 ^ r547;
  wire _4138 = r596 ^ r643;
  wire _4139 = _4137 ^ _4138;
  wire _4140 = r696 ^ r824;
  wire _4141 = r857 ^ r939;
  wire _4142 = _4140 ^ _4141;
  wire _4143 = _4139 ^ _4142;
  wire _4144 = _4136 ^ _4143;
  wire _4145 = r954 ^ r1053;
  wire _4146 = r1107 ^ r1119;
  wire _4147 = _4145 ^ _4146;
  wire _4148 = r1209 ^ r1220;
  wire _4149 = r1291 ^ r1371;
  wire _4150 = _4148 ^ _4149;
  wire _4151 = _4147 ^ _4150;
  wire _4152 = r1413 ^ r1429;
  wire _4153 = r1499 ^ r1586;
  wire _4154 = _4152 ^ _4153;
  wire _4155 = r1617 ^ r1655;
  wire _4156 = r1705 ^ r1756;
  wire _4157 = _4155 ^ _4156;
  wire _4158 = _4154 ^ _4157;
  wire _4159 = _4151 ^ _4158;
  wire _4160 = _4144 ^ _4159;
  wire _4161 = _4129 | _4160;
  wire _4162 = r50 ^ r73;
  wire _4163 = r140 ^ r188;
  wire _4164 = _4162 ^ _4163;
  wire _4165 = r245 ^ r285;
  wire _4166 = r385 ^ r398;
  wire _4167 = _4165 ^ _4166;
  wire _4168 = _4164 ^ _4167;
  wire _4169 = r477 ^ r520;
  wire _4170 = r586 ^ r654;
  wire _4171 = _4169 ^ _4170;
  wire _4172 = r706 ^ r756;
  wire _4173 = r786 ^ r835;
  wire _4174 = _4172 ^ _4173;
  wire _4175 = _4171 ^ _4174;
  wire _4176 = _4168 ^ _4175;
  wire _4177 = r981 ^ r1014;
  wire _4178 = r1099 ^ r1189;
  wire _4179 = _4177 ^ _4178;
  wire _4180 = r1230 ^ r1292;
  wire _4181 = r1359 ^ r1401;
  wire _4182 = _4180 ^ _4181;
  wire _4183 = _4179 ^ _4182;
  wire _4184 = r1439 ^ r1465;
  wire _4185 = r1513 ^ r1556;
  wire _4186 = _4184 ^ _4185;
  wire _4187 = r1620 ^ r1718;
  wire _4188 = r1773 ^ r1832;
  wire _4189 = _4187 ^ _4188;
  wire _4190 = _4186 ^ _4189;
  wire _4191 = _4183 ^ _4190;
  wire _4192 = _4176 ^ _4191;
  wire _4193 = r65 ^ r154;
  wire _4194 = r206 ^ r243;
  wire _4195 = _4193 ^ _4194;
  wire _4196 = r307 ^ r334;
  wire _4197 = r403 ^ r479;
  wire _4198 = _4196 ^ _4197;
  wire _4199 = _4195 ^ _4198;
  wire _4200 = r530 ^ r608;
  wire _4201 = r665 ^ r700;
  wire _4202 = _4200 ^ _4201;
  wire _4203 = r750 ^ r791;
  wire _4204 = r870 ^ r887;
  wire _4205 = _4203 ^ _4204;
  wire _4206 = _4202 ^ _4205;
  wire _4207 = _4199 ^ _4206;
  wire _4208 = r932 ^ r972;
  wire _4209 = r1044 ^ r1064;
  wire _4210 = _4208 ^ _4209;
  wire _4211 = r1143 ^ r1173;
  wire _4212 = r1264 ^ r1321;
  wire _4213 = _4211 ^ _4212;
  wire _4214 = _4210 ^ _4213;
  wire _4215 = r1377 ^ r1551;
  wire _4216 = r1572 ^ r1605;
  wire _4217 = _4215 ^ _4216;
  wire _4218 = r1608 ^ r1674;
  wire _4219 = r1792 ^ r1833;
  wire _4220 = _4218 ^ _4219;
  wire _4221 = _4217 ^ _4220;
  wire _4222 = _4214 ^ _4221;
  wire _4223 = _4207 ^ _4222;
  wire _4224 = _4192 | _4223;
  wire _4225 = _4161 | _4224;
  wire _4226 = r49 ^ r151;
  wire _4227 = r214 ^ r274;
  wire _4228 = _4226 ^ _4227;
  wire _4229 = r321 ^ r364;
  wire _4230 = r448 ^ r615;
  wire _4231 = _4229 ^ _4230;
  wire _4232 = _4228 ^ _4231;
  wire _4233 = r637 ^ r704;
  wire _4234 = r733 ^ r873;
  wire _4235 = _4233 ^ _4234;
  wire _4236 = r914 ^ r959;
  wire _4237 = r1041 ^ r1185;
  wire _4238 = _4236 ^ _4237;
  wire _4239 = _4235 ^ _4238;
  wire _4240 = _4232 ^ _4239;
  wire _4241 = r1247 ^ r1352;
  wire _4242 = r1404 ^ r1482;
  wire _4243 = _4241 ^ _4242;
  wire _4244 = r1500 ^ r1560;
  wire _4245 = r1635 ^ r1778;
  wire _4246 = _4244 ^ _4245;
  wire _4247 = _4243 ^ _4246;
  wire _4248 = r1809 ^ r1940;
  wire _4249 = r1947 ^ r1982;
  wire _4250 = _4248 ^ _4249;
  wire _4251 = r2017 ^ r2042;
  wire _4252 = r2044 ^ r2047;
  wire _4253 = _4251 ^ _4252;
  wire _4254 = _4250 ^ _4253;
  wire _4255 = _4247 ^ _4254;
  wire _4256 = _4240 ^ _4255;
  wire _4257 = r48 ^ r209;
  wire _4258 = r255 ^ r317;
  wire _4259 = _4257 ^ _4258;
  wire _4260 = r380 ^ r416;
  wire _4261 = r527 ^ r600;
  wire _4262 = _4260 ^ _4261;
  wire _4263 = _4259 ^ _4262;
  wire _4264 = r626 ^ r693;
  wire _4265 = r740 ^ r790;
  wire _4266 = _4264 ^ _4265;
  wire _4267 = r860 ^ r896;
  wire _4268 = r978 ^ r1058;
  wire _4269 = _4267 ^ _4268;
  wire _4270 = _4266 ^ _4269;
  wire _4271 = _4263 ^ _4270;
  wire _4272 = r1147 ^ r1194;
  wire _4273 = r1259 ^ r1349;
  wire _4274 = _4272 ^ _4273;
  wire _4275 = r1423 ^ r1441;
  wire _4276 = r1509 ^ r1528;
  wire _4277 = _4275 ^ _4276;
  wire _4278 = _4274 ^ _4277;
  wire _4279 = r1555 ^ r1577;
  wire _4280 = r1675 ^ r1878;
  wire _4281 = _4279 ^ _4280;
  wire _4282 = r1929 ^ r1938;
  wire _4283 = r1945 ^ r1952;
  wire _4284 = _4282 ^ _4283;
  wire _4285 = _4281 ^ _4284;
  wire _4286 = _4278 ^ _4285;
  wire _4287 = _4271 ^ _4286;
  wire _4288 = _4256 | _4287;
  wire _4289 = r47 ^ r100;
  wire _4290 = r134 ^ r258;
  wire _4291 = _4289 ^ _4290;
  wire _4292 = r423 ^ r497;
  wire _4293 = r518 ^ r763;
  wire _4294 = _4292 ^ _4293;
  wire _4295 = _4291 ^ _4294;
  wire _4296 = r950 ^ r1050;
  wire _4297 = r1068 ^ r1151;
  wire _4298 = _4296 ^ _4297;
  wire _4299 = r1271 ^ r1281;
  wire _4300 = r1284 ^ r1607;
  wire _4301 = _4299 ^ _4300;
  wire _4302 = _4298 ^ _4301;
  wire _4303 = _4295 ^ _4302;
  wire _4304 = r1628 ^ r1668;
  wire _4305 = r1694 ^ r1750;
  wire _4306 = _4304 ^ _4305;
  wire _4307 = r1787 ^ r1850;
  wire _4308 = r1856 ^ r1869;
  wire _4309 = _4307 ^ _4308;
  wire _4310 = _4306 ^ _4309;
  wire _4311 = r1880 ^ r1941;
  wire _4312 = r1964 ^ r1965;
  wire _4313 = _4311 ^ _4312;
  wire _4314 = r2001 ^ r2008;
  wire _4315 = r2014 ^ r2023;
  wire _4316 = _4314 ^ _4315;
  wire _4317 = _4313 ^ _4316;
  wire _4318 = _4310 ^ _4317;
  wire _4319 = _4303 ^ _4318;
  wire _4320 = r46 ^ r103;
  wire _4321 = r135 ^ r205;
  wire _4322 = _4320 ^ _4321;
  wire _4323 = r388 ^ r449;
  wire _4324 = r555 ^ r571;
  wire _4325 = _4323 ^ _4324;
  wire _4326 = _4322 ^ _4325;
  wire _4327 = r712 ^ r761;
  wire _4328 = r821 ^ r920;
  wire _4329 = _4327 ^ _4328;
  wire _4330 = r947 ^ r1062;
  wire _4331 = r1140 ^ r1211;
  wire _4332 = _4330 ^ _4331;
  wire _4333 = _4329 ^ _4332;
  wire _4334 = _4326 ^ _4333;
  wire _4335 = r1357 ^ r1387;
  wire _4336 = r1447 ^ r1487;
  wire _4337 = _4335 ^ _4336;
  wire _4338 = r1532 ^ r1537;
  wire _4339 = r1686 ^ r1816;
  wire _4340 = _4338 ^ _4339;
  wire _4341 = _4337 ^ _4340;
  wire _4342 = r1817 ^ r1824;
  wire _4343 = r1846 ^ r1851;
  wire _4344 = _4342 ^ _4343;
  wire _4345 = r1886 ^ r1994;
  wire _4346 = r2005 ^ r2010;
  wire _4347 = _4345 ^ _4346;
  wire _4348 = _4344 ^ _4347;
  wire _4349 = _4341 ^ _4348;
  wire _4350 = _4334 ^ _4349;
  wire _4351 = _4319 | _4350;
  wire _4352 = _4288 | _4351;
  wire _4353 = _4225 | _4352;
  wire _4354 = r45 ^ r94;
  wire _4355 = r111 ^ r175;
  wire _4356 = _4354 ^ _4355;
  wire _4357 = r275 ^ r301;
  wire _4358 = r352 ^ r408;
  wire _4359 = _4357 ^ _4358;
  wire _4360 = _4356 ^ _4359;
  wire _4361 = r478 ^ r537;
  wire _4362 = r607 ^ r649;
  wire _4363 = _4361 ^ _4362;
  wire _4364 = r670 ^ r738;
  wire _4365 = r827 ^ r882;
  wire _4366 = _4364 ^ _4365;
  wire _4367 = _4363 ^ _4366;
  wire _4368 = _4360 ^ _4367;
  wire _4369 = r890 ^ r1097;
  wire _4370 = r1120 ^ r1197;
  wire _4371 = _4369 ^ _4370;
  wire _4372 = r1232 ^ r1283;
  wire _4373 = r1451 ^ r1480;
  wire _4374 = _4372 ^ _4373;
  wire _4375 = _4371 ^ _4374;
  wire _4376 = r1540 ^ r1636;
  wire _4377 = r1777 ^ r1845;
  wire _4378 = _4376 ^ _4377;
  wire _4379 = r1894 ^ r1939;
  wire _4380 = r1949 ^ r1953;
  wire _4381 = _4379 ^ _4380;
  wire _4382 = _4378 ^ _4381;
  wire _4383 = _4375 ^ _4382;
  wire _4384 = _4368 ^ _4383;
  wire _4385 = r44 ^ r74;
  wire _4386 = r161 ^ r182;
  wire _4387 = _4385 ^ _4386;
  wire _4388 = r242 ^ r282;
  wire _4389 = r366 ^ r434;
  wire _4390 = _4388 ^ _4389;
  wire _4391 = _4387 ^ _4390;
  wire _4392 = r492 ^ r551;
  wire _4393 = r564 ^ r656;
  wire _4394 = _4392 ^ _4393;
  wire _4395 = r679 ^ r774;
  wire _4396 = r796 ^ r934;
  wire _4397 = _4395 ^ _4396;
  wire _4398 = _4394 ^ _4397;
  wire _4399 = _4391 ^ _4398;
  wire _4400 = r956 ^ r1028;
  wire _4401 = r1103 ^ r1160;
  wire _4402 = _4400 ^ _4401;
  wire _4403 = r1213 ^ r1274;
  wire _4404 = r1341 ^ r1422;
  wire _4405 = _4403 ^ _4404;
  wire _4406 = _4402 ^ _4405;
  wire _4407 = r1427 ^ r1526;
  wire _4408 = r1678 ^ r1693;
  wire _4409 = _4407 ^ _4408;
  wire _4410 = r1724 ^ r1731;
  wire _4411 = r1893 ^ r1909;
  wire _4412 = _4410 ^ _4411;
  wire _4413 = _4409 ^ _4412;
  wire _4414 = _4406 ^ _4413;
  wire _4415 = _4399 ^ _4414;
  wire _4416 = _4384 | _4415;
  wire _4417 = r43 ^ r55;
  wire _4418 = r120 ^ r218;
  wire _4419 = _4417 ^ _4418;
  wire _4420 = r268 ^ r327;
  wire _4421 = r362 ^ r414;
  wire _4422 = _4420 ^ _4421;
  wire _4423 = _4419 ^ _4422;
  wire _4424 = r466 ^ r506;
  wire _4425 = r572 ^ r653;
  wire _4426 = _4424 ^ _4425;
  wire _4427 = r707 ^ r776;
  wire _4428 = r794 ^ r837;
  wire _4429 = _4427 ^ _4428;
  wire _4430 = _4426 ^ _4429;
  wire _4431 = _4423 ^ _4430;
  wire _4432 = r922 ^ r989;
  wire _4433 = r1031 ^ r1074;
  wire _4434 = _4432 ^ _4433;
  wire _4435 = r1115 ^ r1177;
  wire _4436 = r1310 ^ r1431;
  wire _4437 = _4435 ^ _4436;
  wire _4438 = _4434 ^ _4437;
  wire _4439 = r1450 ^ r1461;
  wire _4440 = r1618 ^ r1680;
  wire _4441 = _4439 ^ _4440;
  wire _4442 = r1712 ^ r1744;
  wire _4443 = r1794 ^ r1834;
  wire _4444 = _4442 ^ _4443;
  wire _4445 = _4441 ^ _4444;
  wire _4446 = _4438 ^ _4445;
  wire _4447 = _4431 ^ _4446;
  wire _4448 = r42 ^ r69;
  wire _4449 = r124 ^ r220;
  wire _4450 = _4448 ^ _4449;
  wire _4451 = r252 ^ r289;
  wire _4452 = r383 ^ r426;
  wire _4453 = _4451 ^ _4452;
  wire _4454 = _4450 ^ _4453;
  wire _4455 = r500 ^ r531;
  wire _4456 = r601 ^ r657;
  wire _4457 = _4455 ^ _4456;
  wire _4458 = r695 ^ r884;
  wire _4459 = r937 ^ r999;
  wire _4460 = _4458 ^ _4459;
  wire _4461 = _4457 ^ _4460;
  wire _4462 = _4454 ^ _4461;
  wire _4463 = r1022 ^ r1072;
  wire _4464 = r1126 ^ r1186;
  wire _4465 = _4463 ^ _4464;
  wire _4466 = r1253 ^ r1317;
  wire _4467 = r1338 ^ r1386;
  wire _4468 = _4466 ^ _4467;
  wire _4469 = _4465 ^ _4468;
  wire _4470 = r1396 ^ r1445;
  wire _4471 = r1582 ^ r1633;
  wire _4472 = _4470 ^ _4471;
  wire _4473 = r1746 ^ r1779;
  wire _4474 = r1815 ^ r1881;
  wire _4475 = _4473 ^ _4474;
  wire _4476 = _4472 ^ _4475;
  wire _4477 = _4469 ^ _4476;
  wire _4478 = _4462 ^ _4477;
  wire _4479 = _4447 | _4478;
  wire _4480 = _4416 | _4479;
  wire _4481 = r41 ^ r80;
  wire _4482 = r170 ^ r191;
  wire _4483 = _4481 ^ _4482;
  wire _4484 = r277 ^ r293;
  wire _4485 = r346 ^ r435;
  wire _4486 = _4484 ^ _4485;
  wire _4487 = _4483 ^ _4486;
  wire _4488 = r467 ^ r519;
  wire _4489 = r614 ^ r648;
  wire _4490 = _4488 ^ _4489;
  wire _4491 = r681 ^ r739;
  wire _4492 = r806 ^ r871;
  wire _4493 = _4491 ^ _4492;
  wire _4494 = _4490 ^ _4493;
  wire _4495 = _4487 ^ _4494;
  wire _4496 = r902 ^ r992;
  wire _4497 = r1101 ^ r1154;
  wire _4498 = _4496 ^ _4497;
  wire _4499 = r1182 ^ r1261;
  wire _4500 = r1278 ^ r1287;
  wire _4501 = _4499 ^ _4500;
  wire _4502 = _4498 ^ _4501;
  wire _4503 = r1467 ^ r1504;
  wire _4504 = r1533 ^ r1544;
  wire _4505 = _4503 ^ _4504;
  wire _4506 = r1580 ^ r1611;
  wire _4507 = r1708 ^ r1757;
  wire _4508 = _4506 ^ _4507;
  wire _4509 = _4505 ^ _4508;
  wire _4510 = _4502 ^ _4509;
  wire _4511 = _4495 ^ _4510;
  wire _4512 = r123 ^ r173;
  wire _4513 = r269 ^ r332;
  wire _4514 = _4512 ^ _4513;
  wire _4515 = r347 ^ r407;
  wire _4516 = r480 ^ r508;
  wire _4517 = _4515 ^ _4516;
  wire _4518 = _4514 ^ _4517;
  wire _4519 = r618 ^ r698;
  wire _4520 = r760 ^ r809;
  wire _4521 = _4519 ^ _4520;
  wire _4522 = r834 ^ r911;
  wire _4523 = r996 ^ r1040;
  wire _4524 = _4522 ^ _4523;
  wire _4525 = _4521 ^ _4524;
  wire _4526 = _4518 ^ _4525;
  wire _4527 = r1085 ^ r1142;
  wire _4528 = r1187 ^ r1332;
  wire _4529 = _4527 ^ _4528;
  wire _4530 = r1364 ^ r1459;
  wire _4531 = r1474 ^ r1546;
  wire _4532 = _4530 ^ _4531;
  wire _4533 = _4529 ^ _4532;
  wire _4534 = r1741 ^ r1788;
  wire _4535 = r1810 ^ r1814;
  wire _4536 = _4534 ^ _4535;
  wire _4537 = r1848 ^ r1872;
  wire _4538 = r1879 ^ r1910;
  wire _4539 = _4537 ^ _4538;
  wire _4540 = _4536 ^ _4539;
  wire _4541 = _4533 ^ _4540;
  wire _4542 = _4526 ^ _4541;
  wire _4543 = _4511 | _4542;
  wire _4544 = r40 ^ r96;
  wire _4545 = r118 ^ r256;
  wire _4546 = _4544 ^ _4545;
  wire _4547 = r382 ^ r422;
  wire _4548 = r522 ^ r567;
  wire _4549 = _4547 ^ _4548;
  wire _4550 = _4546 ^ _4549;
  wire _4551 = r623 ^ r907;
  wire _4552 = r986 ^ r1054;
  wire _4553 = _4551 ^ _4552;
  wire _4554 = r1129 ^ r1262;
  wire _4555 = r1315 ^ r1348;
  wire _4556 = _4554 ^ _4555;
  wire _4557 = _4553 ^ _4556;
  wire _4558 = _4550 ^ _4557;
  wire _4559 = r1408 ^ r1623;
  wire _4560 = r1658 ^ r1747;
  wire _4561 = _4559 ^ _4560;
  wire _4562 = r1797 ^ r1818;
  wire _4563 = r1827 ^ r1873;
  wire _4564 = _4562 ^ _4563;
  wire _4565 = _4561 ^ _4564;
  wire _4566 = r1899 ^ r1902;
  wire _4567 = r1918 ^ r1955;
  wire _4568 = _4566 ^ _4567;
  wire _4569 = r1973 ^ r1989;
  wire _4570 = r1998 ^ r2003;
  wire _4571 = _4569 ^ _4570;
  wire _4572 = _4568 ^ _4571;
  wire _4573 = _4565 ^ _4572;
  wire _4574 = _4558 ^ _4573;
  wire _4575 = r39 ^ r83;
  wire _4576 = r158 ^ r192;
  wire _4577 = _4575 ^ _4576;
  wire _4578 = r273 ^ r287;
  wire _4579 = r373 ^ r394;
  wire _4580 = _4578 ^ _4579;
  wire _4581 = _4577 ^ _4580;
  wire _4582 = r495 ^ r543;
  wire _4583 = r589 ^ r661;
  wire _4584 = _4582 ^ _4583;
  wire _4585 = r671 ^ r771;
  wire _4586 = r862 ^ r912;
  wire _4587 = _4585 ^ _4586;
  wire _4588 = _4584 ^ _4587;
  wire _4589 = _4581 ^ _4588;
  wire _4590 = r964 ^ r1008;
  wire _4591 = r1075 ^ r1145;
  wire _4592 = _4590 ^ _4591;
  wire _4593 = r1199 ^ r1252;
  wire _4594 = r1299 ^ r1360;
  wire _4595 = _4593 ^ _4594;
  wire _4596 = _4592 ^ _4595;
  wire _4597 = r1391 ^ r1436;
  wire _4598 = r1455 ^ r1592;
  wire _4599 = _4597 ^ _4598;
  wire _4600 = r1615 ^ r1679;
  wire _4601 = r1688 ^ r1758;
  wire _4602 = _4600 ^ _4601;
  wire _4603 = _4599 ^ _4602;
  wire _4604 = _4596 ^ _4603;
  wire _4605 = _4589 ^ _4604;
  wire _4606 = _4574 | _4605;
  wire _4607 = _4543 | _4606;
  wire _4608 = _4480 | _4607;
  wire _4609 = _4353 | _4608;
  wire _4610 = r38 ^ r98;
  wire _4611 = r166 ^ r219;
  wire _4612 = _4610 ^ _4611;
  wire _4613 = r249 ^ r324;
  wire _4614 = r333 ^ r429;
  wire _4615 = _4613 ^ _4614;
  wire _4616 = _4612 ^ _4615;
  wire _4617 = r462 ^ r553;
  wire _4618 = r602 ^ r663;
  wire _4619 = _4617 ^ _4618;
  wire _4620 = r720 ^ r741;
  wire _4621 = r793 ^ r876;
  wire _4622 = _4620 ^ _4621;
  wire _4623 = _4619 ^ _4622;
  wire _4624 = _4616 ^ _4623;
  wire _4625 = r901 ^ r946;
  wire _4626 = r1034 ^ r1102;
  wire _4627 = _4625 ^ _4626;
  wire _4628 = r1206 ^ r1301;
  wire _4629 = r1330 ^ r1370;
  wire _4630 = _4628 ^ _4629;
  wire _4631 = _4627 ^ _4630;
  wire _4632 = r1400 ^ r1511;
  wire _4633 = r1520 ^ r1566;
  wire _4634 = _4632 ^ _4633;
  wire _4635 = r1583 ^ r1643;
  wire _4636 = r1785 ^ r1835;
  wire _4637 = _4635 ^ _4636;
  wire _4638 = _4634 ^ _4637;
  wire _4639 = _4631 ^ _4638;
  wire _4640 = _4624 ^ _4639;
  wire _4641 = r37 ^ r61;
  wire _4642 = r130 ^ r181;
  wire _4643 = _4641 ^ _4642;
  wire _4644 = r247 ^ r331;
  wire _4645 = r336 ^ r396;
  wire _4646 = _4644 ^ _4645;
  wire _4647 = _4643 ^ _4646;
  wire _4648 = r463 ^ r548;
  wire _4649 = r599 ^ r631;
  wire _4650 = _4648 ^ _4649;
  wire _4651 = r672 ^ r732;
  wire _4652 = r819 ^ r868;
  wire _4653 = _4651 ^ _4652;
  wire _4654 = _4650 ^ _4653;
  wire _4655 = _4647 ^ _4654;
  wire _4656 = r925 ^ r960;
  wire _4657 = r1024 ^ r1071;
  wire _4658 = _4656 ^ _4657;
  wire _4659 = r1117 ^ r1165;
  wire _4660 = r1191 ^ r1227;
  wire _4661 = _4659 ^ _4660;
  wire _4662 = _4658 ^ _4661;
  wire _4663 = r1288 ^ r1342;
  wire _4664 = r1409 ^ r1442;
  wire _4665 = _4663 ^ _4664;
  wire _4666 = r1460 ^ r1492;
  wire _4667 = r1669 ^ r1759;
  wire _4668 = _4666 ^ _4667;
  wire _4669 = _4665 ^ _4668;
  wire _4670 = _4662 ^ _4669;
  wire _4671 = _4655 ^ _4670;
  wire _4672 = _4640 | _4671;
  wire _4673 = r36 ^ r71;
  wire _4674 = r128 ^ r261;
  wire _4675 = _4673 ^ _4674;
  wire _4676 = r299 ^ r494;
  wire _4677 = r562 ^ r716;
  wire _4678 = _4676 ^ _4677;
  wire _4679 = _4675 ^ _4678;
  wire _4680 = r775 ^ r803;
  wire _4681 = r845 ^ r971;
  wire _4682 = _4680 ^ _4681;
  wire _4683 = r1011 ^ r1266;
  wire _4684 = r1316 ^ r1457;
  wire _4685 = _4683 ^ _4684;
  wire _4686 = _4682 ^ _4685;
  wire _4687 = _4679 ^ _4686;
  wire _4688 = r1496 ^ r1535;
  wire _4689 = r1545 ^ r1646;
  wire _4690 = _4688 ^ _4689;
  wire _4691 = r1654 ^ r1689;
  wire _4692 = r1854 ^ r1890;
  wire _4693 = _4691 ^ _4692;
  wire _4694 = _4690 ^ _4693;
  wire _4695 = r1946 ^ r1948;
  wire _4696 = r1972 ^ r1980;
  wire _4697 = _4695 ^ _4696;
  wire _4698 = r1991 ^ r1997;
  wire _4699 = r2032 ^ r2039;
  wire _4700 = _4698 ^ _4699;
  wire _4701 = _4697 ^ _4700;
  wire _4702 = _4694 ^ _4701;
  wire _4703 = _4687 ^ _4702;
  wire _4704 = r35 ^ r66;
  wire _4705 = r164 ^ r187;
  wire _4706 = _4704 ^ _4705;
  wire _4707 = r253 ^ r297;
  wire _4708 = r335 ^ r406;
  wire _4709 = _4707 ^ _4708;
  wire _4710 = _4706 ^ _4709;
  wire _4711 = r485 ^ r542;
  wire _4712 = r583 ^ r625;
  wire _4713 = _4711 ^ _4712;
  wire _4714 = r684 ^ r722;
  wire _4715 = r737 ^ r828;
  wire _4716 = _4714 ^ _4715;
  wire _4717 = _4713 ^ _4716;
  wire _4718 = _4710 ^ _4717;
  wire _4719 = r855 ^ r915;
  wire _4720 = r1026 ^ r1081;
  wire _4721 = _4719 ^ _4720;
  wire _4722 = r1118 ^ r1215;
  wire _4723 = r1268 ^ r1285;
  wire _4724 = _4722 ^ _4723;
  wire _4725 = _4721 ^ _4724;
  wire _4726 = r1373 ^ r1489;
  wire _4727 = r1567 ^ r1600;
  wire _4728 = _4726 ^ _4727;
  wire _4729 = r1739 ^ r1752;
  wire _4730 = r1807 ^ r1836;
  wire _4731 = _4729 ^ _4730;
  wire _4732 = _4728 ^ _4731;
  wire _4733 = _4725 ^ _4732;
  wire _4734 = _4718 ^ _4733;
  wire _4735 = _4703 | _4734;
  wire _4736 = _4672 | _4735;
  wire _4737 = r34 ^ r72;
  wire _4738 = r143 ^ r207;
  wire _4739 = _4737 ^ _4738;
  wire _4740 = r231 ^ r329;
  wire _4741 = r390 ^ r424;
  wire _4742 = _4740 ^ _4741;
  wire _4743 = _4739 ^ _4742;
  wire _4744 = r504 ^ r510;
  wire _4745 = r584 ^ r632;
  wire _4746 = _4744 ^ _4745;
  wire _4747 = r690 ^ r768;
  wire _4748 = r820 ^ r849;
  wire _4749 = _4747 ^ _4748;
  wire _4750 = _4746 ^ _4749;
  wire _4751 = _4743 ^ _4750;
  wire _4752 = r917 ^ r988;
  wire _4753 = r1046 ^ r1104;
  wire _4754 = _4752 ^ _4753;
  wire _4755 = r1198 ^ r1238;
  wire _4756 = r1308 ^ r1331;
  wire _4757 = _4755 ^ _4756;
  wire _4758 = _4754 ^ _4757;
  wire _4759 = r1335 ^ r1424;
  wire _4760 = r1435 ^ r1510;
  wire _4761 = _4759 ^ _4760;
  wire _4762 = r1589 ^ r1640;
  wire _4763 = r1803 ^ r1837;
  wire _4764 = _4762 ^ _4763;
  wire _4765 = _4761 ^ _4764;
  wire _4766 = _4758 ^ _4765;
  wire _4767 = _4751 ^ _4766;
  wire _4768 = r33 ^ r60;
  wire _4769 = r146 ^ r221;
  wire _4770 = _4768 ^ _4769;
  wire _4771 = r241 ^ r309;
  wire _4772 = r370 ^ r446;
  wire _4773 = _4771 ^ _4772;
  wire _4774 = _4770 ^ _4773;
  wire _4775 = r452 ^ r516;
  wire _4776 = r561 ^ r662;
  wire _4777 = _4775 ^ _4776;
  wire _4778 = r675 ^ r765;
  wire _4779 = r807 ^ r853;
  wire _4780 = _4778 ^ _4779;
  wire _4781 = _4777 ^ _4780;
  wire _4782 = _4774 ^ _4781;
  wire _4783 = r941 ^ r974;
  wire _4784 = r1056 ^ r1096;
  wire _4785 = _4783 ^ _4784;
  wire _4786 = r1131 ^ r1210;
  wire _4787 = r1275 ^ r1296;
  wire _4788 = _4786 ^ _4787;
  wire _4789 = _4785 ^ _4788;
  wire _4790 = r1354 ^ r1403;
  wire _4791 = r1454 ^ r1462;
  wire _4792 = _4790 ^ _4791;
  wire _4793 = r1473 ^ r1624;
  wire _4794 = r1726 ^ r1838;
  wire _4795 = _4793 ^ _4794;
  wire _4796 = _4792 ^ _4795;
  wire _4797 = _4789 ^ _4796;
  wire _4798 = _4782 ^ _4797;
  wire _4799 = _4767 | _4798;
  wire _4800 = r32 ^ r86;
  wire _4801 = r131 ^ r217;
  wire _4802 = _4800 ^ _4801;
  wire _4803 = r312 ^ r378;
  wire _4804 = r392 ^ r505;
  wire _4805 = _4803 ^ _4804;
  wire _4806 = _4802 ^ _4805;
  wire _4807 = r557 ^ r622;
  wire _4808 = r826 ^ r842;
  wire _4809 = _4807 ^ _4808;
  wire _4810 = r923 ^ r991;
  wire _4811 = r1051 ^ r1086;
  wire _4812 = _4810 ^ _4811;
  wire _4813 = _4809 ^ _4812;
  wire _4814 = _4806 ^ _4813;
  wire _4815 = r1138 ^ r1216;
  wire _4816 = r1231 ^ r1276;
  wire _4817 = _4815 ^ _4816;
  wire _4818 = r1318 ^ r1362;
  wire _4819 = r1388 ^ r1602;
  wire _4820 = _4818 ^ _4819;
  wire _4821 = _4817 ^ _4820;
  wire _4822 = r1749 ^ r1805;
  wire _4823 = r1847 ^ r1858;
  wire _4824 = _4822 ^ _4823;
  wire _4825 = r1859 ^ r1911;
  wire _4826 = r1925 ^ r1930;
  wire _4827 = _4825 ^ _4826;
  wire _4828 = _4824 ^ _4827;
  wire _4829 = _4821 ^ _4828;
  wire _4830 = _4814 ^ _4829;
  wire _4831 = r31 ^ r92;
  wire _4832 = r165 ^ r184;
  wire _4833 = _4831 ^ _4832;
  wire _4834 = r238 ^ r342;
  wire _4835 = r451 ^ r570;
  wire _4836 = _4834 ^ _4835;
  wire _4837 = _4833 ^ _4836;
  wire _4838 = r650 ^ r702;
  wire _4839 = r800 ^ r933;
  wire _4840 = _4838 ^ _4839;
  wire _4841 = r952 ^ r1057;
  wire _4842 = r1110 ^ r1192;
  wire _4843 = _4841 ^ _4842;
  wire _4844 = _4840 ^ _4843;
  wire _4845 = _4837 ^ _4844;
  wire _4846 = r1239 ^ r1547;
  wire _4847 = r1562 ^ r1619;
  wire _4848 = _4846 ^ _4847;
  wire _4849 = r1667 ^ r1714;
  wire _4850 = r1822 ^ r1864;
  wire _4851 = _4849 ^ _4850;
  wire _4852 = _4848 ^ _4851;
  wire _4853 = r1867 ^ r1912;
  wire _4854 = r1950 ^ r2021;
  wire _4855 = _4853 ^ _4854;
  wire _4856 = r2029 ^ r2031;
  wire _4857 = r2034 ^ r2041;
  wire _4858 = _4856 ^ _4857;
  wire _4859 = _4855 ^ _4858;
  wire _4860 = _4852 ^ _4859;
  wire _4861 = _4845 ^ _4860;
  wire _4862 = _4830 | _4861;
  wire _4863 = _4799 | _4862;
  wire _4864 = _4736 | _4863;
  wire _4865 = r30 ^ r76;
  wire _4866 = r127 ^ r202;
  wire _4867 = _4865 ^ _4866;
  wire _4868 = r228 ^ r330;
  wire _4869 = r340 ^ r415;
  wire _4870 = _4868 ^ _4869;
  wire _4871 = _4867 ^ _4870;
  wire _4872 = r502 ^ r525;
  wire _4873 = r575 ^ r628;
  wire _4874 = _4872 ^ _4873;
  wire _4875 = r682 ^ r748;
  wire _4876 = r798 ^ r861;
  wire _4877 = _4875 ^ _4876;
  wire _4878 = _4874 ^ _4877;
  wire _4879 = _4871 ^ _4878;
  wire _4880 = r942 ^ r962;
  wire _4881 = r1045 ^ r1079;
  wire _4882 = _4880 ^ _4881;
  wire _4883 = r1123 ^ r1205;
  wire _4884 = r1267 ^ r1300;
  wire _4885 = _4883 ^ _4884;
  wire _4886 = _4882 ^ _4885;
  wire _4887 = r1363 ^ r1390;
  wire _4888 = r1458 ^ r1543;
  wire _4889 = _4887 ^ _4888;
  wire _4890 = r1711 ^ r1742;
  wire _4891 = r1802 ^ r1839;
  wire _4892 = _4890 ^ _4891;
  wire _4893 = _4889 ^ _4892;
  wire _4894 = _4886 ^ _4893;
  wire _4895 = _4879 ^ _4894;
  wire _4896 = r29 ^ r78;
  wire _4897 = r155 ^ r203;
  wire _4898 = _4896 ^ _4897;
  wire _4899 = r262 ^ r296;
  wire _4900 = r376 ^ r433;
  wire _4901 = _4899 ^ _4900;
  wire _4902 = _4898 ^ _4901;
  wire _4903 = r509 ^ r616;
  wire _4904 = r652 ^ r694;
  wire _4905 = _4903 ^ _4904;
  wire _4906 = r758 ^ r812;
  wire _4907 = r872 ^ r916;
  wire _4908 = _4906 ^ _4907;
  wire _4909 = _4905 ^ _4908;
  wire _4910 = _4902 ^ _4909;
  wire _4911 = r957 ^ r1077;
  wire _4912 = r1149 ^ r1178;
  wire _4913 = _4911 ^ _4912;
  wire _4914 = r1226 ^ r1314;
  wire _4915 = r1353 ^ r1398;
  wire _4916 = _4914 ^ _4915;
  wire _4917 = _4913 ^ _4916;
  wire _4918 = r1437 ^ r1484;
  wire _4919 = r1553 ^ r1587;
  wire _4920 = _4918 ^ _4919;
  wire _4921 = r1651 ^ r1699;
  wire _4922 = r1729 ^ r1840;
  wire _4923 = _4921 ^ _4922;
  wire _4924 = _4920 ^ _4923;
  wire _4925 = _4917 ^ _4924;
  wire _4926 = _4910 ^ _4925;
  wire _4927 = _4895 | _4926;
  wire _4928 = r28 ^ r139;
  wire _4929 = r183 ^ r246;
  wire _4930 = _4928 ^ _4929;
  wire _4931 = r322 ^ r490;
  wire _4932 = r574 ^ r703;
  wire _4933 = _4931 ^ _4932;
  wire _4934 = _4930 ^ _4933;
  wire _4935 = r751 ^ r805;
  wire _4936 = r883 ^ r930;
  wire _4937 = _4935 ^ _4936;
  wire _4938 = r963 ^ r1020;
  wire _4939 = r1166 ^ r1254;
  wire _4940 = _4938 ^ _4939;
  wire _4941 = _4937 ^ _4940;
  wire _4942 = _4934 ^ _4941;
  wire _4943 = r1376 ^ r1420;
  wire _4944 = r1434 ^ r1584;
  wire _4945 = _4943 ^ _4944;
  wire _4946 = r1642 ^ r1685;
  wire _4947 = r1706 ^ r1855;
  wire _4948 = _4946 ^ _4947;
  wire _4949 = _4945 ^ _4948;
  wire _4950 = r1868 ^ r1891;
  wire _4951 = r1942 ^ r1999;
  wire _4952 = _4950 ^ _4951;
  wire _4953 = r2013 ^ r2015;
  wire _4954 = r2045 ^ r2046;
  wire _4955 = _4953 ^ _4954;
  wire _4956 = _4952 ^ _4955;
  wire _4957 = _4949 ^ _4956;
  wire _4958 = _4942 ^ _4957;
  wire _4959 = r27 ^ r84;
  wire _4960 = r167 ^ r174;
  wire _4961 = _4959 ^ _4960;
  wire _4962 = r257 ^ r306;
  wire _4963 = r357 ^ r447;
  wire _4964 = _4962 ^ _4963;
  wire _4965 = _4961 ^ _4964;
  wire _4966 = r458 ^ r526;
  wire _4967 = r569 ^ r660;
  wire _4968 = _4966 ^ _4967;
  wire _4969 = r676 ^ r755;
  wire _4970 = r782 ^ r856;
  wire _4971 = _4969 ^ _4970;
  wire _4972 = _4968 ^ _4971;
  wire _4973 = _4965 ^ _4972;
  wire _4974 = r903 ^ r951;
  wire _4975 = r1005 ^ r1083;
  wire _4976 = _4974 ^ _4975;
  wire _4977 = r1141 ^ r1180;
  wire _4978 = r1234 ^ r1290;
  wire _4979 = _4977 ^ _4978;
  wire _4980 = _4976 ^ _4979;
  wire _4981 = r1329 ^ r1382;
  wire _4982 = r1421 ^ r1456;
  wire _4983 = _4981 ^ _4982;
  wire _4984 = r1595 ^ r1657;
  wire _4985 = r1702 ^ r1760;
  wire _4986 = _4984 ^ _4985;
  wire _4987 = _4983 ^ _4986;
  wire _4988 = _4980 ^ _4987;
  wire _4989 = _4973 ^ _4988;
  wire _4990 = _4958 | _4989;
  wire _4991 = _4927 | _4990;
  wire _4992 = r26 ^ r95;
  wire _4993 = r157 ^ r343;
  wire _4994 = _4992 ^ _4993;
  wire _4995 = r437 ^ r456;
  wire _4996 = r558 ^ r605;
  wire _4997 = _4995 ^ _4996;
  wire _4998 = _4994 ^ _4997;
  wire _4999 = r745 ^ r844;
  wire _5000 = r936 ^ r977;
  wire _5001 = _4999 ^ _5000;
  wire _5002 = r1003 ^ r1006;
  wire _5003 = r1150 ^ r1255;
  wire _5004 = _5002 ^ _5003;
  wire _5005 = _5001 ^ _5004;
  wire _5006 = _4998 ^ _5005;
  wire _5007 = r1303 ^ r1366;
  wire _5008 = r1397 ^ r1508;
  wire _5009 = _5007 ^ _5008;
  wire _5010 = r1644 ^ r1661;
  wire _5011 = r1728 ^ r1789;
  wire _5012 = _5010 ^ _5011;
  wire _5013 = _5009 ^ _5012;
  wire _5014 = r1913 ^ r1921;
  wire _5015 = r1936 ^ r1971;
  wire _5016 = _5014 ^ _5015;
  wire _5017 = r1975 ^ r1984;
  wire _5018 = r2019 ^ r2022;
  wire _5019 = _5017 ^ _5018;
  wire _5020 = _5016 ^ _5019;
  wire _5021 = _5013 ^ _5020;
  wire _5022 = _5006 ^ _5021;
  wire _5023 = r25 ^ r102;
  wire _5024 = r144 ^ r194;
  wire _5025 = _5023 ^ _5024;
  wire _5026 = r323 ^ r377;
  wire _5027 = r431 ^ r488;
  wire _5028 = _5026 ^ _5027;
  wire _5029 = _5025 ^ _5028;
  wire _5030 = r515 ^ r612;
  wire _5031 = r645 ^ r717;
  wire _5032 = _5030 ^ _5031;
  wire _5033 = r725 ^ r785;
  wire _5034 = r830 ^ r886;
  wire _5035 = _5033 ^ _5034;
  wire _5036 = _5032 ^ _5035;
  wire _5037 = _5029 ^ _5036;
  wire _5038 = r905 ^ r983;
  wire _5039 = r1029 ^ r1069;
  wire _5040 = _5038 ^ _5039;
  wire _5041 = r1122 ^ r1190;
  wire _5042 = r1269 ^ r1297;
  wire _5043 = _5041 ^ _5042;
  wire _5044 = _5040 ^ _5043;
  wire _5045 = r1368 ^ r1384;
  wire _5046 = r1392 ^ r1477;
  wire _5047 = _5045 ^ _5046;
  wire _5048 = r1612 ^ r1687;
  wire _5049 = r1696 ^ r1761;
  wire _5050 = _5048 ^ _5049;
  wire _5051 = _5047 ^ _5050;
  wire _5052 = _5044 ^ _5051;
  wire _5053 = _5037 ^ _5052;
  wire _5054 = _5022 | _5053;
  wire _5055 = r24 ^ r77;
  wire _5056 = r163 ^ r224;
  wire _5057 = _5055 ^ _5056;
  wire _5058 = r230 ^ r310;
  wire _5059 = r339 ^ r412;
  wire _5060 = _5058 ^ _5059;
  wire _5061 = _5057 ^ _5060;
  wire _5062 = r470 ^ r544;
  wire _5063 = r580 ^ r646;
  wire _5064 = _5062 ^ _5063;
  wire _5065 = r697 ^ r764;
  wire _5066 = r789 ^ r847;
  wire _5067 = _5065 ^ _5066;
  wire _5068 = _5064 ^ _5067;
  wire _5069 = _5061 ^ _5068;
  wire _5070 = r918 ^ r966;
  wire _5071 = r1012 ^ r1063;
  wire _5072 = _5070 ^ _5071;
  wire _5073 = r1137 ^ r1208;
  wire _5074 = r1218 ^ r1265;
  wire _5075 = _5073 ^ _5074;
  wire _5076 = _5072 ^ _5075;
  wire _5077 = r1326 ^ r1337;
  wire _5078 = r1407 ^ r1475;
  wire _5079 = _5077 ^ _5078;
  wire _5080 = r1578 ^ r1621;
  wire _5081 = r1660 ^ r1762;
  wire _5082 = _5080 ^ _5081;
  wire _5083 = _5079 ^ _5082;
  wire _5084 = _5076 ^ _5083;
  wire _5085 = _5069 ^ _5084;
  wire _5086 = r23 ^ r91;
  wire _5087 = r136 ^ r271;
  wire _5088 = _5086 ^ _5087;
  wire _5089 = r367 ^ r420;
  wire _5090 = r473 ^ r521;
  wire _5091 = _5089 ^ _5090;
  wire _5092 = _5088 ^ _5091;
  wire _5093 = r578 ^ r624;
  wire _5094 = r866 ^ r968;
  wire _5095 = _5093 ^ _5094;
  wire _5096 = r1023 ^ r1067;
  wire _5097 = r1113 ^ r1229;
  wire _5098 = _5096 ^ _5097;
  wire _5099 = _5095 ^ _5098;
  wire _5100 = _5092 ^ _5099;
  wire _5101 = r1374 ^ r1481;
  wire _5102 = r1512 ^ r1616;
  wire _5103 = _5101 ^ _5102;
  wire _5104 = r1735 ^ r1755;
  wire _5105 = r1775 ^ r1900;
  wire _5106 = _5104 ^ _5105;
  wire _5107 = _5103 ^ _5106;
  wire _5108 = r1951 ^ r1956;
  wire _5109 = r1958 ^ r1967;
  wire _5110 = _5108 ^ _5109;
  wire _5111 = r1969 ^ r1974;
  wire _5112 = r1985 ^ r1987;
  wire _5113 = _5111 ^ _5112;
  wire _5114 = _5110 ^ _5113;
  wire _5115 = _5107 ^ _5114;
  wire _5116 = _5100 ^ _5115;
  wire _5117 = _5085 | _5116;
  wire _5118 = _5054 | _5117;
  wire _5119 = _4991 | _5118;
  wire _5120 = _4864 | _5119;
  wire _5121 = _4609 | _5120;
  wire _5122 = r22 ^ r62;
  wire _5123 = r133 ^ r189;
  wire _5124 = _5122 ^ _5123;
  wire _5125 = r233 ^ r302;
  wire _5126 = r351 ^ r442;
  wire _5127 = _5125 ^ _5126;
  wire _5128 = _5124 ^ _5127;
  wire _5129 = r459 ^ r546;
  wire _5130 = r610 ^ r617;
  wire _5131 = _5129 ^ _5130;
  wire _5132 = r677 ^ r731;
  wire _5133 = r813 ^ r874;
  wire _5134 = _5132 ^ _5133;
  wire _5135 = _5131 ^ _5134;
  wire _5136 = _5128 ^ _5135;
  wire _5137 = r931 ^ r994;
  wire _5138 = r1030 ^ r1109;
  wire _5139 = _5137 ^ _5138;
  wire _5140 = r1144 ^ r1175;
  wire _5141 = r1249 ^ r1443;
  wire _5142 = _5140 ^ _5141;
  wire _5143 = _5139 ^ _5142;
  wire _5144 = r1527 ^ r1534;
  wire _5145 = r1552 ^ r1565;
  wire _5146 = _5144 ^ _5145;
  wire _5147 = r1576 ^ r1622;
  wire _5148 = r1683 ^ r1763;
  wire _5149 = _5147 ^ _5148;
  wire _5150 = _5146 ^ _5149;
  wire _5151 = _5143 ^ _5150;
  wire _5152 = _5136 ^ _5151;
  wire _5153 = r21 ^ r97;
  wire _5154 = r149 ^ r171;
  wire _5155 = _5153 ^ _5154;
  wire _5156 = r250 ^ r300;
  wire _5157 = r379 ^ r440;
  wire _5158 = _5156 ^ _5157;
  wire _5159 = _5155 ^ _5158;
  wire _5160 = r489 ^ r559;
  wire _5161 = r630 ^ r674;
  wire _5162 = _5160 ^ _5161;
  wire _5163 = r759 ^ r797;
  wire _5164 = r869 ^ r898;
  wire _5165 = _5163 ^ _5164;
  wire _5166 = _5162 ^ _5165;
  wire _5167 = _5159 ^ _5166;
  wire _5168 = r975 ^ r1207;
  wire _5169 = r1250 ^ r1411;
  wire _5170 = _5168 ^ _5169;
  wire _5171 = r1452 ^ r1531;
  wire _5172 = r1570 ^ r1650;
  wire _5173 = _5171 ^ _5172;
  wire _5174 = _5170 ^ _5173;
  wire _5175 = r1743 ^ r1745;
  wire _5176 = r1784 ^ r1790;
  wire _5177 = _5175 ^ _5176;
  wire _5178 = r1823 ^ r1830;
  wire _5179 = r1861 ^ r1882;
  wire _5180 = _5178 ^ _5179;
  wire _5181 = _5177 ^ _5180;
  wire _5182 = _5174 ^ _5181;
  wire _5183 = _5167 ^ _5182;
  wire _5184 = _5152 | _5183;
  wire _5185 = r20 ^ r64;
  wire _5186 = r141 ^ r179;
  wire _5187 = _5185 ^ _5186;
  wire _5188 = r259 ^ r315;
  wire _5189 = r369 ^ r418;
  wire _5190 = _5188 ^ _5189;
  wire _5191 = _5187 ^ _5190;
  wire _5192 = r455 ^ r556;
  wire _5193 = r594 ^ r635;
  wire _5194 = _5192 ^ _5193;
  wire _5195 = r692 ^ r747;
  wire _5196 = r808 ^ r875;
  wire _5197 = _5195 ^ _5196;
  wire _5198 = _5194 ^ _5197;
  wire _5199 = _5191 ^ _5198;
  wire _5200 = r899 ^ r987;
  wire _5201 = r1019 ^ r1076;
  wire _5202 = _5200 ^ _5201;
  wire _5203 = r1124 ^ r1228;
  wire _5204 = r1323 ^ r1367;
  wire _5205 = _5203 ^ _5204;
  wire _5206 = _5202 ^ _5205;
  wire _5207 = r1405 ^ r1446;
  wire _5208 = r1575 ^ r1632;
  wire _5209 = _5207 ^ _5208;
  wire _5210 = r1664 ^ r1725;
  wire _5211 = r1919 ^ r1923;
  wire _5212 = _5210 ^ _5211;
  wire _5213 = _5209 ^ _5212;
  wire _5214 = _5206 ^ _5213;
  wire _5215 = _5199 ^ _5214;
  wire _5216 = r19 ^ r79;
  wire _5217 = r115 ^ r254;
  wire _5218 = _5216 ^ _5217;
  wire _5219 = r355 ^ r399;
  wire _5220 = r481 ^ r517;
  wire _5221 = _5219 ^ _5220;
  wire _5222 = _5218 ^ _5221;
  wire _5223 = r581 ^ r668;
  wire _5224 = r734 ^ r865;
  wire _5225 = _5223 ^ _5224;
  wire _5226 = r995 ^ r1047;
  wire _5227 = r1087 ^ r1121;
  wire _5228 = _5226 ^ _5227;
  wire _5229 = _5225 ^ _5228;
  wire _5230 = _5222 ^ _5229;
  wire _5231 = r1381 ^ r1550;
  wire _5232 = r1569 ^ r1637;
  wire _5233 = _5231 ^ _5232;
  wire _5234 = r1663 ^ r1698;
  wire _5235 = r1801 ^ r1874;
  wire _5236 = _5234 ^ _5235;
  wire _5237 = _5233 ^ _5236;
  wire _5238 = r1896 ^ r1907;
  wire _5239 = r1915 ^ r1960;
  wire _5240 = _5238 ^ _5239;
  wire _5241 = r1976 ^ r1979;
  wire _5242 = r2006 ^ r2011;
  wire _5243 = _5241 ^ _5242;
  wire _5244 = _5240 ^ _5243;
  wire _5245 = _5237 ^ _5244;
  wire _5246 = _5230 ^ _5245;
  wire _5247 = _5215 | _5246;
  wire _5248 = _5184 | _5247;
  wire _5249 = r18 ^ r75;
  wire _5250 = r125 ^ r197;
  wire _5251 = _5249 ^ _5250;
  wire _5252 = r260 ^ r375;
  wire _5253 = r401 ^ r539;
  wire _5254 = _5252 ^ _5253;
  wire _5255 = _5251 ^ _5254;
  wire _5256 = r611 ^ r634;
  wire _5257 = r714 ^ r749;
  wire _5258 = _5256 ^ _5257;
  wire _5259 = r792 ^ r833;
  wire _5260 = r924 ^ r967;
  wire _5261 = _5259 ^ _5260;
  wire _5262 = _5258 ^ _5261;
  wire _5263 = _5255 ^ _5262;
  wire _5264 = r1025 ^ r1095;
  wire _5265 = r1139 ^ r1237;
  wire _5266 = _5264 ^ _5265;
  wire _5267 = r1289 ^ r1394;
  wire _5268 = r1494 ^ r1516;
  wire _5269 = _5267 ^ _5268;
  wire _5270 = _5266 ^ _5269;
  wire _5271 = r1557 ^ r1563;
  wire _5272 = r1690 ^ r1732;
  wire _5273 = _5271 ^ _5272;
  wire _5274 = r1826 ^ r1897;
  wire _5275 = r1914 ^ r1916;
  wire _5276 = _5274 ^ _5275;
  wire _5277 = _5273 ^ _5276;
  wire _5278 = _5270 ^ _5277;
  wire _5279 = _5263 ^ _5278;
  wire _5280 = r17 ^ r93;
  wire _5281 = r119 ^ r177;
  wire _5282 = _5280 ^ _5281;
  wire _5283 = r294 ^ r348;
  wire _5284 = r443 ^ r491;
  wire _5285 = _5283 ^ _5284;
  wire _5286 = _5282 ^ _5285;
  wire _5287 = r540 ^ r629;
  wire _5288 = r691 ^ r769;
  wire _5289 = _5287 ^ _5288;
  wire _5290 = r781 ^ r839;
  wire _5291 = r940 ^ r982;
  wire _5292 = _5290 ^ _5291;
  wire _5293 = _5289 ^ _5292;
  wire _5294 = _5286 ^ _5293;
  wire _5295 = r1049 ^ r1070;
  wire _5296 = r1162 ^ r1219;
  wire _5297 = _5295 ^ _5296;
  wire _5298 = r1416 ^ r1440;
  wire _5299 = r1519 ^ r1601;
  wire _5300 = _5298 ^ _5299;
  wire _5301 = _5297 ^ _5300;
  wire _5302 = r1701 ^ r1780;
  wire _5303 = r1806 ^ r1811;
  wire _5304 = _5302 ^ _5303;
  wire _5305 = r1906 ^ r1917;
  wire _5306 = r2018 ^ r2026;
  wire _5307 = _5305 ^ _5306;
  wire _5308 = _5304 ^ _5307;
  wire _5309 = _5301 ^ _5308;
  wire _5310 = _5294 ^ _5309;
  wire _5311 = _5279 | _5310;
  wire _5312 = r16 ^ r57;
  wire _5313 = r122 ^ r210;
  wire _5314 = _5312 ^ _5313;
  wire _5315 = r288 ^ r345;
  wire _5316 = r419 ^ r483;
  wire _5317 = _5315 ^ _5316;
  wire _5318 = _5314 ^ _5317;
  wire _5319 = r667 ^ r683;
  wire _5320 = r723 ^ r777;
  wire _5321 = _5319 ^ _5320;
  wire _5322 = r822 ^ r878;
  wire _5323 = r888 ^ r953;
  wire _5324 = _5322 ^ _5323;
  wire _5325 = _5321 ^ _5324;
  wire _5326 = _5318 ^ _5325;
  wire _5327 = r1007 ^ r1111;
  wire _5328 = r1163 ^ r1309;
  wire _5329 = _5327 ^ _5328;
  wire _5330 = r1356 ^ r1415;
  wire _5331 = r1471 ^ r1515;
  wire _5332 = _5330 ^ _5331;
  wire _5333 = _5329 ^ _5332;
  wire _5334 = r1525 ^ r1579;
  wire _5335 = r1673 ^ r1709;
  wire _5336 = _5334 ^ _5335;
  wire _5337 = r1808 ^ r1862;
  wire _5338 = r1863 ^ r1883;
  wire _5339 = _5337 ^ _5338;
  wire _5340 = _5336 ^ _5339;
  wire _5341 = _5333 ^ _5340;
  wire _5342 = _5326 ^ _5341;
  wire _5343 = r15 ^ r58;
  wire _5344 = r112 ^ r213;
  wire _5345 = _5343 ^ _5344;
  wire _5346 = r225 ^ r292;
  wire _5347 = r360 ^ r471;
  wire _5348 = _5346 ^ _5347;
  wire _5349 = _5345 ^ _5348;
  wire _5350 = r588 ^ r701;
  wire _5351 = r773 ^ r784;
  wire _5352 = _5350 ^ _5351;
  wire _5353 = r880 ^ r990;
  wire _5354 = r1004 ^ r1167;
  wire _5355 = _5353 ^ _5354;
  wire _5356 = _5352 ^ _5355;
  wire _5357 = _5349 ^ _5356;
  wire _5358 = r1214 ^ r1240;
  wire _5359 = r1369 ^ r1393;
  wire _5360 = _5358 ^ _5359;
  wire _5361 = r1502 ^ r1574;
  wire _5362 = r1630 ^ r1665;
  wire _5363 = _5361 ^ _5362;
  wire _5364 = _5360 ^ _5363;
  wire _5365 = r1791 ^ r1895;
  wire _5366 = r1927 ^ r1990;
  wire _5367 = _5365 ^ _5366;
  wire _5368 = r2030 ^ r2035;
  wire _5369 = r2037 ^ r2043;
  wire _5370 = _5368 ^ _5369;
  wire _5371 = _5367 ^ _5370;
  wire _5372 = _5364 ^ _5371;
  wire _5373 = _5357 ^ _5372;
  wire _5374 = _5342 | _5373;
  wire _5375 = _5311 | _5374;
  wire _5376 = _5248 | _5375;
  wire _5377 = r14 ^ r150;
  wire _5378 = r199 ^ r264;
  wire _5379 = _5377 ^ _5378;
  wire _5380 = r283 ^ r353;
  wire _5381 = r409 ^ r487;
  wire _5382 = _5380 ^ _5381;
  wire _5383 = _5379 ^ _5382;
  wire _5384 = r524 ^ r613;
  wire _5385 = r641 ^ r705;
  wire _5386 = _5384 ^ _5385;
  wire _5387 = r724 ^ r801;
  wire _5388 = r851 ^ r943;
  wire _5389 = _5387 ^ _5388;
  wire _5390 = _5386 ^ _5389;
  wire _5391 = _5383 ^ _5390;
  wire _5392 = r955 ^ r1021;
  wire _5393 = r1061 ^ r1130;
  wire _5394 = _5392 ^ _5393;
  wire _5395 = r1196 ^ r1235;
  wire _5396 = r1277 ^ r1325;
  wire _5397 = _5395 ^ _5396;
  wire _5398 = _5394 ^ _5397;
  wire _5399 = r1365 ^ r1603;
  wire _5400 = r1641 ^ r1649;
  wire _5401 = _5399 ^ _5400;
  wire _5402 = r1734 ^ r1786;
  wire _5403 = r1996 ^ r2000;
  wire _5404 = _5402 ^ _5403;
  wire _5405 = _5401 ^ _5404;
  wire _5406 = _5398 ^ _5405;
  wire _5407 = _5391 ^ _5406;
  wire _5408 = r13 ^ r85;
  wire _5409 = r132 ^ r178;
  wire _5410 = _5408 ^ _5409;
  wire _5411 = r266 ^ r316;
  wire _5412 = r387 ^ r395;
  wire _5413 = _5411 ^ _5412;
  wire _5414 = _5410 ^ _5413;
  wire _5415 = r529 ^ r604;
  wire _5416 = r639 ^ r810;
  wire _5417 = _5415 ^ _5416;
  wire _5418 = r831 ^ r938;
  wire _5419 = r969 ^ r1042;
  wire _5420 = _5418 ^ _5419;
  wire _5421 = _5417 ^ _5420;
  wire _5422 = _5414 ^ _5421;
  wire _5423 = r1148 ^ r1203;
  wire _5424 = r1273 ^ r1311;
  wire _5425 = _5423 ^ _5424;
  wire _5426 = r1453 ^ r1469;
  wire _5427 = r1479 ^ r1488;
  wire _5428 = _5426 ^ _5427;
  wire _5429 = _5425 ^ _5428;
  wire _5430 = r1498 ^ r1539;
  wire _5431 = r1713 ^ r1751;
  wire _5432 = _5430 ^ _5431;
  wire _5433 = r1819 ^ r1961;
  wire _5434 = r1962 ^ r1977;
  wire _5435 = _5433 ^ _5434;
  wire _5436 = _5432 ^ _5435;
  wire _5437 = _5429 ^ _5436;
  wire _5438 = _5422 ^ _5437;
  wire _5439 = _5407 | _5438;
  wire _5440 = r12 ^ r101;
  wire _5441 = r145 ^ r236;
  wire _5442 = _5440 ^ _5441;
  wire _5443 = r337 ^ r421;
  wire _5444 = r461 ^ r592;
  wire _5445 = _5443 ^ _5444;
  wire _5446 = _5442 ^ _5445;
  wire _5447 = r620 ^ r843;
  wire _5448 = r965 ^ r1043;
  wire _5449 = _5447 ^ _5448;
  wire _5450 = r1088 ^ r1153;
  wire _5451 = r1171 ^ r1328;
  wire _5452 = _5450 ^ _5451;
  wire _5453 = _5449 ^ _5452;
  wire _5454 = _5446 ^ _5453;
  wire _5455 = r1350 ^ r1417;
  wire _5456 = r1497 ^ r1524;
  wire _5457 = _5455 ^ _5456;
  wire _5458 = r1588 ^ r1626;
  wire _5459 = r1681 ^ r1800;
  wire _5460 = _5458 ^ _5459;
  wire _5461 = _5457 ^ _5460;
  wire _5462 = r1804 ^ r1898;
  wire _5463 = r1924 ^ r1959;
  wire _5464 = _5462 ^ _5463;
  wire _5465 = r1986 ^ r1993;
  wire _5466 = r2020 ^ r2025;
  wire _5467 = _5465 ^ _5466;
  wire _5468 = _5464 ^ _5467;
  wire _5469 = _5461 ^ _5468;
  wire _5470 = _5454 ^ _5469;
  wire _5471 = r105 ^ r156;
  wire _5472 = r222 ^ r311;
  wire _5473 = _5471 ^ _5472;
  wire _5474 = r411 ^ r476;
  wire _5475 = r528 ^ r609;
  wire _5476 = _5474 ^ _5475;
  wire _5477 = _5473 ^ _5476;
  wire _5478 = r699 ^ r743;
  wire _5479 = r811 ^ r852;
  wire _5480 = _5478 ^ _5479;
  wire _5481 = r928 ^ r985;
  wire _5482 = r1084 ^ r1245;
  wire _5483 = _5481 ^ _5482;
  wire _5484 = _5480 ^ _5483;
  wire _5485 = _5477 ^ _5484;
  wire _5486 = r1279 ^ r1294;
  wire _5487 = r1351 ^ r1430;
  wire _5488 = _5486 ^ _5487;
  wire _5489 = r1514 ^ r1518;
  wire _5490 = r1593 ^ r1692;
  wire _5491 = _5489 ^ _5490;
  wire _5492 = _5488 ^ _5491;
  wire _5493 = r1730 ^ r1798;
  wire _5494 = r1857 ^ r1889;
  wire _5495 = _5493 ^ _5494;
  wire _5496 = r1892 ^ r1922;
  wire _5497 = r1933 ^ r1937;
  wire _5498 = _5496 ^ _5497;
  wire _5499 = _5495 ^ _5498;
  wire _5500 = _5492 ^ _5499;
  wire _5501 = _5485 ^ _5500;
  wire _5502 = _5470 | _5501;
  wire _5503 = _5439 | _5502;
  wire _5504 = r11 ^ r110;
  wire _5505 = r126 ^ r229;
  wire _5506 = _5504 ^ _5505;
  wire _5507 = r400 ^ r468;
  wire _5508 = r523 ^ r585;
  wire _5509 = _5507 ^ _5508;
  wire _5510 = _5506 ^ _5509;
  wire _5511 = r655 ^ r727;
  wire _5512 = r879 ^ r894;
  wire _5513 = _5511 ^ _5512;
  wire _5514 = r948 ^ r1013;
  wire _5515 = r1089 ^ r1152;
  wire _5516 = _5514 ^ _5515;
  wire _5517 = _5513 ^ _5516;
  wire _5518 = _5510 ^ _5517;
  wire _5519 = r1201 ^ r1243;
  wire _5520 = r1383 ^ r1414;
  wire _5521 = _5519 ^ _5520;
  wire _5522 = r1591 ^ r1613;
  wire _5523 = r1754 ^ r1795;
  wire _5524 = _5522 ^ _5523;
  wire _5525 = _5521 ^ _5524;
  wire _5526 = r1866 ^ r1875;
  wire _5527 = r1908 ^ r1957;
  wire _5528 = _5526 ^ _5527;
  wire _5529 = r1983 ^ r2009;
  wire _5530 = r2027 ^ r2033;
  wire _5531 = _5529 ^ _5530;
  wire _5532 = _5528 ^ _5531;
  wire _5533 = _5525 ^ _5532;
  wire _5534 = _5518 ^ _5533;
  wire _5535 = r10 ^ r104;
  wire _5536 = r114 ^ r180;
  wire _5537 = _5535 ^ _5536;
  wire _5538 = r237 ^ r295;
  wire _5539 = r384 ^ r417;
  wire _5540 = _5538 ^ _5539;
  wire _5541 = _5537 ^ _5540;
  wire _5542 = r499 ^ r642;
  wire _5543 = r688 ^ r729;
  wire _5544 = _5542 ^ _5543;
  wire _5545 = r825 ^ r838;
  wire _5546 = r892 ^ r949;
  wire _5547 = _5545 ^ _5546;
  wire _5548 = _5544 ^ _5547;
  wire _5549 = _5541 ^ _5548;
  wire _5550 = r1060 ^ r1146;
  wire _5551 = r1183 ^ r1298;
  wire _5552 = _5550 ^ _5551;
  wire _5553 = r1375 ^ r1470;
  wire _5554 = r1522 ^ r1594;
  wire _5555 = _5553 ^ _5554;
  wire _5556 = _5552 ^ _5555;
  wire _5557 = r1682 ^ r1716;
  wire _5558 = r1727 ^ r1820;
  wire _5559 = _5557 ^ _5558;
  wire _5560 = r1829 ^ r1853;
  wire _5561 = r1934 ^ r1944;
  wire _5562 = _5560 ^ _5561;
  wire _5563 = _5559 ^ _5562;
  wire _5564 = _5556 ^ _5563;
  wire _5565 = _5549 ^ _5564;
  wire _5566 = _5534 | _5565;
  wire _5567 = r9 ^ r99;
  wire _5568 = r159 ^ r265;
  wire _5569 = _5567 ^ _5568;
  wire _5570 = r361 ^ r453;
  wire _5571 = r514 ^ r597;
  wire _5572 = _5570 ^ _5571;
  wire _5573 = _5569 ^ _5572;
  wire _5574 = r753 ^ r984;
  wire _5575 = r1033 ^ r1100;
  wire _5576 = _5574 ^ _5575;
  wire _5577 = r1128 ^ r1168;
  wire _5578 = r1257 ^ r1302;
  wire _5579 = _5577 ^ _5578;
  wire _5580 = _5576 ^ _5579;
  wire _5581 = _5573 ^ _5580;
  wire _5582 = r1336 ^ r1425;
  wire _5583 = r1614 ^ r1671;
  wire _5584 = _5582 ^ _5583;
  wire _5585 = r1736 ^ r1770;
  wire _5586 = r1799 ^ r1849;
  wire _5587 = _5585 ^ _5586;
  wire _5588 = _5584 ^ _5587;
  wire _5589 = r1877 ^ r1887;
  wire _5590 = r1904 ^ r1966;
  wire _5591 = _5589 ^ _5590;
  wire _5592 = r1970 ^ r1988;
  wire _5593 = r1992 ^ r1995;
  wire _5594 = _5592 ^ _5593;
  wire _5595 = _5591 ^ _5594;
  wire _5596 = _5588 ^ _5595;
  wire _5597 = _5581 ^ _5596;
  wire _5598 = r8 ^ r82;
  wire _5599 = r117 ^ r211;
  wire _5600 = _5598 ^ _5599;
  wire _5601 = r278 ^ r325;
  wire _5602 = r344 ^ r445;
  wire _5603 = _5601 ^ _5602;
  wire _5604 = _5600 ^ _5603;
  wire _5605 = r503 ^ r535;
  wire _5606 = r590 ^ r638;
  wire _5607 = _5605 ^ _5606;
  wire _5608 = r709 ^ r735;
  wire _5609 = r815 ^ r846;
  wire _5610 = _5608 ^ _5609;
  wire _5611 = _5607 ^ _5610;
  wire _5612 = _5604 ^ _5611;
  wire _5613 = r908 ^ r976;
  wire _5614 = r1106 ^ r1135;
  wire _5615 = _5613 ^ _5614;
  wire _5616 = r1164 ^ r1172;
  wire _5617 = r1260 ^ r1293;
  wire _5618 = _5616 ^ _5617;
  wire _5619 = _5615 ^ _5618;
  wire _5620 = r1340 ^ r1395;
  wire _5621 = r1438 ^ r1495;
  wire _5622 = _5620 ^ _5621;
  wire _5623 = r1505 ^ r1606;
  wire _5624 = r1627 ^ r1764;
  wire _5625 = _5623 ^ _5624;
  wire _5626 = _5622 ^ _5625;
  wire _5627 = _5619 ^ _5626;
  wire _5628 = _5612 ^ _5627;
  wire _5629 = _5597 | _5628;
  wire _5630 = _5566 | _5629;
  wire _5631 = _5503 | _5630;
  wire _5632 = _5376 | _5631;
  wire _5633 = r7 ^ r89;
  wire _5634 = r137 ^ r176;
  wire _5635 = _5633 ^ _5634;
  wire _5636 = r251 ^ r286;
  wire _5637 = r356 ^ r404;
  wire _5638 = _5636 ^ _5637;
  wire _5639 = _5635 ^ _5638;
  wire _5640 = r450 ^ r533;
  wire _5641 = r566 ^ r664;
  wire _5642 = _5640 ^ _5641;
  wire _5643 = r686 ^ r746;
  wire _5644 = r817 ^ r867;
  wire _5645 = _5643 ^ _5644;
  wire _5646 = _5642 ^ _5645;
  wire _5647 = _5639 ^ _5646;
  wire _5648 = r910 ^ r993;
  wire _5649 = r1032 ^ r1091;
  wire _5650 = _5648 ^ _5649;
  wire _5651 = r1158 ^ r1169;
  wire _5652 = r1202 ^ r1246;
  wire _5653 = _5651 ^ _5652;
  wire _5654 = _5650 ^ _5653;
  wire _5655 = r1313 ^ r1389;
  wire _5656 = r1464 ^ r1536;
  wire _5657 = _5655 ^ _5656;
  wire _5658 = r1549 ^ r1625;
  wire _5659 = r1691 ^ r1765;
  wire _5660 = _5658 ^ _5659;
  wire _5661 = _5657 ^ _5660;
  wire _5662 = _5654 ^ _5661;
  wire _5663 = _5647 ^ _5662;
  wire _5664 = r6 ^ r109;
  wire _5665 = r147 ^ r204;
  wire _5666 = _5664 ^ _5665;
  wire _5667 = r232 ^ r304;
  wire _5668 = r368 ^ r397;
  wire _5669 = _5667 ^ _5668;
  wire _5670 = _5666 ^ _5669;
  wire _5671 = r496 ^ r512;
  wire _5672 = r576 ^ r651;
  wire _5673 = _5671 ^ _5672;
  wire _5674 = r721 ^ r754;
  wire _5675 = r787 ^ r881;
  wire _5676 = _5674 ^ _5675;
  wire _5677 = _5673 ^ _5676;
  wire _5678 = _5670 ^ _5677;
  wire _5679 = r895 ^ r998;
  wire _5680 = r1027 ^ r1059;
  wire _5681 = _5679 ^ _5680;
  wire _5682 = r1093 ^ r1156;
  wire _5683 = r1320 ^ r1339;
  wire _5684 = _5682 ^ _5683;
  wire _5685 = _5681 ^ _5684;
  wire _5686 = r1472 ^ r1517;
  wire _5687 = r1523 ^ r1538;
  wire _5688 = _5686 ^ _5687;
  wire _5689 = r1597 ^ r1639;
  wire _5690 = r1697 ^ r1766;
  wire _5691 = _5689 ^ _5690;
  wire _5692 = _5688 ^ _5691;
  wire _5693 = _5685 ^ _5692;
  wire _5694 = _5678 ^ _5693;
  wire _5695 = _5663 | _5694;
  wire _5696 = r5 ^ r107;
  wire _5697 = r142 ^ r201;
  wire _5698 = _5696 ^ _5697;
  wire _5699 = r313 ^ r338;
  wire _5700 = r428 ^ r549;
  wire _5701 = _5699 ^ _5700;
  wire _5702 = _5698 ^ _5701;
  wire _5703 = r621 ^ r728;
  wire _5704 = r823 ^ r877;
  wire _5705 = _5703 ^ _5704;
  wire _5706 = r927 ^ r1010;
  wire _5707 = r1065 ^ r1133;
  wire _5708 = _5706 ^ _5707;
  wire _5709 = _5705 ^ _5708;
  wire _5710 = _5702 ^ _5709;
  wire _5711 = r1193 ^ r1242;
  wire _5712 = r1282 ^ r1304;
  wire _5713 = _5711 ^ _5712;
  wire _5714 = r1503 ^ r1599;
  wire _5715 = r1609 ^ r1676;
  wire _5716 = _5714 ^ _5715;
  wire _5717 = _5713 ^ _5716;
  wire _5718 = r1704 ^ r1796;
  wire _5719 = r1813 ^ r1871;
  wire _5720 = _5718 ^ _5719;
  wire _5721 = r1888 ^ r1920;
  wire _5722 = r1963 ^ r1978;
  wire _5723 = _5721 ^ _5722;
  wire _5724 = _5720 ^ _5723;
  wire _5725 = _5717 ^ _5724;
  wire _5726 = _5710 ^ _5725;
  wire _5727 = r4 ^ r87;
  wire _5728 = r148 ^ r215;
  wire _5729 = _5727 ^ _5728;
  wire _5730 = r267 ^ r308;
  wire _5731 = r386 ^ r438;
  wire _5732 = _5730 ^ _5731;
  wire _5733 = _5729 ^ _5732;
  wire _5734 = r460 ^ r552;
  wire _5735 = r573 ^ r666;
  wire _5736 = _5734 ^ _5735;
  wire _5737 = r711 ^ r742;
  wire _5738 = r780 ^ r841;
  wire _5739 = _5737 ^ _5738;
  wire _5740 = _5736 ^ _5739;
  wire _5741 = _5733 ^ _5740;
  wire _5742 = r891 ^ r997;
  wire _5743 = r1017 ^ r1098;
  wire _5744 = _5742 ^ _5743;
  wire _5745 = r1114 ^ r1179;
  wire _5746 = r1270 ^ r1306;
  wire _5747 = _5745 ^ _5746;
  wire _5748 = _5744 ^ _5747;
  wire _5749 = r1372 ^ r1428;
  wire _5750 = r1483 ^ r1610;
  wire _5751 = _5749 ^ _5750;
  wire _5752 = r1670 ^ r1717;
  wire _5753 = r1771 ^ r1841;
  wire _5754 = _5752 ^ _5753;
  wire _5755 = _5751 ^ _5754;
  wire _5756 = _5748 ^ _5755;
  wire _5757 = _5741 ^ _5756;
  wire _5758 = _5726 | _5757;
  wire _5759 = _5695 | _5758;
  wire _5760 = r67 ^ r208;
  wire _5761 = r263 ^ r314;
  wire _5762 = _5760 ^ _5761;
  wire _5763 = r371 ^ r432;
  wire _5764 = r472 ^ r536;
  wire _5765 = _5763 ^ _5764;
  wire _5766 = _5762 ^ _5765;
  wire _5767 = r563 ^ r687;
  wire _5768 = r770 ^ r788;
  wire _5769 = _5767 ^ _5768;
  wire _5770 = r863 ^ r919;
  wire _5771 = r1038 ^ r1116;
  wire _5772 = _5770 ^ _5771;
  wire _5773 = _5769 ^ _5772;
  wire _5774 = _5766 ^ _5773;
  wire _5775 = r1204 ^ r1221;
  wire _5776 = r1379 ^ r1419;
  wire _5777 = _5775 ^ _5776;
  wire _5778 = r1468 ^ r1507;
  wire _5779 = r1529 ^ r1604;
  wire _5780 = _5778 ^ _5779;
  wire _5781 = _5777 ^ _5780;
  wire _5782 = r1638 ^ r1695;
  wire _5783 = r1738 ^ r1885;
  wire _5784 = _5782 ^ _5783;
  wire _5785 = r1901 ^ r1935;
  wire _5786 = r2016 ^ r2024;
  wire _5787 = _5785 ^ _5786;
  wire _5788 = _5784 ^ _5787;
  wire _5789 = _5781 ^ _5788;
  wire _5790 = _5774 ^ _5789;
  wire _5791 = r3 ^ r70;
  wire _5792 = r162 ^ r186;
  wire _5793 = _5791 ^ _5792;
  wire _5794 = r227 ^ r303;
  wire _5795 = r389 ^ r436;
  wire _5796 = _5794 ^ _5795;
  wire _5797 = _5793 ^ _5796;
  wire _5798 = r482 ^ r513;
  wire _5799 = r598 ^ r619;
  wire _5800 = _5798 ^ _5799;
  wire _5801 = r708 ^ r816;
  wire _5802 = r864 ^ r904;
  wire _5803 = _5801 ^ _5802;
  wire _5804 = _5800 ^ _5803;
  wire _5805 = _5797 ^ _5804;
  wire _5806 = r973 ^ r1036;
  wire _5807 = r1066 ^ r1159;
  wire _5808 = _5806 ^ _5807;
  wire _5809 = r1195 ^ r1223;
  wire _5810 = r1225 ^ r1312;
  wire _5811 = _5809 ^ _5810;
  wire _5812 = _5808 ^ _5811;
  wire _5813 = r1346 ^ r1385;
  wire _5814 = r1476 ^ r1541;
  wire _5815 = _5813 ^ _5814;
  wire _5816 = r1631 ^ r1710;
  wire _5817 = r1733 ^ r1842;
  wire _5818 = _5816 ^ _5817;
  wire _5819 = _5815 ^ _5818;
  wire _5820 = _5812 ^ _5819;
  wire _5821 = _5805 ^ _5820;
  wire _5822 = _5790 | _5821;
  wire _5823 = r2 ^ r54;
  wire _5824 = r169 ^ r195;
  wire _5825 = _5823 ^ _5824;
  wire _5826 = r248 ^ r328;
  wire _5827 = r350 ^ r425;
  wire _5828 = _5826 ^ _5827;
  wire _5829 = _5825 ^ _5828;
  wire _5830 = r454 ^ r532;
  wire _5831 = r582 ^ r647;
  wire _5832 = _5830 ^ _5831;
  wire _5833 = r678 ^ r772;
  wire _5834 = r829 ^ r840;
  wire _5835 = _5833 ^ _5834;
  wire _5836 = _5832 ^ _5835;
  wire _5837 = _5829 ^ _5836;
  wire _5838 = r929 ^ r1015;
  wire _5839 = r1092 ^ r1134;
  wire _5840 = _5838 ^ _5839;
  wire _5841 = r1184 ^ r1272;
  wire _5842 = r1324 ^ r1334;
  wire _5843 = _5841 ^ _5842;
  wire _5844 = _5840 ^ _5843;
  wire _5845 = r1344 ^ r1448;
  wire _5846 = r1486 ^ r1647;
  wire _5847 = _5845 ^ _5846;
  wire _5848 = r1656 ^ r1700;
  wire _5849 = r1772 ^ r1843;
  wire _5850 = _5848 ^ _5849;
  wire _5851 = _5847 ^ _5850;
  wire _5852 = _5844 ^ _5851;
  wire _5853 = _5837 ^ _5852;
  wire _5854 = r1 ^ r88;
  wire _5855 = r190 ^ r281;
  wire _5856 = _5854 ^ _5855;
  wire _5857 = r358 ^ r405;
  wire _5858 = r498 ^ r560;
  wire _5859 = _5857 ^ _5858;
  wire _5860 = _5856 ^ _5859;
  wire _5861 = r593 ^ r644;
  wire _5862 = r718 ^ r730;
  wire _5863 = _5861 ^ _5862;
  wire _5864 = r802 ^ r832;
  wire _5865 = r921 ^ r944;
  wire _5866 = _5864 ^ _5865;
  wire _5867 = _5863 ^ _5866;
  wire _5868 = _5860 ^ _5867;
  wire _5869 = r1052 ^ r1105;
  wire _5870 = r1155 ^ r1200;
  wire _5871 = _5869 ^ _5870;
  wire _5872 = r1258 ^ r1280;
  wire _5873 = r1402 ^ r1432;
  wire _5874 = _5872 ^ _5873;
  wire _5875 = _5871 ^ _5874;
  wire _5876 = r1491 ^ r1530;
  wire _5877 = r1598 ^ r1659;
  wire _5878 = _5876 ^ _5877;
  wire _5879 = r1776 ^ r1860;
  wire _5880 = r1926 ^ r1931;
  wire _5881 = _5879 ^ _5880;
  wire _5882 = _5878 ^ _5881;
  wire _5883 = _5875 ^ _5882;
  wire _5884 = _5868 ^ _5883;
  wire _5885 = _5853 | _5884;
  wire _5886 = _5822 | _5885;
  wire _5887 = _5759 | _5886;
  wire _5888 = r0 ^ r106;
  wire _5889 = r153 ^ r193;
  wire _5890 = _5888 ^ _5889;
  wire _5891 = r226 ^ r318;
  wire _5892 = r354 ^ r444;
  wire _5893 = _5891 ^ _5892;
  wire _5894 = _5890 ^ _5893;
  wire _5895 = r484 ^ r545;
  wire _5896 = r603 ^ r658;
  wire _5897 = _5895 ^ _5896;
  wire _5898 = r689 ^ r726;
  wire _5899 = r783 ^ r850;
  wire _5900 = _5898 ^ _5899;
  wire _5901 = _5897 ^ _5900;
  wire _5902 = _5894 ^ _5901;
  wire _5903 = r909 ^ r1001;
  wire _5904 = r1055 ^ r1080;
  wire _5905 = _5903 ^ _5904;
  wire _5906 = r1125 ^ r1176;
  wire _5907 = r1305 ^ r1358;
  wire _5908 = _5906 ^ _5907;
  wire _5909 = _5905 ^ _5908;
  wire _5910 = r1412 ^ r1426;
  wire _5911 = r1463 ^ r1521;
  wire _5912 = _5910 ^ _5911;
  wire _5913 = r1558 ^ r1648;
  wire _5914 = r1652 ^ r1767;
  wire _5915 = _5913 ^ _5914;
  wire _5916 = _5912 ^ _5915;
  wire _5917 = _5909 ^ _5916;
  wire _5918 = _5902 ^ _5917;
  wire _5919 = r121 ^ r272;
  wire _5920 = r320 ^ r359;
  wire _5921 = _5919 ^ _5920;
  wire _5922 = r501 ^ r577;
  wire _5923 = r680 ^ r804;
  wire _5924 = _5922 ^ _5923;
  wire _5925 = _5921 ^ _5924;
  wire _5926 = r926 ^ r979;
  wire _5927 = r1039 ^ r1174;
  wire _5928 = _5926 ^ _5927;
  wire _5929 = r1251 ^ r1319;
  wire _5930 = r1361 ^ r1406;
  wire _5931 = _5929 ^ _5930;
  wire _5932 = _5928 ^ _5931;
  wire _5933 = _5925 ^ _5932;
  wire _5934 = r1449 ^ r1490;
  wire _5935 = r1561 ^ r1677;
  wire _5936 = _5934 ^ _5935;
  wire _5937 = r1715 ^ r1723;
  wire _5938 = r1865 ^ r1876;
  wire _5939 = _5937 ^ _5938;
  wire _5940 = _5936 ^ _5939;
  wire _5941 = r1903 ^ r1943;
  wire _5942 = r1954 ^ r1981;
  wire _5943 = _5941 ^ _5942;
  wire _5944 = r2007 ^ r2012;
  wire _5945 = r2028 ^ r2036;
  wire _5946 = _5944 ^ _5945;
  wire _5947 = _5943 ^ _5946;
  wire _5948 = _5940 ^ _5947;
  wire _5949 = _5933 ^ _5948;
  wire _5950 = _5918 | _5949;
  wire _5951 = r63 ^ r160;
  wire _5952 = r216 ^ r235;
  wire _5953 = _5951 ^ _5952;
  wire _5954 = r290 ^ r349;
  wire _5955 = r410 ^ r465;
  wire _5956 = _5954 ^ _5955;
  wire _5957 = _5953 ^ _5956;
  wire _5958 = r507 ^ r565;
  wire _5959 = r627 ^ r669;
  wire _5960 = _5958 ^ _5959;
  wire _5961 = r766 ^ r818;
  wire _5962 = r900 ^ r958;
  wire _5963 = _5961 ^ _5962;
  wire _5964 = _5960 ^ _5963;
  wire _5965 = _5957 ^ _5964;
  wire _5966 = r1016 ^ r1082;
  wire _5967 = r1136 ^ r1188;
  wire _5968 = _5966 ^ _5967;
  wire _5969 = r1222 ^ r1248;
  wire _5970 = r1295 ^ r1347;
  wire _5971 = _5969 ^ _5970;
  wire _5972 = _5968 ^ _5971;
  wire _5973 = r1410 ^ r1478;
  wire _5974 = r1501 ^ r1571;
  wire _5975 = _5973 ^ _5974;
  wire _5976 = r1645 ^ r1666;
  wire _5977 = r1928 ^ r1932;
  wire _5978 = _5976 ^ _5977;
  wire _5979 = _5975 ^ _5978;
  wire _5980 = _5972 ^ _5979;
  wire _5981 = _5965 ^ _5980;
  wire _5982 = r90 ^ r113;
  wire _5983 = r200 ^ r240;
  wire _5984 = _5982 ^ _5983;
  wire _5985 = r326 ^ r374;
  wire _5986 = r439 ^ r474;
  wire _5987 = _5985 ^ _5986;
  wire _5988 = _5984 ^ _5987;
  wire _5989 = r550 ^ r606;
  wire _5990 = r636 ^ r685;
  wire _5991 = _5989 ^ _5990;
  wire _5992 = r767 ^ r814;
  wire _5993 = r854 ^ r897;
  wire _5994 = _5992 ^ _5993;
  wire _5995 = _5991 ^ _5994;
  wire _5996 = _5988 ^ _5995;
  wire _5997 = r961 ^ r1035;
  wire _5998 = r1094 ^ r1127;
  wire _5999 = _5997 ^ _5998;
  wire _6000 = r1181 ^ r1263;
  wire _6001 = r1327 ^ r1378;
  wire _6002 = _6000 ^ _6001;
  wire _6003 = _5999 ^ _6002;
  wire _6004 = r1399 ^ r1554;
  wire _6005 = r1564 ^ r1590;
  wire _6006 = _6004 ^ _6005;
  wire _6007 = r1629 ^ r1672;
  wire _6008 = r1722 ^ r1768;
  wire _6009 = _6007 ^ _6008;
  wire _6010 = _6006 ^ _6009;
  wire _6011 = _6003 ^ _6010;
  wire _6012 = _5996 ^ _6011;
  wire _6013 = _5981 | _6012;
  wire _6014 = _5950 | _6013;
  wire _6015 = r81 ^ r212;
  wire _6016 = r279 ^ r284;
  wire _6017 = _6015 ^ _6016;
  wire _6018 = r381 ^ r427;
  wire _6019 = r469 ^ r511;
  wire _6020 = _6018 ^ _6019;
  wire _6021 = _6017 ^ _6020;
  wire _6022 = r568 ^ r715;
  wire _6023 = r744 ^ r779;
  wire _6024 = _6022 ^ _6023;
  wire _6025 = r848 ^ r913;
  wire _6026 = r945 ^ r1090;
  wire _6027 = _6025 ^ _6026;
  wire _6028 = _6024 ^ _6027;
  wire _6029 = _6021 ^ _6028;
  wire _6030 = r1108 ^ r1212;
  wire _6031 = r1256 ^ r1343;
  wire _6032 = _6030 ^ _6031;
  wire _6033 = r1542 ^ r1568;
  wire _6034 = r1721 ^ r1737;
  wire _6035 = _6033 ^ _6034;
  wire _6036 = _6032 ^ _6035;
  wire _6037 = r1774 ^ r1783;
  wire _6038 = r1812 ^ r1825;
  wire _6039 = _6037 ^ _6038;
  wire _6040 = r1828 ^ r1852;
  wire _6041 = r1870 ^ r1884;
  wire _6042 = _6040 ^ _6041;
  wire _6043 = _6039 ^ _6042;
  wire _6044 = _6036 ^ _6043;
  wire _6045 = _6029 ^ _6044;
  wire _6046 = r68 ^ r152;
  wire _6047 = r223 ^ r239;
  wire _6048 = _6046 ^ _6047;
  wire _6049 = r291 ^ r363;
  wire _6050 = r413 ^ r475;
  wire _6051 = _6049 ^ _6050;
  wire _6052 = _6048 ^ _6051;
  wire _6053 = r541 ^ r587;
  wire _6054 = r633 ^ r713;
  wire _6055 = _6053 ^ _6054;
  wire _6056 = r736 ^ r799;
  wire _6057 = r885 ^ r906;
  wire _6058 = _6056 ^ _6057;
  wire _6059 = _6055 ^ _6058;
  wire _6060 = _6052 ^ _6059;
  wire _6061 = r980 ^ r1048;
  wire _6062 = r1132 ^ r1233;
  wire _6063 = _6061 ^ _6062;
  wire _6064 = r1307 ^ r1418;
  wire _6065 = r1444 ^ r1506;
  wire _6066 = _6064 ^ _6065;
  wire _6067 = _6063 ^ _6066;
  wire _6068 = r1559 ^ r1596;
  wire _6069 = r1662 ^ r1719;
  wire _6070 = _6068 ^ _6069;
  wire _6071 = r1740 ^ r1748;
  wire _6072 = r1793 ^ r1844;
  wire _6073 = _6071 ^ _6072;
  wire _6074 = _6070 ^ _6073;
  wire _6075 = _6067 ^ _6074;
  wire _6076 = _6060 ^ _6075;
  wire _6077 = _6045 | _6076;
  wire _6078 = r168 ^ r196;
  wire _6079 = r234 ^ r319;
  wire _6080 = _6078 ^ _6079;
  wire _6081 = r365 ^ r430;
  wire _6082 = r464 ^ r538;
  wire _6083 = _6081 ^ _6082;
  wire _6084 = _6080 ^ _6083;
  wire _6085 = r595 ^ r673;
  wire _6086 = r752 ^ r836;
  wire _6087 = _6085 ^ _6086;
  wire _6088 = r935 ^ r1000;
  wire _6089 = r1018 ^ r1112;
  wire _6090 = _6088 ^ _6089;
  wire _6091 = _6087 ^ _6090;
  wire _6092 = _6084 ^ _6091;
  wire _6093 = r1241 ^ r1355;
  wire _6094 = r1433 ^ r1466;
  wire _6095 = _6093 ^ _6094;
  wire _6096 = r1485 ^ r1653;
  wire _6097 = r1720 ^ r1753;
  wire _6098 = _6096 ^ _6097;
  wire _6099 = _6095 ^ _6098;
  wire _6100 = r1782 ^ r1821;
  wire _6101 = r1905 ^ r1968;
  wire _6102 = _6100 ^ _6101;
  wire _6103 = r2002 ^ r2004;
  wire _6104 = r2038 ^ r2040;
  wire _6105 = _6103 ^ _6104;
  wire _6106 = _6102 ^ _6105;
  wire _6107 = _6099 ^ _6106;
  wire _6108 = _6092 ^ _6107;
  wire _6109 = r52 ^ r59;
  wire _6110 = r138 ^ r185;
  wire _6111 = _6109 ^ _6110;
  wire _6112 = r270 ^ r280;
  wire _6113 = r393 ^ r486;
  wire _6114 = _6112 ^ _6113;
  wire _6115 = _6111 ^ _6114;
  wire _6116 = r554 ^ r591;
  wire _6117 = r659 ^ r719;
  wire _6118 = _6116 ^ _6117;
  wire _6119 = r757 ^ r778;
  wire _6120 = r859 ^ r889;
  wire _6121 = _6119 ^ _6120;
  wire _6122 = _6118 ^ _6121;
  wire _6123 = _6115 ^ _6122;
  wire _6124 = r970 ^ r1009;
  wire _6125 = r1078 ^ r1161;
  wire _6126 = _6124 ^ _6125;
  wire _6127 = r1217 ^ r1224;
  wire _6128 = r1236 ^ r1322;
  wire _6129 = _6127 ^ _6128;
  wire _6130 = _6126 ^ _6129;
  wire _6131 = r1333 ^ r1380;
  wire _6132 = r1548 ^ r1585;
  wire _6133 = _6131 ^ _6132;
  wire _6134 = r1634 ^ r1684;
  wire _6135 = r1703 ^ r1769;
  wire _6136 = _6134 ^ _6135;
  wire _6137 = _6133 ^ _6136;
  wire _6138 = _6130 ^ _6137;
  wire _6139 = _6123 ^ _6138;
  wire _6140 = _6108 | _6139;
  wire _6141 = _6077 | _6140;
  wire _6142 = _6014 | _6141;
  wire _6143 = _5887 | _6142;
  wire _6144 = _5632 | _6143;
  wire _6145 = _5121 | _6144;
  wire _6146 = r53 ^ r107;
  wire _6147 = r128 ^ r197;
  wire _6148 = _6146 ^ _6147;
  wire _6149 = r243 ^ r297;
  wire _6150 = r340 ^ r440;
  wire _6151 = _6149 ^ _6150;
  wire _6152 = _6148 ^ _6151;
  wire _6153 = r456 ^ r533;
  wire _6154 = r578 ^ r639;
  wire _6155 = _6153 ^ _6154;
  wire _6156 = r709 ^ r761;
  wire _6157 = r794 ^ r857;
  wire _6158 = _6156 ^ _6157;
  wire _6159 = _6155 ^ _6158;
  wire _6160 = _6152 ^ _6159;
  wire _6161 = r892 ^ r1001;
  wire _6162 = r1036 ^ r1072;
  wire _6163 = _6161 ^ _6162;
  wire _6164 = r1156 ^ r1243;
  wire _6165 = r1344 ^ r1415;
  wire _6166 = _6164 ^ _6165;
  wire _6167 = _6163 ^ _6166;
  wire _6168 = r1455 ^ r1485;
  wire _6169 = r1518 ^ r1580;
  wire _6170 = _6168 ^ _6169;
  wire _6171 = r1663 ^ r1734;
  wire _6172 = r1788 ^ r1845;
  wire _6173 = _6171 ^ _6172;
  wire _6174 = _6170 ^ _6173;
  wire _6175 = _6167 ^ _6174;
  wire _6176 = _6160 ^ _6175;
  wire _6177 = r51 ^ r58;
  wire _6178 = r137 ^ r269;
  wire _6179 = _6177 ^ _6178;
  wire _6180 = r333 ^ r485;
  wire _6181 = r590 ^ r658;
  wire _6182 = _6180 ^ _6181;
  wire _6183 = _6179 ^ _6182;
  wire _6184 = r756 ^ r858;
  wire _6185 = r888 ^ r969;
  wire _6186 = _6184 ^ _6185;
  wire _6187 = r1008 ^ r1160;
  wire _6188 = r1216 ^ r1223;
  wire _6189 = _6187 ^ _6188;
  wire _6190 = _6186 ^ _6189;
  wire _6191 = _6183 ^ _6190;
  wire _6192 = r1235 ^ r1321;
  wire _6193 = r1379 ^ r1584;
  wire _6194 = _6192 ^ _6193;
  wire _6195 = r1633 ^ r1683;
  wire _6196 = r1702 ^ r1877;
  wire _6197 = _6195 ^ _6196;
  wire _6198 = _6194 ^ _6197;
  wire _6199 = r1899 ^ r1944;
  wire _6200 = r1985 ^ r2022;
  wire _6201 = _6199 ^ _6200;
  wire _6202 = r2027 ^ r2032;
  wire _6203 = r2040 ^ r2042;
  wire _6204 = _6202 ^ _6203;
  wire _6205 = _6201 ^ _6204;
  wire _6206 = _6198 ^ _6205;
  wire _6207 = _6191 ^ _6206;
  wire _6208 = _6176 | _6207;
  wire _6209 = r50 ^ r55;
  wire _6210 = r115 ^ r171;
  wire _6211 = _6209 ^ _6210;
  wire _6212 = r275 ^ r304;
  wire _6213 = r371 ^ r401;
  wire _6214 = _6212 ^ _6213;
  wire _6215 = _6211 ^ _6214;
  wire _6216 = r492 ^ r546;
  wire _6217 = r595 ^ r642;
  wire _6218 = _6216 ^ _6217;
  wire _6219 = r695 ^ r823;
  wire _6220 = r938 ^ r953;
  wire _6221 = _6219 ^ _6220;
  wire _6222 = _6218 ^ _6221;
  wire _6223 = _6215 ^ _6222;
  wire _6224 = r1052 ^ r1106;
  wire _6225 = r1118 ^ r1208;
  wire _6226 = _6224 ^ _6225;
  wire _6227 = r1219 ^ r1239;
  wire _6228 = r1290 ^ r1370;
  wire _6229 = _6227 ^ _6228;
  wire _6230 = _6226 ^ _6229;
  wire _6231 = r1412 ^ r1428;
  wire _6232 = r1499 ^ r1585;
  wire _6233 = _6231 ^ _6232;
  wire _6234 = r1616 ^ r1654;
  wire _6235 = r1792 ^ r1846;
  wire _6236 = _6234 ^ _6235;
  wire _6237 = _6233 ^ _6236;
  wire _6238 = _6230 ^ _6237;
  wire _6239 = _6223 ^ _6238;
  wire _6240 = r72 ^ r139;
  wire _6241 = r187 ^ r244;
  wire _6242 = _6240 ^ _6241;
  wire _6243 = r384 ^ r397;
  wire _6244 = r519 ^ r585;
  wire _6245 = _6243 ^ _6244;
  wire _6246 = _6242 ^ _6245;
  wire _6247 = r705 ^ r755;
  wire _6248 = r785 ^ r834;
  wire _6249 = _6247 ^ _6248;
  wire _6250 = r942 ^ r1098;
  wire _6251 = r1188 ^ r1229;
  wire _6252 = _6250 ^ _6251;
  wire _6253 = _6249 ^ _6252;
  wire _6254 = _6246 ^ _6253;
  wire _6255 = r1291 ^ r1358;
  wire _6256 = r1400 ^ r1438;
  wire _6257 = _6255 ^ _6256;
  wire _6258 = r1464 ^ r1555;
  wire _6259 = r1619 ^ r1668;
  wire _6260 = _6258 ^ _6259;
  wire _6261 = _6257 ^ _6260;
  wire _6262 = r1718 ^ r1729;
  wire _6263 = r1732 ^ r1790;
  wire _6264 = _6262 ^ _6263;
  wire _6265 = r1827 ^ r1833;
  wire _6266 = r1843 ^ r1885;
  wire _6267 = _6265 ^ _6266;
  wire _6268 = _6264 ^ _6267;
  wire _6269 = _6261 ^ _6268;
  wire _6270 = _6254 ^ _6269;
  wire _6271 = _6239 | _6270;
  wire _6272 = _6208 | _6271;
  wire _6273 = r49 ^ r64;
  wire _6274 = r153 ^ r205;
  wire _6275 = _6273 ^ _6274;
  wire _6276 = r242 ^ r306;
  wire _6277 = r402 ^ r478;
  wire _6278 = _6276 ^ _6277;
  wire _6279 = _6275 ^ _6278;
  wire _6280 = r529 ^ r664;
  wire _6281 = r699 ^ r749;
  wire _6282 = _6280 ^ _6281;
  wire _6283 = r790 ^ r830;
  wire _6284 = r869 ^ r931;
  wire _6285 = _6283 ^ _6284;
  wire _6286 = _6282 ^ _6285;
  wire _6287 = _6279 ^ _6286;
  wire _6288 = r971 ^ r1043;
  wire _6289 = r1063 ^ r1142;
  wire _6290 = _6288 ^ _6289;
  wire _6291 = r1172 ^ r1263;
  wire _6292 = r1320 ^ r1376;
  wire _6293 = _6291 ^ _6292;
  wire _6294 = _6290 ^ _6293;
  wire _6295 = r1550 ^ r1571;
  wire _6296 = r1604 ^ r1673;
  wire _6297 = _6295 ^ _6296;
  wire _6298 = r1728 ^ r1740;
  wire _6299 = r1769 ^ r1847;
  wire _6300 = _6298 ^ _6299;
  wire _6301 = _6297 ^ _6300;
  wire _6302 = _6294 ^ _6301;
  wire _6303 = _6287 ^ _6302;
  wire _6304 = r48 ^ r96;
  wire _6305 = r150 ^ r213;
  wire _6306 = _6304 ^ _6305;
  wire _6307 = r273 ^ r320;
  wire _6308 = r363 ^ r504;
  wire _6309 = _6307 ^ _6308;
  wire _6310 = _6306 ^ _6309;
  wire _6311 = r523 ^ r614;
  wire _6312 = r636 ^ r703;
  wire _6313 = _6311 ^ _6312;
  wire _6314 = r732 ^ r872;
  wire _6315 = r887 ^ r913;
  wire _6316 = _6314 ^ _6315;
  wire _6317 = _6313 ^ _6316;
  wire _6318 = _6310 ^ _6317;
  wire _6319 = r958 ^ r1040;
  wire _6320 = r1068 ^ r1153;
  wire _6321 = _6319 ^ _6320;
  wire _6322 = r1184 ^ r1246;
  wire _6323 = r1312 ^ r1351;
  wire _6324 = _6322 ^ _6323;
  wire _6325 = _6321 ^ _6324;
  wire _6326 = r1403 ^ r1457;
  wire _6327 = r1481 ^ r1500;
  wire _6328 = _6326 ^ _6327;
  wire _6329 = r1634 ^ r1670;
  wire _6330 = r1701 ^ r1770;
  wire _6331 = _6329 ^ _6330;
  wire _6332 = _6328 ^ _6331;
  wire _6333 = _6325 ^ _6332;
  wire _6334 = _6318 ^ _6333;
  wire _6335 = _6303 | _6334;
  wire _6336 = r47 ^ r105;
  wire _6337 = r111 ^ r208;
  wire _6338 = _6336 ^ _6337;
  wire _6339 = r254 ^ r316;
  wire _6340 = r379 ^ r415;
  wire _6341 = _6339 ^ _6340;
  wire _6342 = _6338 ^ _6341;
  wire _6343 = r484 ^ r526;
  wire _6344 = r599 ^ r625;
  wire _6345 = _6343 ^ _6344;
  wire _6346 = r692 ^ r739;
  wire _6347 = r789 ^ r859;
  wire _6348 = _6346 ^ _6347;
  wire _6349 = _6345 ^ _6348;
  wire _6350 = _6342 ^ _6349;
  wire _6351 = r895 ^ r977;
  wire _6352 = r1057 ^ r1146;
  wire _6353 = _6351 ^ _6352;
  wire _6354 = r1193 ^ r1258;
  wire _6355 = r1348 ^ r1422;
  wire _6356 = _6354 ^ _6355;
  wire _6357 = _6353 ^ _6356;
  wire _6358 = r1440 ^ r1484;
  wire _6359 = r1487 ^ r1509;
  wire _6360 = _6358 ^ _6359;
  wire _6361 = r1527 ^ r1674;
  wire _6362 = r1689 ^ r1771;
  wire _6363 = _6361 ^ _6362;
  wire _6364 = _6360 ^ _6363;
  wire _6365 = _6357 ^ _6364;
  wire _6366 = _6350 ^ _6365;
  wire _6367 = r46 ^ r99;
  wire _6368 = r133 ^ r214;
  wire _6369 = _6367 ^ _6368;
  wire _6370 = r257 ^ r282;
  wire _6371 = r350 ^ r422;
  wire _6372 = _6370 ^ _6371;
  wire _6373 = _6369 ^ _6372;
  wire _6374 = r496 ^ r517;
  wire _6375 = r601 ^ r667;
  wire _6376 = _6374 ^ _6375;
  wire _6377 = r673 ^ r762;
  wire _6378 = r784 ^ r835;
  wire _6379 = _6377 ^ _6378;
  wire _6380 = _6376 ^ _6379;
  wire _6381 = _6373 ^ _6380;
  wire _6382 = r909 ^ r949;
  wire _6383 = r1049 ^ r1067;
  wire _6384 = _6382 ^ _6383;
  wire _6385 = r1150 ^ r1270;
  wire _6386 = r1280 ^ r1283;
  wire _6387 = _6385 ^ _6386;
  wire _6388 = _6384 ^ _6387;
  wire _6389 = r1363 ^ r1539;
  wire _6390 = r1562 ^ r1607;
  wire _6391 = _6389 ^ _6390;
  wire _6392 = r1627 ^ r1748;
  wire _6393 = r1765 ^ r1848;
  wire _6394 = _6392 ^ _6393;
  wire _6395 = _6391 ^ _6394;
  wire _6396 = _6388 ^ _6395;
  wire _6397 = _6381 ^ _6396;
  wire _6398 = _6366 | _6397;
  wire _6399 = _6335 | _6398;
  wire _6400 = _6272 | _6399;
  wire _6401 = r45 ^ r102;
  wire _6402 = r134 ^ r204;
  wire _6403 = _6401 ^ _6402;
  wire _6404 = r245 ^ r300;
  wire _6405 = r387 ^ r406;
  wire _6406 = _6404 ^ _6405;
  wire _6407 = _6403 ^ _6406;
  wire _6408 = r448 ^ r554;
  wire _6409 = r570 ^ r628;
  wire _6410 = _6408 ^ _6409;
  wire _6411 = r711 ^ r760;
  wire _6412 = r820 ^ r856;
  wire _6413 = _6411 ^ _6412;
  wire _6414 = _6410 ^ _6413;
  wire _6415 = _6407 ^ _6414;
  wire _6416 = r919 ^ r946;
  wire _6417 = r1024 ^ r1061;
  wire _6418 = _6416 ^ _6417;
  wire _6419 = r1139 ^ r1210;
  wire _6420 = r1241 ^ r1356;
  wire _6421 = _6419 ^ _6420;
  wire _6422 = _6418 ^ _6421;
  wire _6423 = r1386 ^ r1446;
  wire _6424 = r1532 ^ r1576;
  wire _6425 = _6423 ^ _6424;
  wire _6426 = r1613 ^ r1685;
  wire _6427 = r1707 ^ r1772;
  wire _6428 = _6426 ^ _6427;
  wire _6429 = _6425 ^ _6428;
  wire _6430 = _6422 ^ _6429;
  wire _6431 = _6415 ^ _6430;
  wire _6432 = r44 ^ r93;
  wire _6433 = r169 ^ r174;
  wire _6434 = _6432 ^ _6433;
  wire _6435 = r274 ^ r351;
  wire _6436 = r407 ^ r477;
  wire _6437 = _6435 ^ _6436;
  wire _6438 = _6434 ^ _6437;
  wire _6439 = r536 ^ r606;
  wire _6440 = r648 ^ r669;
  wire _6441 = _6439 ^ _6440;
  wire _6442 = r737 ^ r881;
  wire _6443 = r889 ^ r963;
  wire _6444 = _6442 ^ _6443;
  wire _6445 = _6441 ^ _6444;
  wire _6446 = _6438 ^ _6445;
  wire _6447 = r1033 ^ r1096;
  wire _6448 = r1119 ^ r1196;
  wire _6449 = _6447 ^ _6448;
  wire _6450 = r1231 ^ r1430;
  wire _6451 = r1450 ^ r1479;
  wire _6452 = _6450 ^ _6451;
  wire _6453 = _6449 ^ _6452;
  wire _6454 = r1531 ^ r1535;
  wire _6455 = r1747 ^ r1750;
  wire _6456 = _6454 ^ _6455;
  wire _6457 = r1758 ^ r1812;
  wire _6458 = r1835 ^ r1886;
  wire _6459 = _6457 ^ _6458;
  wire _6460 = _6456 ^ _6459;
  wire _6461 = _6453 ^ _6460;
  wire _6462 = _6446 ^ _6461;
  wire _6463 = _6431 | _6462;
  wire _6464 = r43 ^ r73;
  wire _6465 = r160 ^ r181;
  wire _6466 = _6464 ^ _6465;
  wire _6467 = r281 ^ r365;
  wire _6468 = r433 ^ r491;
  wire _6469 = _6467 ^ _6468;
  wire _6470 = _6466 ^ _6469;
  wire _6471 = r550 ^ r563;
  wire _6472 = r655 ^ r678;
  wire _6473 = _6471 ^ _6472;
  wire _6474 = r773 ^ r795;
  wire _6475 = r933 ^ r955;
  wire _6476 = _6474 ^ _6475;
  wire _6477 = _6473 ^ _6476;
  wire _6478 = _6470 ^ _6477;
  wire _6479 = r1027 ^ r1102;
  wire _6480 = r1159 ^ r1273;
  wire _6481 = _6479 ^ _6480;
  wire _6482 = r1328 ^ r1340;
  wire _6483 = r1426 ^ r1602;
  wire _6484 = _6482 ^ _6483;
  wire _6485 = _6481 ^ _6484;
  wire _6486 = r1724 ^ r1726;
  wire _6487 = r1761 ^ r1803;
  wire _6488 = _6486 ^ _6487;
  wire _6489 = r1839 ^ r1841;
  wire _6490 = r1868 ^ r1887;
  wire _6491 = _6489 ^ _6490;
  wire _6492 = _6488 ^ _6491;
  wire _6493 = _6485 ^ _6492;
  wire _6494 = _6478 ^ _6493;
  wire _6495 = r42 ^ r54;
  wire _6496 = r119 ^ r217;
  wire _6497 = _6495 ^ _6496;
  wire _6498 = r267 ^ r326;
  wire _6499 = r361 ^ r413;
  wire _6500 = _6498 ^ _6499;
  wire _6501 = _6497 ^ _6500;
  wire _6502 = r465 ^ r560;
  wire _6503 = r571 ^ r706;
  wire _6504 = _6502 ^ _6503;
  wire _6505 = r793 ^ r836;
  wire _6506 = r988 ^ r1030;
  wire _6507 = _6505 ^ _6506;
  wire _6508 = _6504 ^ _6507;
  wire _6509 = _6501 ^ _6508;
  wire _6510 = r1073 ^ r1234;
  wire _6511 = r1392 ^ r1460;
  wire _6512 = _6510 ^ _6511;
  wire _6513 = r1617 ^ r1679;
  wire _6514 = r1828 ^ r1871;
  wire _6515 = _6513 ^ _6514;
  wire _6516 = _6512 ^ _6515;
  wire _6517 = r1903 ^ r1912;
  wire _6518 = r1924 ^ r1953;
  wire _6519 = _6517 ^ _6518;
  wire _6520 = r1955 ^ r1956;
  wire _6521 = r2000 ^ r2006;
  wire _6522 = _6520 ^ _6521;
  wire _6523 = _6519 ^ _6522;
  wire _6524 = _6516 ^ _6523;
  wire _6525 = _6509 ^ _6524;
  wire _6526 = _6494 | _6525;
  wire _6527 = _6463 | _6526;
  wire _6528 = r41 ^ r68;
  wire _6529 = r123 ^ r219;
  wire _6530 = _6528 ^ _6529;
  wire _6531 = r251 ^ r288;
  wire _6532 = r382 ^ r425;
  wire _6533 = _6531 ^ _6532;
  wire _6534 = _6530 ^ _6533;
  wire _6535 = r499 ^ r530;
  wire _6536 = r600 ^ r656;
  wire _6537 = _6535 ^ _6536;
  wire _6538 = r694 ^ r763;
  wire _6539 = r826 ^ r883;
  wire _6540 = _6538 ^ _6539;
  wire _6541 = _6537 ^ _6540;
  wire _6542 = _6534 ^ _6541;
  wire _6543 = r936 ^ r998;
  wire _6544 = r1021 ^ r1071;
  wire _6545 = _6543 ^ _6544;
  wire _6546 = r1125 ^ r1252;
  wire _6547 = r1316 ^ r1385;
  wire _6548 = _6546 ^ _6547;
  wire _6549 = _6545 ^ _6548;
  wire _6550 = r1581 ^ r1632;
  wire _6551 = r1657 ^ r1745;
  wire _6552 = _6550 ^ _6551;
  wire _6553 = r1752 ^ r1763;
  wire _6554 = r1795 ^ r1849;
  wire _6555 = _6553 ^ _6554;
  wire _6556 = _6552 ^ _6555;
  wire _6557 = _6549 ^ _6556;
  wire _6558 = _6542 ^ _6557;
  wire _6559 = r170 ^ r276;
  wire _6560 = r345 ^ r434;
  wire _6561 = _6559 ^ _6560;
  wire _6562 = r613 ^ r647;
  wire _6563 = r738 ^ r870;
  wire _6564 = _6562 ^ _6563;
  wire _6565 = _6561 ^ _6564;
  wire _6566 = r901 ^ r1058;
  wire _6567 = r1181 ^ r1260;
  wire _6568 = _6566 ^ _6567;
  wire _6569 = r1286 ^ r1543;
  wire _6570 = r1553 ^ r1610;
  wire _6571 = _6569 ^ _6570;
  wire _6572 = _6568 ^ _6571;
  wire _6573 = _6565 ^ _6572;
  wire _6574 = r1684 ^ r1810;
  wire _6575 = r1914 ^ r1967;
  wire _6576 = _6574 ^ _6575;
  wire _6577 = r1977 ^ r1984;
  wire _6578 = r1989 ^ r1994;
  wire _6579 = _6577 ^ _6578;
  wire _6580 = _6576 ^ _6579;
  wire _6581 = r1997 ^ r2009;
  wire _6582 = r2015 ^ r2016;
  wire _6583 = _6581 ^ _6582;
  wire _6584 = r2025 ^ r2029;
  wire _6585 = r2036 ^ r2044;
  wire _6586 = _6584 ^ _6585;
  wire _6587 = _6583 ^ _6586;
  wire _6588 = _6580 ^ _6587;
  wire _6589 = _6573 ^ _6588;
  wire _6590 = _6558 | _6589;
  wire _6591 = r40 ^ r122;
  wire _6592 = r172 ^ r332;
  wire _6593 = _6591 ^ _6592;
  wire _6594 = r346 ^ r479;
  wire _6595 = r587 ^ r617;
  wire _6596 = _6594 ^ _6595;
  wire _6597 = _6593 ^ _6596;
  wire _6598 = r697 ^ r759;
  wire _6599 = r808 ^ r833;
  wire _6600 = _6598 ^ _6599;
  wire _6601 = r910 ^ r995;
  wire _6602 = r1039 ^ r1084;
  wire _6603 = _6601 ^ _6602;
  wire _6604 = _6600 ^ _6603;
  wire _6605 = _6597 ^ _6604;
  wire _6606 = r1141 ^ r1186;
  wire _6607 = r1256 ^ r1285;
  wire _6608 = _6606 ^ _6607;
  wire _6609 = r1331 ^ r1458;
  wire _6610 = r1473 ^ r1545;
  wire _6611 = _6609 ^ _6610;
  wire _6612 = _6608 ^ _6611;
  wire _6613 = r1652 ^ r1693;
  wire _6614 = r1824 ^ r1829;
  wire _6615 = _6613 ^ _6614;
  wire _6616 = r1869 ^ r1921;
  wire _6617 = r1930 ^ r1938;
  wire _6618 = _6616 ^ _6617;
  wire _6619 = _6615 ^ _6618;
  wire _6620 = _6612 ^ _6619;
  wire _6621 = _6605 ^ _6620;
  wire _6622 = r39 ^ r95;
  wire _6623 = r117 ^ r255;
  wire _6624 = _6622 ^ _6623;
  wire _6625 = r292 ^ r381;
  wire _6626 = r391 ^ r421;
  wire _6627 = _6625 ^ _6626;
  wire _6628 = _6624 ^ _6627;
  wire _6629 = r521 ^ r566;
  wire _6630 = r622 ^ r716;
  wire _6631 = _6629 ^ _6630;
  wire _6632 = r730 ^ r796;
  wire _6633 = r864 ^ r906;
  wire _6634 = _6632 ^ _6633;
  wire _6635 = _6631 ^ _6634;
  wire _6636 = _6628 ^ _6635;
  wire _6637 = r985 ^ r1053;
  wire _6638 = r1087 ^ r1128;
  wire _6639 = _6637 ^ _6638;
  wire _6640 = r1176 ^ r1261;
  wire _6641 = r1314 ^ r1347;
  wire _6642 = _6640 ^ _6641;
  wire _6643 = _6639 ^ _6642;
  wire _6644 = r1407 ^ r1434;
  wire _6645 = r1591 ^ r1622;
  wire _6646 = _6644 ^ _6645;
  wire _6647 = r1725 ^ r1881;
  wire _6648 = r1954 ^ r1963;
  wire _6649 = _6647 ^ _6648;
  wire _6650 = _6646 ^ _6649;
  wire _6651 = _6643 ^ _6650;
  wire _6652 = _6636 ^ _6651;
  wire _6653 = _6621 | _6652;
  wire _6654 = _6590 | _6653;
  wire _6655 = _6527 | _6654;
  wire _6656 = _6400 | _6655;
  wire _6657 = r38 ^ r82;
  wire _6658 = r157 ^ r191;
  wire _6659 = _6657 ^ _6658;
  wire _6660 = r286 ^ r372;
  wire _6661 = r393 ^ r494;
  wire _6662 = _6660 ^ _6661;
  wire _6663 = _6659 ^ _6662;
  wire _6664 = r542 ^ r588;
  wire _6665 = r660 ^ r770;
  wire _6666 = _6664 ^ _6665;
  wire _6667 = r861 ^ r911;
  wire _6668 = r1074 ^ r1144;
  wire _6669 = _6667 ^ _6668;
  wire _6670 = _6666 ^ _6669;
  wire _6671 = _6663 ^ _6670;
  wire _6672 = r1251 ^ r1298;
  wire _6673 = r1359 ^ r1435;
  wire _6674 = _6672 ^ _6673;
  wire _6675 = r1454 ^ r1551;
  wire _6676 = r1614 ^ r1678;
  wire _6677 = _6675 ^ _6676;
  wire _6678 = _6674 ^ _6677;
  wire _6679 = r1767 ^ r1813;
  wire _6680 = r1815 ^ r1862;
  wire _6681 = _6679 ^ _6680;
  wire _6682 = r1884 ^ r1894;
  wire _6683 = r1916 ^ r1919;
  wire _6684 = _6682 ^ _6683;
  wire _6685 = _6681 ^ _6684;
  wire _6686 = _6678 ^ _6685;
  wire _6687 = _6671 ^ _6686;
  wire _6688 = r37 ^ r97;
  wire _6689 = r165 ^ r218;
  wire _6690 = _6688 ^ _6689;
  wire _6691 = r323 ^ r428;
  wire _6692 = r461 ^ r552;
  wire _6693 = _6691 ^ _6692;
  wire _6694 = _6690 ^ _6693;
  wire _6695 = r662 ^ r719;
  wire _6696 = r740 ^ r792;
  wire _6697 = _6695 ^ _6696;
  wire _6698 = r875 ^ r900;
  wire _6699 = r945 ^ r1101;
  wire _6700 = _6698 ^ _6699;
  wire _6701 = _6697 ^ _6700;
  wire _6702 = _6694 ^ _6701;
  wire _6703 = r1205 ^ r1329;
  wire _6704 = r1399 ^ r1510;
  wire _6705 = _6703 ^ _6704;
  wire _6706 = r1565 ^ r1582;
  wire _6707 = r1642 ^ r1710;
  wire _6708 = _6706 ^ _6707;
  wire _6709 = _6705 ^ _6708;
  wire _6710 = r1844 ^ r1880;
  wire _6711 = r1907 ^ r1908;
  wire _6712 = _6710 ^ _6711;
  wire _6713 = r1917 ^ r1922;
  wire _6714 = r1931 ^ r1939;
  wire _6715 = _6713 ^ _6714;
  wire _6716 = _6712 ^ _6715;
  wire _6717 = _6709 ^ _6716;
  wire _6718 = _6702 ^ _6717;
  wire _6719 = _6687 | _6718;
  wire _6720 = r36 ^ r60;
  wire _6721 = r129 ^ r180;
  wire _6722 = _6720 ^ _6721;
  wire _6723 = r246 ^ r330;
  wire _6724 = r335 ^ r395;
  wire _6725 = _6723 ^ _6724;
  wire _6726 = _6722 ^ _6725;
  wire _6727 = r462 ^ r547;
  wire _6728 = r598 ^ r630;
  wire _6729 = _6727 ^ _6728;
  wire _6730 = r671 ^ r731;
  wire _6731 = r818 ^ r867;
  wire _6732 = _6730 ^ _6731;
  wire _6733 = _6729 ^ _6732;
  wire _6734 = _6726 ^ _6733;
  wire _6735 = r924 ^ r959;
  wire _6736 = r1023 ^ r1070;
  wire _6737 = _6735 ^ _6736;
  wire _6738 = r1116 ^ r1164;
  wire _6739 = r1190 ^ r1226;
  wire _6740 = _6738 ^ _6739;
  wire _6741 = _6737 ^ _6740;
  wire _6742 = r1287 ^ r1341;
  wire _6743 = r1408 ^ r1441;
  wire _6744 = _6742 ^ _6743;
  wire _6745 = r1459 ^ r1491;
  wire _6746 = r1694 ^ r1773;
  wire _6747 = _6745 ^ _6746;
  wire _6748 = _6744 ^ _6747;
  wire _6749 = _6741 ^ _6748;
  wire _6750 = _6734 ^ _6749;
  wire _6751 = r35 ^ r70;
  wire _6752 = r127 ^ r206;
  wire _6753 = _6751 ^ _6752;
  wire _6754 = r260 ^ r298;
  wire _6755 = r408 ^ r493;
  wire _6756 = _6754 ^ _6755;
  wire _6757 = _6753 ^ _6756;
  wire _6758 = r553 ^ r561;
  wire _6759 = r715 ^ r774;
  wire _6760 = _6758 ^ _6759;
  wire _6761 = r802 ^ r844;
  wire _6762 = r930 ^ r970;
  wire _6763 = _6761 ^ _6762;
  wire _6764 = _6760 ^ _6763;
  wire _6765 = _6757 ^ _6764;
  wire _6766 = r1010 ^ r1094;
  wire _6767 = r1167 ^ r1192;
  wire _6768 = _6766 ^ _6767;
  wire _6769 = r1265 ^ r1315;
  wire _6770 = r1496 ^ r1513;
  wire _6771 = _6769 ^ _6770;
  wire _6772 = _6768 ^ _6771;
  wire _6773 = r1534 ^ r1544;
  wire _6774 = r1559 ^ r1579;
  wire _6775 = _6773 ^ _6774;
  wire _6776 = r1645 ^ r1738;
  wire _6777 = r1743 ^ r1850;
  wire _6778 = _6776 ^ _6777;
  wire _6779 = _6775 ^ _6778;
  wire _6780 = _6772 ^ _6779;
  wire _6781 = _6765 ^ _6780;
  wire _6782 = _6750 | _6781;
  wire _6783 = _6719 | _6782;
  wire _6784 = r34 ^ r65;
  wire _6785 = r163 ^ r186;
  wire _6786 = _6784 ^ _6785;
  wire _6787 = r296 ^ r405;
  wire _6788 = r541 ^ r683;
  wire _6789 = _6787 ^ _6788;
  wire _6790 = _6786 ^ _6789;
  wire _6791 = r827 ^ r999;
  wire _6792 = r1025 ^ r1080;
  wire _6793 = _6791 ^ _6792;
  wire _6794 = r1117 ^ r1267;
  wire _6795 = r1372 ^ r1395;
  wire _6796 = _6794 ^ _6795;
  wire _6797 = _6793 ^ _6796;
  wire _6798 = _6790 ^ _6797;
  wire _6799 = r1488 ^ r1566;
  wire _6800 = r1712 ^ r1730;
  wire _6801 = _6799 ^ _6800;
  wire _6802 = r1737 ^ r1796;
  wire _6803 = r1865 ^ r1875;
  wire _6804 = _6802 ^ _6803;
  wire _6805 = _6801 ^ _6804;
  wire _6806 = r1895 ^ r1896;
  wire _6807 = r1898 ^ r1900;
  wire _6808 = _6806 ^ _6807;
  wire _6809 = r1902 ^ r1905;
  wire _6810 = r1934 ^ r1945;
  wire _6811 = _6809 ^ _6810;
  wire _6812 = _6808 ^ _6811;
  wire _6813 = _6805 ^ _6812;
  wire _6814 = _6798 ^ _6813;
  wire _6815 = r33 ^ r71;
  wire _6816 = r142 ^ r230;
  wire _6817 = _6815 ^ _6816;
  wire _6818 = r389 ^ r503;
  wire _6819 = r583 ^ r631;
  wire _6820 = _6818 ^ _6819;
  wire _6821 = _6817 ^ _6820;
  wire _6822 = r767 ^ r848;
  wire _6823 = r916 ^ r987;
  wire _6824 = _6822 ^ _6823;
  wire _6825 = r1045 ^ r1103;
  wire _6826 = r1197 ^ r1237;
  wire _6827 = _6825 ^ _6826;
  wire _6828 = _6824 ^ _6827;
  wire _6829 = _6821 ^ _6828;
  wire _6830 = r1307 ^ r1330;
  wire _6831 = r1423 ^ r1639;
  wire _6832 = _6830 ^ _6831;
  wire _6833 = r1680 ^ r1692;
  wire _6834 = r1915 ^ r1918;
  wire _6835 = _6833 ^ _6834;
  wire _6836 = _6832 ^ _6835;
  wire _6837 = r1957 ^ r1974;
  wire _6838 = r1975 ^ r2002;
  wire _6839 = _6837 ^ _6838;
  wire _6840 = r2012 ^ r2018;
  wire _6841 = r2021 ^ r2037;
  wire _6842 = _6840 ^ _6841;
  wire _6843 = _6839 ^ _6842;
  wire _6844 = _6836 ^ _6843;
  wire _6845 = _6829 ^ _6844;
  wire _6846 = _6814 | _6845;
  wire _6847 = r32 ^ r59;
  wire _6848 = r145 ^ r220;
  wire _6849 = _6847 ^ _6848;
  wire _6850 = r240 ^ r308;
  wire _6851 = r369 ^ r445;
  wire _6852 = _6850 ^ _6851;
  wire _6853 = _6849 ^ _6852;
  wire _6854 = r451 ^ r515;
  wire _6855 = r615 ^ r661;
  wire _6856 = _6854 ^ _6855;
  wire _6857 = r674 ^ r764;
  wire _6858 = r806 ^ r852;
  wire _6859 = _6857 ^ _6858;
  wire _6860 = _6856 ^ _6859;
  wire _6861 = _6853 ^ _6860;
  wire _6862 = r940 ^ r973;
  wire _6863 = r1055 ^ r1095;
  wire _6864 = _6862 ^ _6863;
  wire _6865 = r1130 ^ r1209;
  wire _6866 = r1274 ^ r1295;
  wire _6867 = _6865 ^ _6866;
  wire _6868 = _6864 ^ _6867;
  wire _6869 = r1353 ^ r1402;
  wire _6870 = r1453 ^ r1461;
  wire _6871 = _6869 ^ _6870;
  wire _6872 = r1472 ^ r1623;
  wire _6873 = r1677 ^ r1774;
  wire _6874 = _6872 ^ _6873;
  wire _6875 = _6871 ^ _6874;
  wire _6876 = _6868 ^ _6875;
  wire _6877 = _6861 ^ _6876;
  wire _6878 = r31 ^ r85;
  wire _6879 = r130 ^ r216;
  wire _6880 = _6878 ^ _6879;
  wire _6881 = r234 ^ r311;
  wire _6882 = r377 ^ r446;
  wire _6883 = _6881 ^ _6882;
  wire _6884 = _6880 ^ _6883;
  wire _6885 = r505 ^ r556;
  wire _6886 = r607 ^ r621;
  wire _6887 = _6885 ^ _6886;
  wire _6888 = r676 ^ r724;
  wire _6889 = r825 ^ r841;
  wire _6890 = _6888 ^ _6889;
  wire _6891 = _6887 ^ _6890;
  wire _6892 = _6884 ^ _6891;
  wire _6893 = r922 ^ r990;
  wire _6894 = r1050 ^ r1085;
  wire _6895 = _6893 ^ _6894;
  wire _6896 = r1137 ^ r1215;
  wire _6897 = r1224 ^ r1230;
  wire _6898 = _6896 ^ _6897;
  wire _6899 = _6895 ^ _6898;
  wire _6900 = r1317 ^ r1361;
  wire _6901 = r1387 ^ r1425;
  wire _6902 = _6900 ^ _6901;
  wire _6903 = r1601 ^ r1608;
  wire _6904 = r1651 ^ r1775;
  wire _6905 = _6903 ^ _6904;
  wire _6906 = _6902 ^ _6905;
  wire _6907 = _6899 ^ _6906;
  wire _6908 = _6892 ^ _6907;
  wire _6909 = _6877 | _6908;
  wire _6910 = _6846 | _6909;
  wire _6911 = _6783 | _6910;
  wire _6912 = r30 ^ r91;
  wire _6913 = r164 ^ r183;
  wire _6914 = _6912 ^ _6913;
  wire _6915 = r237 ^ r299;
  wire _6916 = r341 ^ r423;
  wire _6917 = _6915 ^ _6916;
  wire _6918 = _6914 ^ _6917;
  wire _6919 = r450 ^ r558;
  wire _6920 = r649 ^ r701;
  wire _6921 = _6919 ^ _6920;
  wire _6922 = r772 ^ r876;
  wire _6923 = r932 ^ r951;
  wire _6924 = _6922 ^ _6923;
  wire _6925 = _6921 ^ _6924;
  wire _6926 = _6918 ^ _6925;
  wire _6927 = r1056 ^ r1100;
  wire _6928 = r1108 ^ r1121;
  wire _6929 = _6927 ^ _6928;
  wire _6930 = r1191 ^ r1238;
  wire _6931 = r1309 ^ r1357;
  wire _6932 = _6930 ^ _6931;
  wire _6933 = _6929 ^ _6932;
  wire _6934 = r1546 ^ r1561;
  wire _6935 = r1618 ^ r1713;
  wire _6936 = _6934 ^ _6935;
  wire _6937 = r1766 ^ r1797;
  wire _6938 = r1821 ^ r1888;
  wire _6939 = _6937 ^ _6938;
  wire _6940 = _6936 ^ _6939;
  wire _6941 = _6933 ^ _6940;
  wire _6942 = _6926 ^ _6941;
  wire _6943 = r29 ^ r75;
  wire _6944 = r126 ^ r201;
  wire _6945 = _6943 ^ _6944;
  wire _6946 = r227 ^ r329;
  wire _6947 = r339 ^ r414;
  wire _6948 = _6946 ^ _6947;
  wire _6949 = _6945 ^ _6948;
  wire _6950 = r501 ^ r524;
  wire _6951 = r574 ^ r627;
  wire _6952 = _6950 ^ _6951;
  wire _6953 = r681 ^ r747;
  wire _6954 = r797 ^ r860;
  wire _6955 = _6953 ^ _6954;
  wire _6956 = _6952 ^ _6955;
  wire _6957 = _6949 ^ _6956;
  wire _6958 = r941 ^ r961;
  wire _6959 = r1044 ^ r1078;
  wire _6960 = _6958 ^ _6959;
  wire _6961 = r1122 ^ r1204;
  wire _6962 = r1266 ^ r1299;
  wire _6963 = _6961 ^ _6962;
  wire _6964 = _6960 ^ _6963;
  wire _6965 = r1332 ^ r1362;
  wire _6966 = r1389 ^ r1542;
  wire _6967 = _6965 ^ _6966;
  wire _6968 = r1606 ^ r1628;
  wire _6969 = r1667 ^ r1776;
  wire _6970 = _6968 ^ _6969;
  wire _6971 = _6967 ^ _6970;
  wire _6972 = _6964 ^ _6971;
  wire _6973 = _6957 ^ _6972;
  wire _6974 = _6942 | _6973;
  wire _6975 = r28 ^ r77;
  wire _6976 = r154 ^ r202;
  wire _6977 = _6975 ^ _6976;
  wire _6978 = r261 ^ r295;
  wire _6979 = r375 ^ r432;
  wire _6980 = _6978 ^ _6979;
  wire _6981 = _6977 ^ _6980;
  wire _6982 = r483 ^ r508;
  wire _6983 = r616 ^ r651;
  wire _6984 = _6982 ^ _6983;
  wire _6985 = r693 ^ r757;
  wire _6986 = r811 ^ r871;
  wire _6987 = _6985 ^ _6986;
  wire _6988 = _6984 ^ _6987;
  wire _6989 = _6981 ^ _6988;
  wire _6990 = r915 ^ r956;
  wire _6991 = r1013 ^ r1076;
  wire _6992 = _6990 ^ _6991;
  wire _6993 = r1148 ^ r1177;
  wire _6994 = r1225 ^ r1277;
  wire _6995 = _6993 ^ _6994;
  wire _6996 = _6992 ^ _6995;
  wire _6997 = r1313 ^ r1352;
  wire _6998 = r1397 ^ r1436;
  wire _6999 = _6997 ^ _6998;
  wire _7000 = r1492 ^ r1586;
  wire _7001 = r1698 ^ r1777;
  wire _7002 = _7000 ^ _7001;
  wire _7003 = _6999 ^ _7002;
  wire _7004 = _6996 ^ _7003;
  wire _7005 = _6989 ^ _7004;
  wire _7006 = r27 ^ r101;
  wire _7007 = r138 ^ r182;
  wire _7008 = _7006 ^ _7007;
  wire _7009 = r321 ^ r354;
  wire _7010 = r437 ^ r489;
  wire _7011 = _7009 ^ _7010;
  wire _7012 = _7008 ^ _7011;
  wire _7013 = r518 ^ r573;
  wire _7014 = r663 ^ r702;
  wire _7015 = _7013 ^ _7014;
  wire _7016 = r750 ^ r804;
  wire _7017 = r882 ^ r929;
  wire _7018 = _7016 ^ _7017;
  wire _7019 = _7015 ^ _7018;
  wire _7020 = _7012 ^ _7019;
  wire _7021 = r962 ^ r1019;
  wire _7022 = r1089 ^ r1129;
  wire _7023 = _7021 ^ _7022;
  wire _7024 = r1165 ^ r1212;
  wire _7025 = r1253 ^ r1292;
  wire _7026 = _7024 ^ _7025;
  wire _7027 = _7023 ^ _7026;
  wire _7028 = r1375 ^ r1419;
  wire _7029 = r1433 ^ r1641;
  wire _7030 = _7028 ^ _7029;
  wire _7031 = r1705 ^ r1757;
  wire _7032 = r1801 ^ r1851;
  wire _7033 = _7031 ^ _7032;
  wire _7034 = _7030 ^ _7033;
  wire _7035 = _7027 ^ _7034;
  wire _7036 = _7020 ^ _7035;
  wire _7037 = _7005 | _7036;
  wire _7038 = _6974 | _7037;
  wire _7039 = r26 ^ r83;
  wire _7040 = r166 ^ r173;
  wire _7041 = _7039 ^ _7040;
  wire _7042 = r256 ^ r305;
  wire _7043 = r356 ^ r447;
  wire _7044 = _7042 ^ _7043;
  wire _7045 = _7041 ^ _7044;
  wire _7046 = r457 ^ r525;
  wire _7047 = r568 ^ r659;
  wire _7048 = _7046 ^ _7047;
  wire _7049 = r675 ^ r754;
  wire _7050 = r781 ^ r855;
  wire _7051 = _7049 ^ _7050;
  wire _7052 = _7048 ^ _7051;
  wire _7053 = _7045 ^ _7052;
  wire _7054 = r902 ^ r950;
  wire _7055 = r1004 ^ r1082;
  wire _7056 = _7054 ^ _7055;
  wire _7057 = r1140 ^ r1179;
  wire _7058 = r1233 ^ r1282;
  wire _7059 = _7057 ^ _7058;
  wire _7060 = _7056 ^ _7059;
  wire _7061 = r1289 ^ r1381;
  wire _7062 = r1420 ^ r1475;
  wire _7063 = _7061 ^ _7062;
  wire _7064 = r1594 ^ r1629;
  wire _7065 = r1656 ^ r1778;
  wire _7066 = _7064 ^ _7065;
  wire _7067 = _7063 ^ _7066;
  wire _7068 = _7060 ^ _7067;
  wire _7069 = _7053 ^ _7068;
  wire _7070 = r25 ^ r94;
  wire _7071 = r156 ^ r190;
  wire _7072 = _7070 ^ _7071;
  wire _7073 = r268 ^ r331;
  wire _7074 = r342 ^ r436;
  wire _7075 = _7073 ^ _7074;
  wire _7076 = _7072 ^ _7075;
  wire _7077 = r455 ^ r557;
  wire _7078 = r604 ^ r624;
  wire _7079 = _7077 ^ _7078;
  wire _7080 = r689 ^ r791;
  wire _7081 = r843 ^ r935;
  wire _7082 = _7080 ^ _7081;
  wire _7083 = _7079 ^ _7082;
  wire _7084 = _7076 ^ _7083;
  wire _7085 = r976 ^ r1111;
  wire _7086 = r1149 ^ r1302;
  wire _7087 = _7085 ^ _7086;
  wire _7088 = r1334 ^ r1365;
  wire _7089 = r1396 ^ r1590;
  wire _7090 = _7088 ^ _7089;
  wire _7091 = _7087 ^ _7090;
  wire _7092 = r1660 ^ r1704;
  wire _7093 = r1727 ^ r1876;
  wire _7094 = _7092 ^ _7093;
  wire _7095 = r1882 ^ r1935;
  wire _7096 = r1940 ^ r1946;
  wire _7097 = _7095 ^ _7096;
  wire _7098 = _7094 ^ _7097;
  wire _7099 = _7091 ^ _7098;
  wire _7100 = _7084 ^ _7099;
  wire _7101 = _7069 | _7100;
  wire _7102 = r24 ^ r143;
  wire _7103 = r241 ^ r376;
  wire _7104 = _7102 ^ _7103;
  wire _7105 = r430 ^ r487;
  wire _7106 = r611 ^ r644;
  wire _7107 = _7105 ^ _7106;
  wire _7108 = _7104 ^ _7107;
  wire _7109 = r777 ^ r885;
  wire _7110 = r904 ^ r982;
  wire _7111 = _7109 ^ _7110;
  wire _7112 = r1189 ^ r1268;
  wire _7113 = r1367 ^ r1391;
  wire _7114 = _7112 ^ _7113;
  wire _7115 = _7111 ^ _7114;
  wire _7116 = _7108 ^ _7115;
  wire _7117 = r1687 ^ r1749;
  wire _7118 = r1820 ^ r1823;
  wire _7119 = _7117 ^ _7118;
  wire _7120 = r1870 ^ r1913;
  wire _7121 = r1932 ^ r1969;
  wire _7122 = _7120 ^ _7121;
  wire _7123 = _7119 ^ _7122;
  wire _7124 = r1973 ^ r1982;
  wire _7125 = r2007 ^ r2023;
  wire _7126 = _7124 ^ _7125;
  wire _7127 = r2033 ^ r2035;
  wire _7128 = r2041 ^ r2046;
  wire _7129 = _7127 ^ _7128;
  wire _7130 = _7126 ^ _7129;
  wire _7131 = _7123 ^ _7130;
  wire _7132 = _7116 ^ _7131;
  wire _7133 = r23 ^ r76;
  wire _7134 = r162 ^ r224;
  wire _7135 = _7133 ^ _7134;
  wire _7136 = r229 ^ r309;
  wire _7137 = r338 ^ r411;
  wire _7138 = _7136 ^ _7137;
  wire _7139 = _7135 ^ _7138;
  wire _7140 = r469 ^ r543;
  wire _7141 = r579 ^ r645;
  wire _7142 = _7140 ^ _7141;
  wire _7143 = r696 ^ r788;
  wire _7144 = r846 ^ r917;
  wire _7145 = _7143 ^ _7144;
  wire _7146 = _7142 ^ _7145;
  wire _7147 = _7139 ^ _7146;
  wire _7148 = r965 ^ r1011;
  wire _7149 = r1062 ^ r1136;
  wire _7150 = _7148 ^ _7149;
  wire _7151 = r1169 ^ r1207;
  wire _7152 = r1264 ^ r1325;
  wire _7153 = _7151 ^ _7152;
  wire _7154 = _7150 ^ _7153;
  wire _7155 = r1336 ^ r1406;
  wire _7156 = r1474 ^ r1577;
  wire _7157 = _7155 ^ _7156;
  wire _7158 = r1620 ^ r1659;
  wire _7159 = r1714 ^ r1779;
  wire _7160 = _7158 ^ _7159;
  wire _7161 = _7157 ^ _7160;
  wire _7162 = _7154 ^ _7161;
  wire _7163 = _7147 ^ _7162;
  wire _7164 = _7132 | _7163;
  wire _7165 = _7101 | _7164;
  wire _7166 = _7038 | _7165;
  wire _7167 = _6911 | _7166;
  wire _7168 = _6656 | _7167;
  wire _7169 = r22 ^ r90;
  wire _7170 = r135 ^ r193;
  wire _7171 = _7169 ^ _7170;
  wire _7172 = r270 ^ r328;
  wire _7173 = r366 ^ r419;
  wire _7174 = _7172 ^ _7173;
  wire _7175 = _7171 ^ _7174;
  wire _7176 = r472 ^ r520;
  wire _7177 = r623 ^ r718;
  wire _7178 = _7176 ^ _7177;
  wire _7179 = r775 ^ r779;
  wire _7180 = r865 ^ r914;
  wire _7181 = _7179 ^ _7180;
  wire _7182 = _7178 ^ _7181;
  wire _7183 = _7175 ^ _7182;
  wire _7184 = r967 ^ r1022;
  wire _7185 = r1066 ^ r1112;
  wire _7186 = _7184 ^ _7185;
  wire _7187 = r1174 ^ r1228;
  wire _7188 = r1284 ^ r1373;
  wire _7189 = _7187 ^ _7188;
  wire _7190 = _7186 ^ _7189;
  wire _7191 = r1411 ^ r1442;
  wire _7192 = r1480 ^ r1511;
  wire _7193 = _7191 ^ _7192;
  wire _7194 = r1615 ^ r1655;
  wire _7195 = r1708 ^ r1780;
  wire _7196 = _7194 ^ _7195;
  wire _7197 = _7193 ^ _7196;
  wire _7198 = _7190 ^ _7197;
  wire _7199 = _7183 ^ _7198;
  wire _7200 = r21 ^ r61;
  wire _7201 = r132 ^ r188;
  wire _7202 = _7200 ^ _7201;
  wire _7203 = r232 ^ r301;
  wire _7204 = r441 ^ r458;
  wire _7205 = _7203 ^ _7204;
  wire _7206 = _7202 ^ _7205;
  wire _7207 = r545 ^ r609;
  wire _7208 = r812 ^ r873;
  wire _7209 = _7207 ^ _7208;
  wire _7210 = r993 ^ r1029;
  wire _7211 = r1143 ^ r1248;
  wire _7212 = _7210 ^ _7211;
  wire _7213 = _7209 ^ _7212;
  wire _7214 = _7206 ^ _7213;
  wire _7215 = r1486 ^ r1506;
  wire _7216 = r1526 ^ r1533;
  wire _7217 = _7215 ^ _7216;
  wire _7218 = r1552 ^ r1564;
  wire _7219 = r1621 ^ r1682;
  wire _7220 = _7218 ^ _7219;
  wire _7221 = _7217 ^ _7220;
  wire _7222 = r1739 ^ r1800;
  wire _7223 = r1873 ^ r1874;
  wire _7224 = _7222 ^ _7223;
  wire _7225 = r1925 ^ r1948;
  wire _7226 = r1958 ^ r1965;
  wire _7227 = _7225 ^ _7226;
  wire _7228 = _7224 ^ _7227;
  wire _7229 = _7221 ^ _7228;
  wire _7230 = _7214 ^ _7229;
  wire _7231 = _7199 | _7230;
  wire _7232 = r20 ^ r148;
  wire _7233 = r378 ^ r488;
  wire _7234 = _7232 ^ _7233;
  wire _7235 = r591 ^ r758;
  wire _7236 = r868 ^ r897;
  wire _7237 = _7235 ^ _7236;
  wire _7238 = _7234 ^ _7237;
  wire _7239 = r974 ^ r1005;
  wire _7240 = r1206 ^ r1249;
  wire _7241 = _7239 ^ _7240;
  wire _7242 = r1337 ^ r1410;
  wire _7243 = r1451 ^ r1466;
  wire _7244 = _7242 ^ _7243;
  wire _7245 = _7241 ^ _7244;
  wire _7246 = _7238 ^ _7245;
  wire _7247 = r1530 ^ r1569;
  wire _7248 = r1611 ^ r1649;
  wire _7249 = _7247 ^ _7248;
  wire _7250 = r1688 ^ r1825;
  wire _7251 = r1943 ^ r1964;
  wire _7252 = _7250 ^ _7251;
  wire _7253 = _7249 ^ _7252;
  wire _7254 = r1970 ^ r1990;
  wire _7255 = r1993 ^ r2003;
  wire _7256 = _7254 ^ _7255;
  wire _7257 = r2017 ^ r2026;
  wire _7258 = r2034 ^ r2045;
  wire _7259 = _7257 ^ _7258;
  wire _7260 = _7256 ^ _7259;
  wire _7261 = _7253 ^ _7260;
  wire _7262 = _7246 ^ _7261;
  wire _7263 = r19 ^ r63;
  wire _7264 = r140 ^ r178;
  wire _7265 = _7263 ^ _7264;
  wire _7266 = r258 ^ r314;
  wire _7267 = r368 ^ r417;
  wire _7268 = _7266 ^ _7267;
  wire _7269 = _7265 ^ _7268;
  wire _7270 = r454 ^ r555;
  wire _7271 = r593 ^ r634;
  wire _7272 = _7270 ^ _7271;
  wire _7273 = r691 ^ r746;
  wire _7274 = r807 ^ r874;
  wire _7275 = _7273 ^ _7274;
  wire _7276 = _7272 ^ _7275;
  wire _7277 = _7269 ^ _7276;
  wire _7278 = r898 ^ r986;
  wire _7279 = r1018 ^ r1075;
  wire _7280 = _7278 ^ _7279;
  wire _7281 = r1123 ^ r1198;
  wire _7282 = r1227 ^ r1322;
  wire _7283 = _7281 ^ _7282;
  wire _7284 = _7280 ^ _7283;
  wire _7285 = r1366 ^ r1404;
  wire _7286 = r1445 ^ r1575;
  wire _7287 = _7285 ^ _7286;
  wire _7288 = r1595 ^ r1631;
  wire _7289 = r1706 ^ r1781;
  wire _7290 = _7288 ^ _7289;
  wire _7291 = _7287 ^ _7290;
  wire _7292 = _7284 ^ _7291;
  wire _7293 = _7277 ^ _7292;
  wire _7294 = _7262 | _7293;
  wire _7295 = _7231 | _7294;
  wire _7296 = r18 ^ r78;
  wire _7297 = r114 ^ r198;
  wire _7298 = _7296 ^ _7297;
  wire _7299 = r253 ^ r307;
  wire _7300 = r398 ^ r480;
  wire _7301 = _7299 ^ _7300;
  wire _7302 = _7298 ^ _7301;
  wire _7303 = r580 ^ r668;
  wire _7304 = r713 ^ r733;
  wire _7305 = _7303 ^ _7304;
  wire _7306 = r819 ^ r994;
  wire _7307 = r1046 ^ r1086;
  wire _7308 = _7306 ^ _7307;
  wire _7309 = _7305 ^ _7308;
  wire _7310 = _7302 ^ _7309;
  wire _7311 = r1120 ^ r1275;
  wire _7312 = r1303 ^ r1380;
  wire _7313 = _7311 ^ _7312;
  wire _7314 = r1449 ^ r1549;
  wire _7315 = r1568 ^ r1583;
  wire _7316 = _7314 ^ _7315;
  wire _7317 = _7313 ^ _7316;
  wire _7318 = r1697 ^ r1863;
  wire _7319 = r1937 ^ r1942;
  wire _7320 = _7318 ^ _7319;
  wire _7321 = r1962 ^ r1972;
  wire _7322 = r1998 ^ r2004;
  wire _7323 = _7321 ^ _7322;
  wire _7324 = _7320 ^ _7323;
  wire _7325 = _7317 ^ _7324;
  wire _7326 = _7310 ^ _7325;
  wire _7327 = r17 ^ r74;
  wire _7328 = r124 ^ r259;
  wire _7329 = _7327 ^ _7328;
  wire _7330 = r374 ^ r466;
  wire _7331 = r538 ^ r610;
  wire _7332 = _7330 ^ _7331;
  wire _7333 = _7329 ^ _7332;
  wire _7334 = r633 ^ r832;
  wire _7335 = r923 ^ r966;
  wire _7336 = _7334 ^ _7335;
  wire _7337 = r1236 ^ r1288;
  wire _7338 = r1354 ^ r1495;
  wire _7339 = _7337 ^ _7338;
  wire _7340 = _7336 ^ _7339;
  wire _7341 = _7333 ^ _7340;
  wire _7342 = r1515 ^ r1556;
  wire _7343 = r1625 ^ r1798;
  wire _7344 = _7342 ^ _7343;
  wire _7345 = r1842 ^ r1878;
  wire _7346 = r1959 ^ r1976;
  wire _7347 = _7345 ^ _7346;
  wire _7348 = _7344 ^ _7347;
  wire _7349 = r1981 ^ r1988;
  wire _7350 = r1991 ^ r2001;
  wire _7351 = _7349 ^ _7350;
  wire _7352 = r2010 ^ r2019;
  wire _7353 = r2031 ^ r2043;
  wire _7354 = _7352 ^ _7353;
  wire _7355 = _7351 ^ _7354;
  wire _7356 = _7348 ^ _7355;
  wire _7357 = _7341 ^ _7356;
  wire _7358 = _7326 | _7357;
  wire _7359 = r16 ^ r118;
  wire _7360 = r176 ^ r249;
  wire _7361 = _7359 ^ _7360;
  wire _7362 = r293 ^ r347;
  wire _7363 = r442 ^ r490;
  wire _7364 = _7362 ^ _7363;
  wire _7365 = _7361 ^ _7364;
  wire _7366 = r539 ^ r577;
  wire _7367 = r690 ^ r780;
  wire _7368 = _7366 ^ _7367;
  wire _7369 = r838 ^ r939;
  wire _7370 = r981 ^ r1048;
  wire _7371 = _7369 ^ _7370;
  wire _7372 = _7368 ^ _7371;
  wire _7373 = _7365 ^ _7372;
  wire _7374 = r1069 ^ r1161;
  wire _7375 = r1218 ^ r1240;
  wire _7376 = _7374 ^ _7375;
  wire _7377 = r1300 ^ r1519;
  wire _7378 = r1600 ^ r1626;
  wire _7379 = _7377 ^ _7378;
  wire _7380 = _7376 ^ _7379;
  wire _7381 = r1700 ^ r1809;
  wire _7382 = r1819 ^ r1831;
  wire _7383 = _7381 ^ _7382;
  wire _7384 = r1949 ^ r1978;
  wire _7385 = r1996 ^ r2005;
  wire _7386 = _7384 ^ _7385;
  wire _7387 = _7383 ^ _7386;
  wire _7388 = _7380 ^ _7387;
  wire _7389 = _7373 ^ _7388;
  wire _7390 = r15 ^ r56;
  wire _7391 = r209 ^ r272;
  wire _7392 = _7390 ^ _7391;
  wire _7393 = r287 ^ r344;
  wire _7394 = r418 ^ r482;
  wire _7395 = _7393 ^ _7394;
  wire _7396 = _7392 ^ _7395;
  wire _7397 = r516 ^ r602;
  wire _7398 = r666 ^ r682;
  wire _7399 = _7397 ^ _7398;
  wire _7400 = r722 ^ r776;
  wire _7401 = r821 ^ r877;
  wire _7402 = _7400 ^ _7401;
  wire _7403 = _7399 ^ _7402;
  wire _7404 = _7396 ^ _7403;
  wire _7405 = r943 ^ r952;
  wire _7406 = r1006 ^ r1162;
  wire _7407 = _7405 ^ _7406;
  wire _7408 = r1217 ^ r1308;
  wire _7409 = r1355 ^ r1414;
  wire _7410 = _7408 ^ _7409;
  wire _7411 = _7407 ^ _7410;
  wire _7412 = r1470 ^ r1507;
  wire _7413 = r1525 ^ r1578;
  wire _7414 = _7412 ^ _7413;
  wire _7415 = r1647 ^ r1672;
  wire _7416 = r1804 ^ r1852;
  wire _7417 = _7415 ^ _7416;
  wire _7418 = _7414 ^ _7417;
  wire _7419 = _7411 ^ _7418;
  wire _7420 = _7404 ^ _7419;
  wire _7421 = _7389 | _7420;
  wire _7422 = _7358 | _7421;
  wire _7423 = _7295 | _7422;
  wire _7424 = r14 ^ r57;
  wire _7425 = r212 ^ r278;
  wire _7426 = _7424 ^ _7425;
  wire _7427 = r291 ^ r359;
  wire _7428 = r439 ^ r470;
  wire _7429 = _7427 ^ _7428;
  wire _7430 = _7426 ^ _7429;
  wire _7431 = r509 ^ r700;
  wire _7432 = r783 ^ r879;
  wire _7433 = _7431 ^ _7432;
  wire _7434 = r989 ^ r1097;
  wire _7435 = r1138 ^ r1166;
  wire _7436 = _7434 ^ _7435;
  wire _7437 = _7433 ^ _7436;
  wire _7438 = _7430 ^ _7437;
  wire _7439 = r1213 ^ r1368;
  wire _7440 = r1476 ^ r1502;
  wire _7441 = _7439 ^ _7440;
  wire _7442 = r1504 ^ r1573;
  wire _7443 = r1664 ^ r1746;
  wire _7444 = _7442 ^ _7443;
  wire _7445 = _7441 ^ _7444;
  wire _7446 = r1756 ^ r1760;
  wire _7447 = r1864 ^ r1910;
  wire _7448 = _7446 ^ _7447;
  wire _7449 = r1920 ^ r1951;
  wire _7450 = r1952 ^ r1966;
  wire _7451 = _7449 ^ _7450;
  wire _7452 = _7448 ^ _7451;
  wire _7453 = _7445 ^ _7452;
  wire _7454 = _7438 ^ _7453;
  wire _7455 = r13 ^ r92;
  wire _7456 = r149 ^ r263;
  wire _7457 = _7455 ^ _7456;
  wire _7458 = r352 ^ r486;
  wire _7459 = r612 ^ r640;
  wire _7460 = _7458 ^ _7459;
  wire _7461 = _7457 ^ _7460;
  wire _7462 = r723 ^ r850;
  wire _7463 = r954 ^ r1195;
  wire _7464 = _7462 ^ _7463;
  wire _7465 = r1276 ^ r1324;
  wire _7466 = r1364 ^ r1494;
  wire _7467 = _7465 ^ _7466;
  wire _7468 = _7464 ^ _7467;
  wire _7469 = _7461 ^ _7468;
  wire _7470 = r1537 ^ r1640;
  wire _7471 = r1711 ^ r1832;
  wire _7472 = _7470 ^ _7471;
  wire _7473 = r1834 ^ r1892;
  wire _7474 = r1909 ^ r1960;
  wire _7475 = _7473 ^ _7474;
  wire _7476 = _7472 ^ _7475;
  wire _7477 = r1983 ^ r1995;
  wire _7478 = r2008 ^ r2013;
  wire _7479 = _7477 ^ _7478;
  wire _7480 = r2020 ^ r2028;
  wire _7481 = r2039 ^ r2047;
  wire _7482 = _7480 ^ _7481;
  wire _7483 = _7479 ^ _7482;
  wire _7484 = _7476 ^ _7483;
  wire _7485 = _7469 ^ _7484;
  wire _7486 = _7454 | _7485;
  wire _7487 = r12 ^ r84;
  wire _7488 = r131 ^ r177;
  wire _7489 = _7487 ^ _7488;
  wire _7490 = r265 ^ r315;
  wire _7491 = r386 ^ r394;
  wire _7492 = _7490 ^ _7491;
  wire _7493 = _7489 ^ _7492;
  wire _7494 = r463 ^ r528;
  wire _7495 = r603 ^ r638;
  wire _7496 = _7494 ^ _7495;
  wire _7497 = r768 ^ r809;
  wire _7498 = r886 ^ r937;
  wire _7499 = _7497 ^ _7498;
  wire _7500 = _7496 ^ _7499;
  wire _7501 = _7493 ^ _7500;
  wire _7502 = r968 ^ r1041;
  wire _7503 = r1147 ^ r1202;
  wire _7504 = _7502 ^ _7503;
  wire _7505 = r1272 ^ r1310;
  wire _7506 = r1383 ^ r1452;
  wire _7507 = _7505 ^ _7506;
  wire _7508 = _7504 ^ _7507;
  wire _7509 = r1468 ^ r1478;
  wire _7510 = r1498 ^ r1662;
  wire _7511 = _7509 ^ _7510;
  wire _7512 = r1753 ^ r1791;
  wire _7513 = r1808 ^ r1853;
  wire _7514 = _7512 ^ _7513;
  wire _7515 = _7511 ^ _7514;
  wire _7516 = _7508 ^ _7515;
  wire _7517 = _7501 ^ _7516;
  wire _7518 = r100 ^ r144;
  wire _7519 = r196 ^ r235;
  wire _7520 = _7518 ^ _7519;
  wire _7521 = r336 ^ r420;
  wire _7522 = r460 ^ r619;
  wire _7523 = _7521 ^ _7522;
  wire _7524 = _7520 ^ _7523;
  wire _7525 = r704 ^ r736;
  wire _7526 = r805 ^ r842;
  wire _7527 = _7525 ^ _7526;
  wire _7528 = r921 ^ r964;
  wire _7529 = r1042 ^ r1152;
  wire _7530 = _7528 ^ _7529;
  wire _7531 = _7527 ^ _7530;
  wire _7532 = _7524 ^ _7531;
  wire _7533 = r1170 ^ r1327;
  wire _7534 = r1349 ^ r1416;
  wire _7535 = _7533 ^ _7534;
  wire _7536 = r1427 ^ r1497;
  wire _7537 = r1523 ^ r1558;
  wire _7538 = _7536 ^ _7537;
  wire _7539 = _7535 ^ _7538;
  wire _7540 = r1799 ^ r1818;
  wire _7541 = r1826 ^ r1830;
  wire _7542 = _7540 ^ _7541;
  wire _7543 = r1837 ^ r1838;
  wire _7544 = r1867 ^ r1889;
  wire _7545 = _7543 ^ _7544;
  wire _7546 = _7542 ^ _7545;
  wire _7547 = _7539 ^ _7546;
  wire _7548 = _7532 ^ _7547;
  wire _7549 = _7517 | _7548;
  wire _7550 = _7486 | _7549;
  wire _7551 = r11 ^ r104;
  wire _7552 = r155 ^ r221;
  wire _7553 = _7551 ^ _7552;
  wire _7554 = r271 ^ r310;
  wire _7555 = r390 ^ r410;
  wire _7556 = _7554 ^ _7555;
  wire _7557 = _7553 ^ _7556;
  wire _7558 = r475 ^ r527;
  wire _7559 = r608 ^ r653;
  wire _7560 = _7558 ^ _7559;
  wire _7561 = r698 ^ r742;
  wire _7562 = r810 ^ r851;
  wire _7563 = _7561 ^ _7562;
  wire _7564 = _7560 ^ _7563;
  wire _7565 = _7557 ^ _7564;
  wire _7566 = r927 ^ r984;
  wire _7567 = r1020 ^ r1083;
  wire _7568 = _7566 ^ _7567;
  wire _7569 = r1244 ^ r1278;
  wire _7570 = r1293 ^ r1350;
  wire _7571 = _7569 ^ _7570;
  wire _7572 = _7568 ^ _7571;
  wire _7573 = r1393 ^ r1429;
  wire _7574 = r1514 ^ r1517;
  wire _7575 = _7573 ^ _7574;
  wire _7576 = r1592 ^ r1636;
  wire _7577 = r1669 ^ r1782;
  wire _7578 = _7576 ^ _7577;
  wire _7579 = _7575 ^ _7578;
  wire _7580 = _7572 ^ _7579;
  wire _7581 = _7565 ^ _7580;
  wire _7582 = r10 ^ r110;
  wire _7583 = r125 ^ r228;
  wire _7584 = _7582 ^ _7583;
  wire _7585 = r322 ^ r334;
  wire _7586 = r399 ^ r467;
  wire _7587 = _7585 ^ _7586;
  wire _7588 = _7584 ^ _7587;
  wire _7589 = r522 ^ r584;
  wire _7590 = r654 ^ r680;
  wire _7591 = _7589 ^ _7590;
  wire _7592 = r726 ^ r800;
  wire _7593 = r878 ^ r893;
  wire _7594 = _7592 ^ _7593;
  wire _7595 = _7591 ^ _7594;
  wire _7596 = _7588 ^ _7595;
  wire _7597 = r947 ^ r1012;
  wire _7598 = r1088 ^ r1151;
  wire _7599 = _7597 ^ _7598;
  wire _7600 = r1200 ^ r1242;
  wire _7601 = r1301 ^ r1382;
  wire _7602 = _7600 ^ _7601;
  wire _7603 = _7599 ^ _7602;
  wire _7604 = r1413 ^ r1444;
  wire _7605 = r1574 ^ r1612;
  wire _7606 = _7604 ^ _7605;
  wire _7607 = r1650 ^ r1695;
  wire _7608 = r1789 ^ r1854;
  wire _7609 = _7607 ^ _7608;
  wire _7610 = _7606 ^ _7609;
  wire _7611 = _7603 ^ _7610;
  wire _7612 = _7596 ^ _7611;
  wire _7613 = _7581 | _7612;
  wire _7614 = r9 ^ r103;
  wire _7615 = r113 ^ r179;
  wire _7616 = _7614 ^ _7615;
  wire _7617 = r236 ^ r294;
  wire _7618 = r383 ^ r416;
  wire _7619 = _7617 ^ _7618;
  wire _7620 = _7616 ^ _7619;
  wire _7621 = r498 ^ r507;
  wire _7622 = r582 ^ r641;
  wire _7623 = _7621 ^ _7622;
  wire _7624 = r687 ^ r728;
  wire _7625 = r824 ^ r837;
  wire _7626 = _7624 ^ _7625;
  wire _7627 = _7623 ^ _7626;
  wire _7628 = _7620 ^ _7627;
  wire _7629 = r891 ^ r948;
  wire _7630 = r1028 ^ r1059;
  wire _7631 = _7629 ^ _7630;
  wire _7632 = r1079 ^ r1145;
  wire _7633 = r1182 ^ r1297;
  wire _7634 = _7632 ^ _7633;
  wire _7635 = _7631 ^ _7634;
  wire _7636 = r1374 ^ r1469;
  wire _7637 = r1521 ^ r1547;
  wire _7638 = _7636 ^ _7637;
  wire _7639 = r1593 ^ r1643;
  wire _7640 = r1715 ^ r1783;
  wire _7641 = _7639 ^ _7640;
  wire _7642 = _7638 ^ _7641;
  wire _7643 = _7635 ^ _7642;
  wire _7644 = _7628 ^ _7643;
  wire _7645 = r8 ^ r98;
  wire _7646 = r158 ^ r223;
  wire _7647 = _7645 ^ _7646;
  wire _7648 = r264 ^ r284;
  wire _7649 = r360 ^ r392;
  wire _7650 = _7648 ^ _7649;
  wire _7651 = _7647 ^ _7650;
  wire _7652 = r452 ^ r513;
  wire _7653 = r596 ^ r620;
  wire _7654 = _7652 ^ _7653;
  wire _7655 = r710 ^ r752;
  wire _7656 = r829 ^ r866;
  wire _7657 = _7655 ^ _7656;
  wire _7658 = _7654 ^ _7657;
  wire _7659 = _7651 ^ _7658;
  wire _7660 = r926 ^ r983;
  wire _7661 = r1032 ^ r1099;
  wire _7662 = _7660 ^ _7661;
  wire _7663 = r1127 ^ r1185;
  wire _7664 = r1424 ^ r1572;
  wire _7665 = _7663 ^ _7664;
  wire _7666 = _7662 ^ _7665;
  wire _7667 = r1587 ^ r1717;
  wire _7668 = r1794 ^ r1811;
  wire _7669 = _7667 ^ _7668;
  wire _7670 = r1814 ^ r1817;
  wire _7671 = r1866 ^ r1890;
  wire _7672 = _7670 ^ _7671;
  wire _7673 = _7669 ^ _7672;
  wire _7674 = _7666 ^ _7673;
  wire _7675 = _7659 ^ _7674;
  wire _7676 = _7644 | _7675;
  wire _7677 = _7613 | _7676;
  wire _7678 = _7550 | _7677;
  wire _7679 = _7423 | _7678;
  wire _7680 = r7 ^ r81;
  wire _7681 = r116 ^ r210;
  wire _7682 = _7680 ^ _7681;
  wire _7683 = r277 ^ r324;
  wire _7684 = r343 ^ r444;
  wire _7685 = _7683 ^ _7684;
  wire _7686 = _7682 ^ _7685;
  wire _7687 = r502 ^ r534;
  wire _7688 = r589 ^ r637;
  wire _7689 = _7687 ^ _7688;
  wire _7690 = r708 ^ r734;
  wire _7691 = r814 ^ r845;
  wire _7692 = _7690 ^ _7691;
  wire _7693 = _7689 ^ _7692;
  wire _7694 = _7686 ^ _7693;
  wire _7695 = r907 ^ r975;
  wire _7696 = r1105 ^ r1113;
  wire _7697 = _7695 ^ _7696;
  wire _7698 = r1134 ^ r1171;
  wire _7699 = r1259 ^ r1339;
  wire _7700 = _7698 ^ _7699;
  wire _7701 = _7697 ^ _7700;
  wire _7702 = r1394 ^ r1437;
  wire _7703 = r1505 ^ r1605;
  wire _7704 = _7702 ^ _7703;
  wire _7705 = r1686 ^ r1703;
  wire _7706 = r1806 ^ r1855;
  wire _7707 = _7705 ^ _7706;
  wire _7708 = _7704 ^ _7707;
  wire _7709 = _7701 ^ _7708;
  wire _7710 = _7694 ^ _7709;
  wire _7711 = r6 ^ r88;
  wire _7712 = r175 ^ r250;
  wire _7713 = _7711 ^ _7712;
  wire _7714 = r285 ^ r355;
  wire _7715 = r403 ^ r449;
  wire _7716 = _7714 ^ _7715;
  wire _7717 = _7713 ^ _7716;
  wire _7718 = r532 ^ r565;
  wire _7719 = r685 ^ r745;
  wire _7720 = _7718 ^ _7719;
  wire _7721 = r816 ^ r992;
  wire _7722 = r1031 ^ r1090;
  wire _7723 = _7721 ^ _7722;
  wire _7724 = _7720 ^ _7723;
  wire _7725 = _7717 ^ _7724;
  wire _7726 = r1157 ^ r1168;
  wire _7727 = r1201 ^ r1245;
  wire _7728 = _7726 ^ _7727;
  wire _7729 = r1388 ^ r1463;
  wire _7730 = r1536 ^ r1548;
  wire _7731 = _7729 ^ _7730;
  wire _7732 = _7728 ^ _7731;
  wire _7733 = r1624 ^ r1690;
  wire _7734 = r1802 ^ r1891;
  wire _7735 = _7733 ^ _7734;
  wire _7736 = r1893 ^ r1901;
  wire _7737 = r1941 ^ r1947;
  wire _7738 = _7736 ^ _7737;
  wire _7739 = _7735 ^ _7738;
  wire _7740 = _7732 ^ _7739;
  wire _7741 = _7725 ^ _7740;
  wire _7742 = _7710 | _7741;
  wire _7743 = r5 ^ r108;
  wire _7744 = r146 ^ r203;
  wire _7745 = _7743 ^ _7744;
  wire _7746 = r231 ^ r303;
  wire _7747 = r367 ^ r396;
  wire _7748 = _7746 ^ _7747;
  wire _7749 = _7745 ^ _7748;
  wire _7750 = r495 ^ r511;
  wire _7751 = r575 ^ r650;
  wire _7752 = _7750 ^ _7751;
  wire _7753 = r720 ^ r753;
  wire _7754 = r786 ^ r880;
  wire _7755 = _7753 ^ _7754;
  wire _7756 = _7752 ^ _7755;
  wire _7757 = _7749 ^ _7756;
  wire _7758 = r894 ^ r997;
  wire _7759 = r1003 ^ r1026;
  wire _7760 = _7758 ^ _7759;
  wire _7761 = r1092 ^ r1155;
  wire _7762 = r1319 ^ r1338;
  wire _7763 = _7761 ^ _7762;
  wire _7764 = _7760 ^ _7763;
  wire _7765 = r1471 ^ r1522;
  wire _7766 = r1596 ^ r1638;
  wire _7767 = _7765 ^ _7766;
  wire _7768 = r1666 ^ r1696;
  wire _7769 = r1786 ^ r1856;
  wire _7770 = _7768 ^ _7769;
  wire _7771 = _7767 ^ _7770;
  wire _7772 = _7764 ^ _7771;
  wire _7773 = _7757 ^ _7772;
  wire _7774 = r4 ^ r106;
  wire _7775 = r141 ^ r200;
  wire _7776 = _7774 ^ _7775;
  wire _7777 = r252 ^ r312;
  wire _7778 = r337 ^ r427;
  wire _7779 = _7777 ^ _7778;
  wire _7780 = _7776 ^ _7779;
  wire _7781 = r476 ^ r548;
  wire _7782 = r569 ^ r670;
  wire _7783 = _7781 ^ _7782;
  wire _7784 = r727 ^ r822;
  wire _7785 = r1009 ^ r1064;
  wire _7786 = _7784 ^ _7785;
  wire _7787 = _7783 ^ _7786;
  wire _7788 = _7780 ^ _7787;
  wire _7789 = r1132 ^ r1281;
  wire _7790 = r1335 ^ r1439;
  wire _7791 = _7789 ^ _7790;
  wire _7792 = r1503 ^ r1598;
  wire _7793 = r1675 ^ r1744;
  wire _7794 = _7792 ^ _7793;
  wire _7795 = _7791 ^ _7794;
  wire _7796 = r1764 ^ r1816;
  wire _7797 = r1872 ^ r1904;
  wire _7798 = _7796 ^ _7797;
  wire _7799 = r1927 ^ r1950;
  wire _7800 = r1968 ^ r1971;
  wire _7801 = _7799 ^ _7800;
  wire _7802 = _7798 ^ _7801;
  wire _7803 = _7795 ^ _7802;
  wire _7804 = _7788 ^ _7803;
  wire _7805 = _7773 | _7804;
  wire _7806 = _7742 | _7805;
  wire _7807 = r147 ^ r266;
  wire _7808 = r385 ^ r459;
  wire _7809 = _7807 ^ _7808;
  wire _7810 = r551 ^ r572;
  wire _7811 = r665 ^ r741;
  wire _7812 = _7810 ^ _7811;
  wire _7813 = _7809 ^ _7812;
  wire _7814 = r840 ^ r890;
  wire _7815 = r996 ^ r1016;
  wire _7816 = _7814 ^ _7815;
  wire _7817 = r1178 ^ r1269;
  wire _7818 = r1305 ^ r1371;
  wire _7819 = _7817 ^ _7818;
  wire _7820 = _7816 ^ _7819;
  wire _7821 = _7813 ^ _7820;
  wire _7822 = r1421 ^ r1482;
  wire _7823 = r1554 ^ r1609;
  wire _7824 = _7822 ^ _7823;
  wire _7825 = r1716 ^ r1807;
  wire _7826 = r1980 ^ r1986;
  wire _7827 = _7825 ^ _7826;
  wire _7828 = _7824 ^ _7827;
  wire _7829 = r1987 ^ r1992;
  wire _7830 = r1999 ^ r2011;
  wire _7831 = _7829 ^ _7830;
  wire _7832 = r2014 ^ r2024;
  wire _7833 = r2030 ^ r2038;
  wire _7834 = _7832 ^ _7833;
  wire _7835 = _7831 ^ _7834;
  wire _7836 = _7828 ^ _7835;
  wire _7837 = _7821 ^ _7836;
  wire _7838 = r3 ^ r66;
  wire _7839 = r136 ^ r207;
  wire _7840 = _7838 ^ _7839;
  wire _7841 = r262 ^ r313;
  wire _7842 = r370 ^ r431;
  wire _7843 = _7841 ^ _7842;
  wire _7844 = _7840 ^ _7843;
  wire _7845 = r471 ^ r535;
  wire _7846 = r562 ^ r686;
  wire _7847 = _7845 ^ _7846;
  wire _7848 = r769 ^ r787;
  wire _7849 = r862 ^ r918;
  wire _7850 = _7848 ^ _7849;
  wire _7851 = _7847 ^ _7850;
  wire _7852 = _7844 ^ _7851;
  wire _7853 = r991 ^ r1037;
  wire _7854 = r1109 ^ r1115;
  wire _7855 = _7853 ^ _7854;
  wire _7856 = r1203 ^ r1220;
  wire _7857 = r1254 ^ r1378;
  wire _7858 = _7856 ^ _7857;
  wire _7859 = _7855 ^ _7858;
  wire _7860 = r1418 ^ r1467;
  wire _7861 = r1528 ^ r1603;
  wire _7862 = _7860 ^ _7861;
  wire _7863 = r1637 ^ r1653;
  wire _7864 = r1759 ^ r1857;
  wire _7865 = _7863 ^ _7864;
  wire _7866 = _7862 ^ _7865;
  wire _7867 = _7859 ^ _7866;
  wire _7868 = _7852 ^ _7867;
  wire _7869 = _7837 | _7868;
  wire _7870 = r2 ^ r69;
  wire _7871 = r161 ^ r185;
  wire _7872 = _7870 ^ _7871;
  wire _7873 = r226 ^ r302;
  wire _7874 = r388 ^ r435;
  wire _7875 = _7873 ^ _7874;
  wire _7876 = _7872 ^ _7875;
  wire _7877 = r481 ^ r512;
  wire _7878 = r597 ^ r618;
  wire _7879 = _7877 ^ _7878;
  wire _7880 = r707 ^ r748;
  wire _7881 = r815 ^ r863;
  wire _7882 = _7880 ^ _7881;
  wire _7883 = _7879 ^ _7882;
  wire _7884 = _7876 ^ _7883;
  wire _7885 = r903 ^ r972;
  wire _7886 = r1035 ^ r1065;
  wire _7887 = _7885 ^ _7886;
  wire _7888 = r1158 ^ r1194;
  wire _7889 = r1222 ^ r1311;
  wire _7890 = _7888 ^ _7889;
  wire _7891 = _7887 ^ _7890;
  wire _7892 = r1345 ^ r1384;
  wire _7893 = r1524 ^ r1540;
  wire _7894 = _7892 ^ _7893;
  wire _7895 = r1630 ^ r1661;
  wire _7896 = r1709 ^ r1784;
  wire _7897 = _7895 ^ _7896;
  wire _7898 = _7894 ^ _7897;
  wire _7899 = _7891 ^ _7898;
  wire _7900 = _7884 ^ _7899;
  wire _7901 = r1 ^ r109;
  wire _7902 = r168 ^ r194;
  wire _7903 = _7901 ^ _7902;
  wire _7904 = r247 ^ r327;
  wire _7905 = r349 ^ r424;
  wire _7906 = _7904 ^ _7905;
  wire _7907 = _7903 ^ _7906;
  wire _7908 = r453 ^ r531;
  wire _7909 = r581 ^ r646;
  wire _7910 = _7908 ^ _7909;
  wire _7911 = r677 ^ r771;
  wire _7912 = r828 ^ r839;
  wire _7913 = _7911 ^ _7912;
  wire _7914 = _7910 ^ _7913;
  wire _7915 = _7907 ^ _7914;
  wire _7916 = r928 ^ r980;
  wire _7917 = r1014 ^ r1091;
  wire _7918 = _7916 ^ _7917;
  wire _7919 = r1133 ^ r1183;
  wire _7920 = r1271 ^ r1323;
  wire _7921 = _7919 ^ _7920;
  wire _7922 = _7918 ^ _7921;
  wire _7923 = r1333 ^ r1343;
  wire _7924 = r1447 ^ r1483;
  wire _7925 = _7923 ^ _7924;
  wire _7926 = r1646 ^ r1699;
  wire _7927 = r1755 ^ r1858;
  wire _7928 = _7926 ^ _7927;
  wire _7929 = _7925 ^ _7928;
  wire _7930 = _7922 ^ _7929;
  wire _7931 = _7915 ^ _7930;
  wire _7932 = _7900 | _7931;
  wire _7933 = _7869 | _7932;
  wire _7934 = _7806 | _7933;
  wire _7935 = r0 ^ r87;
  wire _7936 = r151 ^ r189;
  wire _7937 = _7935 ^ _7936;
  wire _7938 = r248 ^ r280;
  wire _7939 = r357 ^ r404;
  wire _7940 = _7938 ^ _7939;
  wire _7941 = _7937 ^ _7940;
  wire _7942 = r497 ^ r559;
  wire _7943 = r592 ^ r643;
  wire _7944 = _7942 ^ _7943;
  wire _7945 = r717 ^ r729;
  wire _7946 = r801 ^ r831;
  wire _7947 = _7945 ^ _7946;
  wire _7948 = _7944 ^ _7947;
  wire _7949 = _7941 ^ _7948;
  wire _7950 = r920 ^ r1002;
  wire _7951 = r1051 ^ r1104;
  wire _7952 = _7950 ^ _7951;
  wire _7953 = r1154 ^ r1199;
  wire _7954 = r1257 ^ r1279;
  wire _7955 = _7953 ^ _7954;
  wire _7956 = _7952 ^ _7955;
  wire _7957 = r1377 ^ r1401;
  wire _7958 = r1431 ^ r1490;
  wire _7959 = _7957 ^ _7958;
  wire _7960 = r1529 ^ r1597;
  wire _7961 = r1658 ^ r1785;
  wire _7962 = _7960 ^ _7961;
  wire _7963 = _7959 ^ _7962;
  wire _7964 = _7956 ^ _7963;
  wire _7965 = _7949 ^ _7964;
  wire _7966 = r152 ^ r192;
  wire _7967 = r225 ^ r317;
  wire _7968 = _7966 ^ _7967;
  wire _7969 = r353 ^ r443;
  wire _7970 = r544 ^ r657;
  wire _7971 = _7969 ^ _7970;
  wire _7972 = _7968 ^ _7971;
  wire _7973 = r688 ^ r725;
  wire _7974 = r782 ^ r849;
  wire _7975 = _7973 ^ _7974;
  wire _7976 = r908 ^ r1000;
  wire _7977 = r1054 ^ r1124;
  wire _7978 = _7976 ^ _7977;
  wire _7979 = _7975 ^ _7978;
  wire _7980 = _7972 ^ _7979;
  wire _7981 = r1175 ^ r1304;
  wire _7982 = r1390 ^ r1462;
  wire _7983 = _7981 ^ _7982;
  wire _7984 = r1520 ^ r1557;
  wire _7985 = r1648 ^ r1723;
  wire _7986 = _7984 ^ _7985;
  wire _7987 = _7983 ^ _7986;
  wire _7988 = r1735 ^ r1736;
  wire _7989 = r1741 ^ r1751;
  wire _7990 = _7988 ^ _7989;
  wire _7991 = r1822 ^ r1840;
  wire _7992 = r1883 ^ r1911;
  wire _7993 = _7991 ^ _7992;
  wire _7994 = _7990 ^ _7993;
  wire _7995 = _7987 ^ _7994;
  wire _7996 = _7980 ^ _7995;
  wire _7997 = _7965 | _7996;
  wire _7998 = r79 ^ r120;
  wire _7999 = r184 ^ r319;
  wire _8000 = _7998 ^ _7999;
  wire _8001 = r358 ^ r400;
  wire _8002 = r500 ^ r514;
  wire _8003 = _8001 ^ _8002;
  wire _8004 = _8000 ^ _8003;
  wire _8005 = r576 ^ r652;
  wire _8006 = r679 ^ r744;
  wire _8007 = _8005 ^ _8006;
  wire _8008 = r803 ^ r854;
  wire _8009 = r925 ^ r978;
  wire _8010 = _8008 ^ _8009;
  wire _8011 = _8007 ^ _8010;
  wire _8012 = _8004 ^ _8011;
  wire _8013 = r1038 ^ r1173;
  wire _8014 = r1250 ^ r1318;
  wire _8015 = _8013 ^ _8014;
  wire _8016 = r1360 ^ r1405;
  wire _8017 = r1448 ^ r1489;
  wire _8018 = _8016 ^ _8017;
  wire _8019 = _8015 ^ _8018;
  wire _8020 = r1508 ^ r1512;
  wire _8021 = r1560 ^ r1588;
  wire _8022 = _8020 ^ _8021;
  wire _8023 = r1676 ^ r1762;
  wire _8024 = r1928 ^ r1933;
  wire _8025 = _8023 ^ _8024;
  wire _8026 = _8022 ^ _8025;
  wire _8027 = _8019 ^ _8026;
  wire _8028 = _8012 ^ _8027;
  wire _8029 = r62 ^ r159;
  wire _8030 = r215 ^ r289;
  wire _8031 = _8029 ^ _8030;
  wire _8032 = r348 ^ r409;
  wire _8033 = r464 ^ r506;
  wire _8034 = _8032 ^ _8033;
  wire _8035 = _8031 ^ _8034;
  wire _8036 = r564 ^ r626;
  wire _8037 = r721 ^ r765;
  wire _8038 = _8036 ^ _8037;
  wire _8039 = r817 ^ r899;
  wire _8040 = r957 ^ r1015;
  wire _8041 = _8039 ^ _8040;
  wire _8042 = _8038 ^ _8041;
  wire _8043 = _8035 ^ _8042;
  wire _8044 = r1081 ^ r1135;
  wire _8045 = r1187 ^ r1221;
  wire _8046 = _8044 ^ _8045;
  wire _8047 = r1247 ^ r1294;
  wire _8048 = r1346 ^ r1409;
  wire _8049 = _8047 ^ _8048;
  wire _8050 = _8046 ^ _8049;
  wire _8051 = r1477 ^ r1501;
  wire _8052 = r1570 ^ r1644;
  wire _8053 = _8051 ^ _8052;
  wire _8054 = r1665 ^ r1722;
  wire _8055 = r1793 ^ r1859;
  wire _8056 = _8054 ^ _8055;
  wire _8057 = _8053 ^ _8056;
  wire _8058 = _8050 ^ _8057;
  wire _8059 = _8043 ^ _8058;
  wire _8060 = _8028 | _8059;
  wire _8061 = _7997 | _8060;
  wire _8062 = r89 ^ r112;
  wire _8063 = r199 ^ r239;
  wire _8064 = _8062 ^ _8063;
  wire _8065 = r325 ^ r373;
  wire _8066 = r438 ^ r473;
  wire _8067 = _8065 ^ _8066;
  wire _8068 = _8064 ^ _8067;
  wire _8069 = r549 ^ r605;
  wire _8070 = r635 ^ r684;
  wire _8071 = _8069 ^ _8070;
  wire _8072 = r766 ^ r813;
  wire _8073 = r853 ^ r896;
  wire _8074 = _8072 ^ _8073;
  wire _8075 = _8071 ^ _8074;
  wire _8076 = _8068 ^ _8075;
  wire _8077 = r960 ^ r1034;
  wire _8078 = r1093 ^ r1126;
  wire _8079 = _8077 ^ _8078;
  wire _8080 = r1180 ^ r1262;
  wire _8081 = r1326 ^ r1398;
  wire _8082 = _8080 ^ _8081;
  wire _8083 = _8079 ^ _8082;
  wire _8084 = r1563 ^ r1589;
  wire _8085 = r1671 ^ r1721;
  wire _8086 = _8084 ^ _8085;
  wire _8087 = r1731 ^ r1742;
  wire _8088 = r1805 ^ r1860;
  wire _8089 = _8087 ^ _8088;
  wire _8090 = _8086 ^ _8089;
  wire _8091 = _8083 ^ _8090;
  wire _8092 = _8076 ^ _8091;
  wire _8093 = r80 ^ r121;
  wire _8094 = r211 ^ r279;
  wire _8095 = _8093 ^ _8094;
  wire _8096 = r283 ^ r380;
  wire _8097 = r426 ^ r468;
  wire _8098 = _8096 ^ _8097;
  wire _8099 = _8095 ^ _8098;
  wire _8100 = r510 ^ r567;
  wire _8101 = r629 ^ r714;
  wire _8102 = _8100 ^ _8101;
  wire _8103 = r743 ^ r778;
  wire _8104 = r847 ^ r912;
  wire _8105 = _8103 ^ _8104;
  wire _8106 = _8102 ^ _8105;
  wire _8107 = _8099 ^ _8106;
  wire _8108 = r944 ^ r1007;
  wire _8109 = r1060 ^ r1114;
  wire _8110 = _8108 ^ _8109;
  wire _8111 = r1211 ^ r1255;
  wire _8112 = r1296 ^ r1342;
  wire _8113 = _8111 ^ _8112;
  wire _8114 = _8110 ^ _8113;
  wire _8115 = r1541 ^ r1567;
  wire _8116 = r1599 ^ r1635;
  wire _8117 = _8115 ^ _8116;
  wire _8118 = r1681 ^ r1719;
  wire _8119 = r1768 ^ r1861;
  wire _8120 = _8118 ^ _8119;
  wire _8121 = _8117 ^ _8120;
  wire _8122 = _8114 ^ _8121;
  wire _8123 = _8107 ^ _8122;
  wire _8124 = _8092 | _8123;
  wire _8125 = r67 ^ r222;
  wire _8126 = r238 ^ r290;
  wire _8127 = _8125 ^ _8126;
  wire _8128 = r362 ^ r412;
  wire _8129 = r474 ^ r540;
  wire _8130 = _8128 ^ _8129;
  wire _8131 = _8127 ^ _8130;
  wire _8132 = r586 ^ r632;
  wire _8133 = r712 ^ r735;
  wire _8134 = _8132 ^ _8133;
  wire _8135 = r798 ^ r884;
  wire _8136 = r905 ^ r979;
  wire _8137 = _8135 ^ _8136;
  wire _8138 = _8134 ^ _8137;
  wire _8139 = _8131 ^ _8138;
  wire _8140 = r1047 ^ r1107;
  wire _8141 = r1131 ^ r1232;
  wire _8142 = _8140 ^ _8141;
  wire _8143 = r1306 ^ r1369;
  wire _8144 = r1417 ^ r1443;
  wire _8145 = _8143 ^ _8144;
  wire _8146 = _8142 ^ _8145;
  wire _8147 = r1456 ^ r1493;
  wire _8148 = r1516 ^ r1720;
  wire _8149 = _8147 ^ _8148;
  wire _8150 = r1733 ^ r1754;
  wire _8151 = r1923 ^ r1926;
  wire _8152 = _8150 ^ _8151;
  wire _8153 = _8149 ^ _8152;
  wire _8154 = _8146 ^ _8153;
  wire _8155 = _8139 ^ _8154;
  wire _8156 = r52 ^ r86;
  wire _8157 = r167 ^ r195;
  wire _8158 = _8156 ^ _8157;
  wire _8159 = r233 ^ r318;
  wire _8160 = r364 ^ r429;
  wire _8161 = _8159 ^ _8160;
  wire _8162 = _8158 ^ _8161;
  wire _8163 = r537 ^ r594;
  wire _8164 = r672 ^ r751;
  wire _8165 = _8163 ^ _8164;
  wire _8166 = r799 ^ r934;
  wire _8167 = r1017 ^ r1077;
  wire _8168 = _8166 ^ _8167;
  wire _8169 = _8165 ^ _8168;
  wire _8170 = _8162 ^ _8169;
  wire _8171 = r1110 ^ r1163;
  wire _8172 = r1214 ^ r1432;
  wire _8173 = _8171 ^ _8172;
  wire _8174 = r1465 ^ r1538;
  wire _8175 = r1691 ^ r1787;
  wire _8176 = _8174 ^ _8175;
  wire _8177 = _8173 ^ _8176;
  wire _8178 = r1836 ^ r1879;
  wire _8179 = r1897 ^ r1906;
  wire _8180 = _8178 ^ _8179;
  wire _8181 = r1929 ^ r1936;
  wire _8182 = r1961 ^ r1979;
  wire _8183 = _8181 ^ _8182;
  wire _8184 = _8180 ^ _8183;
  wire _8185 = _8177 ^ _8184;
  wire _8186 = _8170 ^ _8185;
  wire _8187 = _8155 | _8186;
  wire _8188 = _8124 | _8187;
  wire _8189 = _8061 | _8188;
  wire _8190 = _7934 | _8189;
  wire _8191 = _7679 | _8190;
  wire _8192 = _7168 | _8191;
  wire _8193 = _6145 | _8192;
  wire _8194 = _4098 | _8193;
  wire _8195 = r53 ^ r106;
  wire _8196 = r127 ^ r242;
  wire _8197 = _8195 ^ _8196;
  wire _8198 = r296 ^ r339;
  wire _8199 = r455 ^ r532;
  wire _8200 = _8198 ^ _8199;
  wire _8201 = _8197 ^ _8200;
  wire _8202 = r638 ^ r708;
  wire _8203 = r760 ^ r793;
  wire _8204 = _8202 ^ _8203;
  wire _8205 = r891 ^ r1000;
  wire _8206 = r1035 ^ r1071;
  wire _8207 = _8205 ^ _8206;
  wire _8208 = _8204 ^ _8207;
  wire _8209 = _8201 ^ _8208;
  wire _8210 = r1155 ^ r1242;
  wire _8211 = r1285 ^ r1343;
  wire _8212 = _8210 ^ _8211;
  wire _8213 = r1414 ^ r1454;
  wire _8214 = r1517 ^ r1747;
  wire _8215 = _8213 ^ _8214;
  wire _8216 = _8212 ^ _8215;
  wire _8217 = r1780 ^ r1846;
  wire _8218 = r1929 ^ r1959;
  wire _8219 = _8217 ^ _8218;
  wire _8220 = r1962 ^ r1990;
  wire _8221 = r1995 ^ r1997;
  wire _8222 = _8220 ^ _8221;
  wire _8223 = _8219 ^ _8222;
  wire _8224 = _8216 ^ _8223;
  wire _8225 = _8209 ^ _8224;
  wire _8226 = r51 ^ r85;
  wire _8227 = r166 ^ r194;
  wire _8228 = _8226 ^ _8227;
  wire _8229 = r232 ^ r317;
  wire _8230 = r363 ^ r428;
  wire _8231 = _8229 ^ _8230;
  wire _8232 = _8228 ^ _8231;
  wire _8233 = r463 ^ r536;
  wire _8234 = r593 ^ r624;
  wire _8235 = _8233 ^ _8234;
  wire _8236 = r671 ^ r750;
  wire _8237 = r798 ^ r835;
  wire _8238 = _8236 ^ _8237;
  wire _8239 = _8235 ^ _8238;
  wire _8240 = _8232 ^ _8239;
  wire _8241 = r933 ^ r999;
  wire _8242 = r1016 ^ r1076;
  wire _8243 = _8241 ^ _8242;
  wire _8244 = r1108 ^ r1162;
  wire _8245 = r1213 ^ r1240;
  wire _8246 = _8244 ^ _8245;
  wire _8247 = _8243 ^ _8246;
  wire _8248 = r1303 ^ r1354;
  wire _8249 = r1431 ^ r1464;
  wire _8250 = _8248 ^ _8249;
  wire _8251 = r1484 ^ r1652;
  wire _8252 = r1690 ^ r1786;
  wire _8253 = _8251 ^ _8252;
  wire _8254 = _8250 ^ _8253;
  wire _8255 = _8247 ^ _8254;
  wire _8256 = _8240 ^ _8255;
  wire _8257 = _8225 | _8256;
  wire _8258 = r50 ^ r57;
  wire _8259 = r331 ^ r553;
  wire _8260 = _8258 ^ _8259;
  wire _8261 = r589 ^ r657;
  wire _8262 = r718 ^ r755;
  wire _8263 = _8261 ^ _8262;
  wire _8264 = _8260 ^ _8263;
  wire _8265 = r829 ^ r857;
  wire _8266 = r943 ^ r968;
  wire _8267 = _8265 ^ _8266;
  wire _8268 = r1077 ^ r1159;
  wire _8269 = r1215 ^ r1222;
  wire _8270 = _8268 ^ _8269;
  wire _8271 = _8267 ^ _8270;
  wire _8272 = _8264 ^ _8271;
  wire _8273 = r1320 ^ r1378;
  wire _8274 = r1547 ^ r1574;
  wire _8275 = _8273 ^ _8274;
  wire _8276 = r1632 ^ r1682;
  wire _8277 = r1770 ^ r1778;
  wire _8278 = _8276 ^ _8277;
  wire _8279 = _8275 ^ _8278;
  wire _8280 = r1801 ^ r1834;
  wire _8281 = r1884 ^ r1901;
  wire _8282 = _8280 ^ _8281;
  wire _8283 = r1921 ^ r1922;
  wire _8284 = r1945 ^ r1954;
  wire _8285 = _8283 ^ _8284;
  wire _8286 = _8282 ^ _8285;
  wire _8287 = _8279 ^ _8286;
  wire _8288 = _8272 ^ _8287;
  wire _8289 = r54 ^ r114;
  wire _8290 = r274 ^ r303;
  wire _8291 = _8289 ^ _8290;
  wire _8292 = r370 ^ r491;
  wire _8293 = r545 ^ r594;
  wire _8294 = _8292 ^ _8293;
  wire _8295 = _8291 ^ _8294;
  wire _8296 = r641 ^ r694;
  wire _8297 = r822 ^ r856;
  wire _8298 = _8296 ^ _8297;
  wire _8299 = r937 ^ r952;
  wire _8300 = r1051 ^ r1105;
  wire _8301 = _8299 ^ _8300;
  wire _8302 = _8298 ^ _8301;
  wire _8303 = _8295 ^ _8302;
  wire _8304 = r1117 ^ r1207;
  wire _8305 = r1218 ^ r1238;
  wire _8306 = _8304 ^ _8305;
  wire _8307 = r1289 ^ r1499;
  wire _8308 = r1584 ^ r1615;
  wire _8309 = _8307 ^ _8308;
  wire _8310 = _8306 ^ _8309;
  wire _8311 = r1728 ^ r1735;
  wire _8312 = r1738 ^ r1833;
  wire _8313 = _8311 ^ _8312;
  wire _8314 = r1844 ^ r1970;
  wire _8315 = r1981 ^ r1986;
  wire _8316 = _8314 ^ _8315;
  wire _8317 = _8313 ^ _8316;
  wire _8318 = _8310 ^ _8317;
  wire _8319 = _8303 ^ _8318;
  wire _8320 = _8288 | _8319;
  wire _8321 = _8257 | _8320;
  wire _8322 = r49 ^ r71;
  wire _8323 = r138 ^ r186;
  wire _8324 = _8322 ^ _8323;
  wire _8325 = r243 ^ r383;
  wire _8326 = r396 ^ r584;
  wire _8327 = _8325 ^ _8326;
  wire _8328 = _8324 ^ _8327;
  wire _8329 = r754 ^ r833;
  wire _8330 = r941 ^ r980;
  wire _8331 = _8329 ^ _8330;
  wire _8332 = r1013 ^ r1187;
  wire _8333 = r1228 ^ r1290;
  wire _8334 = _8332 ^ _8333;
  wire _8335 = _8331 ^ _8334;
  wire _8336 = _8328 ^ _8335;
  wire _8337 = r1399 ^ r1437;
  wire _8338 = r1463 ^ r1618;
  wire _8339 = _8337 ^ _8338;
  wire _8340 = r1718 ^ r1765;
  wire _8341 = r1771 ^ r1822;
  wire _8342 = _8340 ^ _8341;
  wire _8343 = _8339 ^ _8342;
  wire _8344 = r1857 ^ r1943;
  wire _8345 = r1963 ^ r1988;
  wire _8346 = _8344 ^ _8345;
  wire _8347 = r2015 ^ r2020;
  wire _8348 = r2023 ^ r2030;
  wire _8349 = _8347 ^ _8348;
  wire _8350 = _8346 ^ _8349;
  wire _8351 = _8343 ^ _8350;
  wire _8352 = _8336 ^ _8351;
  wire _8353 = r48 ^ r63;
  wire _8354 = r152 ^ r204;
  wire _8355 = _8353 ^ _8354;
  wire _8356 = r305 ^ r333;
  wire _8357 = r401 ^ r477;
  wire _8358 = _8356 ^ _8357;
  wire _8359 = _8355 ^ _8358;
  wire _8360 = r528 ^ r607;
  wire _8361 = r698 ^ r777;
  wire _8362 = _8360 ^ _8361;
  wire _8363 = r789 ^ r868;
  wire _8364 = r970 ^ r1042;
  wire _8365 = _8363 ^ _8364;
  wire _8366 = _8362 ^ _8365;
  wire _8367 = _8359 ^ _8366;
  wire _8368 = r1062 ^ r1141;
  wire _8369 = r1171 ^ r1262;
  wire _8370 = _8368 ^ _8369;
  wire _8371 = r1319 ^ r1375;
  wire _8372 = r1493 ^ r1549;
  wire _8373 = _8371 ^ _8372;
  wire _8374 = _8370 ^ _8373;
  wire _8375 = r1570 ^ r1603;
  wire _8376 = r1672 ^ r1704;
  wire _8377 = _8375 ^ _8376;
  wire _8378 = r1761 ^ r1842;
  wire _8379 = r1874 ^ r1891;
  wire _8380 = _8378 ^ _8379;
  wire _8381 = _8377 ^ _8380;
  wire _8382 = _8374 ^ _8381;
  wire _8383 = _8367 ^ _8382;
  wire _8384 = _8352 | _8383;
  wire _8385 = r47 ^ r95;
  wire _8386 = r149 ^ r212;
  wire _8387 = _8385 ^ _8386;
  wire _8388 = r319 ^ r362;
  wire _8389 = r392 ^ r503;
  wire _8390 = _8388 ^ _8389;
  wire _8391 = _8387 ^ _8390;
  wire _8392 = r522 ^ r613;
  wire _8393 = r635 ^ r702;
  wire _8394 = _8392 ^ _8393;
  wire _8395 = r731 ^ r830;
  wire _8396 = r871 ^ r912;
  wire _8397 = _8395 ^ _8396;
  wire _8398 = _8394 ^ _8397;
  wire _8399 = _8391 ^ _8398;
  wire _8400 = r957 ^ r1039;
  wire _8401 = r1067 ^ r1152;
  wire _8402 = _8400 ^ _8401;
  wire _8403 = r1183 ^ r1245;
  wire _8404 = r1311 ^ r1350;
  wire _8405 = _8403 ^ _8404;
  wire _8406 = _8402 ^ _8405;
  wire _8407 = r1402 ^ r1480;
  wire _8408 = r1500 ^ r1559;
  wire _8409 = _8407 ^ _8408;
  wire _8410 = r1633 ^ r1700;
  wire _8411 = r1807 ^ r1862;
  wire _8412 = _8410 ^ _8411;
  wire _8413 = _8409 ^ _8412;
  wire _8414 = _8406 ^ _8413;
  wire _8415 = _8399 ^ _8414;
  wire _8416 = r46 ^ r104;
  wire _8417 = r169 ^ r207;
  wire _8418 = _8416 ^ _8417;
  wire _8419 = r253 ^ r315;
  wire _8420 = r378 ^ r414;
  wire _8421 = _8419 ^ _8420;
  wire _8422 = _8418 ^ _8421;
  wire _8423 = r525 ^ r598;
  wire _8424 = r691 ^ r738;
  wire _8425 = _8423 ^ _8424;
  wire _8426 = r788 ^ r858;
  wire _8427 = r894 ^ r976;
  wire _8428 = _8426 ^ _8427;
  wire _8429 = _8425 ^ _8428;
  wire _8430 = _8422 ^ _8429;
  wire _8431 = r1056 ^ r1145;
  wire _8432 = r1257 ^ r1347;
  wire _8433 = _8431 ^ _8432;
  wire _8434 = r1492 ^ r1509;
  wire _8435 = r1526 ^ r1554;
  wire _8436 = _8434 ^ _8435;
  wire _8437 = _8433 ^ _8436;
  wire _8438 = r1576 ^ r1673;
  wire _8439 = r1743 ^ r1840;
  wire _8440 = _8438 ^ _8439;
  wire _8441 = r1841 ^ r1905;
  wire _8442 = r1971 ^ r1978;
  wire _8443 = _8441 ^ _8442;
  wire _8444 = _8440 ^ _8443;
  wire _8445 = _8437 ^ _8444;
  wire _8446 = _8430 ^ _8445;
  wire _8447 = _8415 | _8446;
  wire _8448 = _8384 | _8447;
  wire _8449 = _8321 | _8448;
  wire _8450 = r45 ^ r98;
  wire _8451 = r132 ^ r213;
  wire _8452 = _8450 ^ _8451;
  wire _8453 = r256 ^ r281;
  wire _8454 = r349 ^ r421;
  wire _8455 = _8453 ^ _8454;
  wire _8456 = _8452 ^ _8455;
  wire _8457 = r495 ^ r600;
  wire _8458 = r666 ^ r672;
  wire _8459 = _8457 ^ _8458;
  wire _8460 = r761 ^ r783;
  wire _8461 = r834 ^ r908;
  wire _8462 = _8460 ^ _8461;
  wire _8463 = _8459 ^ _8462;
  wire _8464 = _8456 ^ _8463;
  wire _8465 = r948 ^ r1048;
  wire _8466 = r1066 ^ r1149;
  wire _8467 = _8465 ^ _8466;
  wire _8468 = r1269 ^ r1279;
  wire _8469 = r1362 ^ r1516;
  wire _8470 = _8468 ^ _8469;
  wire _8471 = _8467 ^ _8470;
  wire _8472 = r1531 ^ r1561;
  wire _8473 = r1607 ^ r1693;
  wire _8474 = _8472 ^ _8473;
  wire _8475 = r1753 ^ r1802;
  wire _8476 = r1806 ^ r1863;
  wire _8477 = _8475 ^ _8476;
  wire _8478 = _8474 ^ _8477;
  wire _8479 = _8471 ^ _8478;
  wire _8480 = _8464 ^ _8479;
  wire _8481 = r44 ^ r133;
  wire _8482 = r203 ^ r244;
  wire _8483 = _8481 ^ _8482;
  wire _8484 = r386 ^ r405;
  wire _8485 = r504 ^ r627;
  wire _8486 = _8484 ^ _8485;
  wire _8487 = _8483 ^ _8486;
  wire _8488 = r759 ^ r855;
  wire _8489 = r918 ^ r945;
  wire _8490 = _8488 ^ _8489;
  wire _8491 = r1023 ^ r1209;
  wire _8492 = r1355 ^ r1385;
  wire _8493 = _8491 ^ _8492;
  wire _8494 = _8490 ^ _8493;
  wire _8495 = _8487 ^ _8494;
  wire _8496 = r1445 ^ r1486;
  wire _8497 = r1532 ^ r1612;
  wire _8498 = _8496 ^ _8497;
  wire _8499 = r1757 ^ r1845;
  wire _8500 = r1858 ^ r1888;
  wire _8501 = _8499 ^ _8500;
  wire _8502 = _8498 ^ _8501;
  wire _8503 = r1906 ^ r1915;
  wire _8504 = r1992 ^ r1993;
  wire _8505 = _8503 ^ _8504;
  wire _8506 = r2028 ^ r2032;
  wire _8507 = r2043 ^ r2046;
  wire _8508 = _8506 ^ _8507;
  wire _8509 = _8505 ^ _8508;
  wire _8510 = _8502 ^ _8509;
  wire _8511 = _8495 ^ _8510;
  wire _8512 = _8480 | _8511;
  wire _8513 = r43 ^ r168;
  wire _8514 = r173 ^ r273;
  wire _8515 = _8513 ^ _8514;
  wire _8516 = r300 ^ r535;
  wire _8517 = r605 ^ r647;
  wire _8518 = _8516 ^ _8517;
  wire _8519 = _8515 ^ _8518;
  wire _8520 = r721 ^ r880;
  wire _8521 = r888 ^ r962;
  wire _8522 = _8520 ^ _8521;
  wire _8523 = r1032 ^ r1095;
  wire _8524 = r1118 ^ r1195;
  wire _8525 = _8523 ^ _8524;
  wire _8526 = _8522 ^ _8525;
  wire _8527 = _8519 ^ _8526;
  wire _8528 = r1230 ^ r1429;
  wire _8529 = r1478 ^ r1530;
  wire _8530 = _8528 ^ _8529;
  wire _8531 = r1534 ^ r1539;
  wire _8532 = r1635 ^ r1725;
  wire _8533 = _8531 ^ _8532;
  wire _8534 = _8530 ^ _8533;
  wire _8535 = r1815 ^ r1824;
  wire _8536 = r1827 ^ r1898;
  wire _8537 = _8535 ^ _8536;
  wire _8538 = r1908 ^ r1965;
  wire _8539 = r1996 ^ r2006;
  wire _8540 = _8538 ^ _8539;
  wire _8541 = _8537 ^ _8540;
  wire _8542 = _8534 ^ _8541;
  wire _8543 = _8527 ^ _8542;
  wire _8544 = r42 ^ r72;
  wire _8545 = r159 ^ r180;
  wire _8546 = _8544 ^ _8545;
  wire _8547 = r241 ^ r280;
  wire _8548 = r364 ^ r432;
  wire _8549 = _8547 ^ _8548;
  wire _8550 = _8546 ^ _8549;
  wire _8551 = r490 ^ r549;
  wire _8552 = r562 ^ r654;
  wire _8553 = _8551 ^ _8552;
  wire _8554 = r677 ^ r794;
  wire _8555 = r866 ^ r932;
  wire _8556 = _8554 ^ _8555;
  wire _8557 = _8553 ^ _8556;
  wire _8558 = _8550 ^ _8557;
  wire _8559 = r954 ^ r1026;
  wire _8560 = r1101 ^ r1158;
  wire _8561 = _8559 ^ _8560;
  wire _8562 = r1212 ^ r1272;
  wire _8563 = r1327 ^ r1339;
  wire _8564 = _8562 ^ _8563;
  wire _8565 = _8561 ^ _8564;
  wire _8566 = r1390 ^ r1421;
  wire _8567 = r1601 ^ r1628;
  wire _8568 = _8566 ^ _8567;
  wire _8569 = r1677 ^ r1692;
  wire _8570 = r1724 ^ r1864;
  wire _8571 = _8569 ^ _8570;
  wire _8572 = _8568 ^ _8571;
  wire _8573 = _8565 ^ _8572;
  wire _8574 = _8558 ^ _8573;
  wire _8575 = _8543 | _8574;
  wire _8576 = _8512 | _8575;
  wire _8577 = r41 ^ r109;
  wire _8578 = r118 ^ r216;
  wire _8579 = _8577 ^ _8578;
  wire _8580 = r266 ^ r325;
  wire _8581 = r360 ^ r412;
  wire _8582 = _8580 ^ _8581;
  wire _8583 = _8579 ^ _8582;
  wire _8584 = r464 ^ r559;
  wire _8585 = r570 ^ r652;
  wire _8586 = _8584 ^ _8585;
  wire _8587 = r705 ^ r775;
  wire _8588 = r792 ^ r921;
  wire _8589 = _8587 ^ _8588;
  wire _8590 = _8586 ^ _8589;
  wire _8591 = _8583 ^ _8590;
  wire _8592 = r987 ^ r1029;
  wire _8593 = r1072 ^ r1114;
  wire _8594 = _8592 ^ _8593;
  wire _8595 = r1176 ^ r1233;
  wire _8596 = r1309 ^ r1335;
  wire _8597 = _8595 ^ _8596;
  wire _8598 = _8594 ^ _8597;
  wire _8599 = r1391 ^ r1430;
  wire _8600 = r1449 ^ r1459;
  wire _8601 = _8599 ^ _8600;
  wire _8602 = r1616 ^ r1678;
  wire _8603 = r1711 ^ r1787;
  wire _8604 = _8602 ^ _8603;
  wire _8605 = _8601 ^ _8604;
  wire _8606 = _8598 ^ _8605;
  wire _8607 = _8591 ^ _8606;
  wire _8608 = r67 ^ r122;
  wire _8609 = r218 ^ r250;
  wire _8610 = _8608 ^ _8609;
  wire _8611 = r287 ^ r381;
  wire _8612 = r424 ^ r498;
  wire _8613 = _8611 ^ _8612;
  wire _8614 = _8610 ^ _8613;
  wire _8615 = r529 ^ r599;
  wire _8616 = r655 ^ r693;
  wire _8617 = _8615 ^ _8616;
  wire _8618 = r762 ^ r825;
  wire _8619 = r882 ^ r935;
  wire _8620 = _8618 ^ _8619;
  wire _8621 = _8617 ^ _8620;
  wire _8622 = _8614 ^ _8621;
  wire _8623 = r997 ^ r1070;
  wire _8624 = r1124 ^ r1185;
  wire _8625 = _8623 ^ _8624;
  wire _8626 = r1251 ^ r1315;
  wire _8627 = r1337 ^ r1384;
  wire _8628 = _8626 ^ _8627;
  wire _8629 = _8625 ^ _8628;
  wire _8630 = r1395 ^ r1444;
  wire _8631 = r1580 ^ r1631;
  wire _8632 = _8630 ^ _8631;
  wire _8633 = r1656 ^ r1739;
  wire _8634 = r1810 ^ r1892;
  wire _8635 = _8633 ^ _8634;
  wire _8636 = _8632 ^ _8635;
  wire _8637 = _8629 ^ _8636;
  wire _8638 = _8622 ^ _8637;
  wire _8639 = _8607 | _8638;
  wire _8640 = r40 ^ r79;
  wire _8641 = r170 ^ r190;
  wire _8642 = _8640 ^ _8641;
  wire _8643 = r275 ^ r292;
  wire _8644 = r344 ^ r433;
  wire _8645 = _8643 ^ _8644;
  wire _8646 = _8642 ^ _8645;
  wire _8647 = r466 ^ r518;
  wire _8648 = r612 ^ r646;
  wire _8649 = _8647 ^ _8648;
  wire _8650 = r680 ^ r737;
  wire _8651 = r805 ^ r869;
  wire _8652 = _8650 ^ _8651;
  wire _8653 = _8649 ^ _8652;
  wire _8654 = _8646 ^ _8653;
  wire _8655 = r900 ^ r991;
  wire _8656 = r1057 ^ r1100;
  wire _8657 = _8655 ^ _8656;
  wire _8658 = r1153 ^ r1180;
  wire _8659 = r1259 ^ r1277;
  wire _8660 = _8658 ^ _8659;
  wire _8661 = _8657 ^ _8660;
  wire _8662 = r1383 ^ r1442;
  wire _8663 = r1542 ^ r1579;
  wire _8664 = _8662 ^ _8663;
  wire _8665 = r1609 ^ r1683;
  wire _8666 = r1707 ^ r1788;
  wire _8667 = _8665 ^ _8666;
  wire _8668 = _8664 ^ _8667;
  wire _8669 = _8661 ^ _8668;
  wire _8670 = _8654 ^ _8669;
  wire _8671 = r39 ^ r105;
  wire _8672 = r171 ^ r268;
  wire _8673 = _8671 ^ _8672;
  wire _8674 = r332 ^ r345;
  wire _8675 = r406 ^ r478;
  wire _8676 = _8674 ^ _8675;
  wire _8677 = _8673 ^ _8676;
  wire _8678 = r507 ^ r586;
  wire _8679 = r696 ^ r758;
  wire _8680 = _8678 ^ _8679;
  wire _8681 = r807 ^ r832;
  wire _8682 = r994 ^ r1038;
  wire _8683 = _8681 ^ _8682;
  wire _8684 = _8680 ^ _8683;
  wire _8685 = _8677 ^ _8684;
  wire _8686 = r1083 ^ r1140;
  wire _8687 = r1255 ^ r1330;
  wire _8688 = _8686 ^ _8687;
  wire _8689 = r1363 ^ r1472;
  wire _8690 = r1544 ^ r1606;
  wire _8691 = _8689 ^ _8690;
  wire _8692 = _8688 ^ _8691;
  wire _8693 = r1608 ^ r1803;
  wire _8694 = r1849 ^ r1852;
  wire _8695 = _8693 ^ _8694;
  wire _8696 = r1895 ^ r1911;
  wire _8697 = r1941 ^ r1948;
  wire _8698 = _8696 ^ _8697;
  wire _8699 = _8695 ^ _8698;
  wire _8700 = _8692 ^ _8699;
  wire _8701 = _8685 ^ _8700;
  wire _8702 = _8670 | _8701;
  wire _8703 = _8639 | _8702;
  wire _8704 = _8576 | _8703;
  wire _8705 = _8449 | _8704;
  wire _8706 = r38 ^ r94;
  wire _8707 = r116 ^ r184;
  wire _8708 = _8706 ^ _8707;
  wire _8709 = r254 ^ r291;
  wire _8710 = r380 ^ r420;
  wire _8711 = _8709 ^ _8710;
  wire _8712 = _8708 ^ _8711;
  wire _8713 = r476 ^ r520;
  wire _8714 = r565 ^ r621;
  wire _8715 = _8713 ^ _8714;
  wire _8716 = r715 ^ r729;
  wire _8717 = r795 ^ r863;
  wire _8718 = _8716 ^ _8717;
  wire _8719 = _8715 ^ _8718;
  wire _8720 = _8712 ^ _8719;
  wire _8721 = r905 ^ r984;
  wire _8722 = r1052 ^ r1086;
  wire _8723 = _8721 ^ _8722;
  wire _8724 = r1127 ^ r1175;
  wire _8725 = r1260 ^ r1313;
  wire _8726 = _8724 ^ _8725;
  wire _8727 = _8723 ^ _8726;
  wire _8728 = r1346 ^ r1406;
  wire _8729 = r1433 ^ r1455;
  wire _8730 = _8728 ^ _8729;
  wire _8731 = r1621 ^ r1657;
  wire _8732 = r1706 ^ r1789;
  wire _8733 = _8731 ^ _8732;
  wire _8734 = _8730 ^ _8733;
  wire _8735 = _8727 ^ _8734;
  wire _8736 = _8720 ^ _8735;
  wire _8737 = r37 ^ r81;
  wire _8738 = r156 ^ r272;
  wire _8739 = _8737 ^ _8738;
  wire _8740 = r285 ^ r371;
  wire _8741 = r493 ^ r541;
  wire _8742 = _8740 ^ _8741;
  wire _8743 = _8739 ^ _8742;
  wire _8744 = r659 ^ r670;
  wire _8745 = r769 ^ r826;
  wire _8746 = _8744 ^ _8745;
  wire _8747 = r860 ^ r910;
  wire _8748 = r963 ^ r1007;
  wire _8749 = _8747 ^ _8748;
  wire _8750 = _8746 ^ _8749;
  wire _8751 = _8743 ^ _8750;
  wire _8752 = r1073 ^ r1143;
  wire _8753 = r1198 ^ r1250;
  wire _8754 = _8752 ^ _8753;
  wire _8755 = r1297 ^ r1358;
  wire _8756 = r1453 ^ r1550;
  wire _8757 = _8755 ^ _8756;
  wire _8758 = _8754 ^ _8757;
  wire _8759 = r1726 ^ r1736;
  wire _8760 = r1817 ^ r1910;
  wire _8761 = _8759 ^ _8760;
  wire _8762 = r1918 ^ r1984;
  wire _8763 = r2031 ^ r2042;
  wire _8764 = _8762 ^ _8763;
  wire _8765 = _8761 ^ _8764;
  wire _8766 = _8758 ^ _8765;
  wire _8767 = _8751 ^ _8766;
  wire _8768 = _8736 | _8767;
  wire _8769 = r36 ^ r164;
  wire _8770 = r217 ^ r248;
  wire _8771 = _8769 ^ _8770;
  wire _8772 = r390 ^ r427;
  wire _8773 = r460 ^ r551;
  wire _8774 = _8772 ^ _8773;
  wire _8775 = _8771 ^ _8774;
  wire _8776 = r601 ^ r661;
  wire _8777 = r739 ^ r874;
  wire _8778 = _8776 ^ _8777;
  wire _8779 = r899 ^ r944;
  wire _8780 = r1033 ^ r1204;
  wire _8781 = _8779 ^ _8780;
  wire _8782 = _8778 ^ _8781;
  wire _8783 = _8775 ^ _8782;
  wire _8784 = r1275 ^ r1282;
  wire _8785 = r1300 ^ r1369;
  wire _8786 = _8784 ^ _8785;
  wire _8787 = r1398 ^ r1564;
  wire _8788 = r1581 ^ r1641;
  wire _8789 = _8787 ^ _8788;
  wire _8790 = _8786 ^ _8789;
  wire _8791 = r1650 ^ r1709;
  wire _8792 = r1985 ^ r2002;
  wire _8793 = _8791 ^ _8792;
  wire _8794 = r2017 ^ r2019;
  wire _8795 = r2029 ^ r2033;
  wire _8796 = _8794 ^ _8795;
  wire _8797 = _8793 ^ _8796;
  wire _8798 = _8790 ^ _8797;
  wire _8799 = _8783 ^ _8798;
  wire _8800 = r35 ^ r59;
  wire _8801 = r128 ^ r179;
  wire _8802 = _8800 ^ _8801;
  wire _8803 = r329 ^ r394;
  wire _8804 = r461 ^ r546;
  wire _8805 = _8803 ^ _8804;
  wire _8806 = _8802 ^ _8805;
  wire _8807 = r597 ^ r817;
  wire _8808 = r923 ^ r958;
  wire _8809 = _8807 ^ _8808;
  wire _8810 = r1022 ^ r1069;
  wire _8811 = r1113 ^ r1115;
  wire _8812 = _8810 ^ _8811;
  wire _8813 = _8809 ^ _8812;
  wire _8814 = _8806 ^ _8813;
  wire _8815 = r1189 ^ r1225;
  wire _8816 = r1286 ^ r1340;
  wire _8817 = _8815 ^ _8816;
  wire _8818 = r1407 ^ r1440;
  wire _8819 = r1458 ^ r1490;
  wire _8820 = _8818 ^ _8819;
  wire _8821 = _8817 ^ _8820;
  wire _8822 = r1668 ^ r1813;
  wire _8823 = r1825 ^ r1848;
  wire _8824 = _8822 ^ _8823;
  wire _8825 = r1851 ^ r1873;
  wire _8826 = r1875 ^ r1893;
  wire _8827 = _8825 ^ _8826;
  wire _8828 = _8824 ^ _8827;
  wire _8829 = _8821 ^ _8828;
  wire _8830 = _8814 ^ _8829;
  wire _8831 = _8799 | _8830;
  wire _8832 = _8768 | _8831;
  wire _8833 = r34 ^ r69;
  wire _8834 = r126 ^ r205;
  wire _8835 = _8833 ^ _8834;
  wire _8836 = r259 ^ r297;
  wire _8837 = r407 ^ r492;
  wire _8838 = _8836 ^ _8837;
  wire _8839 = _8835 ^ _8838;
  wire _8840 = r552 ^ r615;
  wire _8841 = r667 ^ r714;
  wire _8842 = _8840 ^ _8841;
  wire _8843 = r773 ^ r801;
  wire _8844 = r843 ^ r929;
  wire _8845 = _8843 ^ _8844;
  wire _8846 = _8842 ^ _8845;
  wire _8847 = _8839 ^ _8846;
  wire _8848 = r969 ^ r1009;
  wire _8849 = r1093 ^ r1166;
  wire _8850 = _8848 ^ _8849;
  wire _8851 = r1191 ^ r1264;
  wire _8852 = r1314 ^ r1456;
  wire _8853 = _8851 ^ _8852;
  wire _8854 = _8850 ^ _8853;
  wire _8855 = r1496 ^ r1533;
  wire _8856 = r1543 ^ r1578;
  wire _8857 = _8855 ^ _8856;
  wire _8858 = r1644 ^ r1653;
  wire _8859 = r1688 ^ r1790;
  wire _8860 = _8858 ^ _8859;
  wire _8861 = _8857 ^ _8860;
  wire _8862 = _8854 ^ _8861;
  wire _8863 = _8847 ^ _8862;
  wire _8864 = r33 ^ r64;
  wire _8865 = r162 ^ r185;
  wire _8866 = _8864 ^ _8865;
  wire _8867 = r252 ^ r295;
  wire _8868 = r334 ^ r391;
  wire _8869 = _8867 ^ _8868;
  wire _8870 = _8866 ^ _8869;
  wire _8871 = r404 ^ r484;
  wire _8872 = r540 ^ r582;
  wire _8873 = _8871 ^ _8872;
  wire _8874 = r682 ^ r736;
  wire _8875 = r854 ^ r914;
  wire _8876 = _8874 ^ _8875;
  wire _8877 = _8873 ^ _8876;
  wire _8878 = _8870 ^ _8877;
  wire _8879 = r998 ^ r1116;
  wire _8880 = r1266 ^ r1371;
  wire _8881 = _8879 ^ _8880;
  wire _8882 = r1394 ^ r1565;
  wire _8883 = r1599 ^ r1669;
  wire _8884 = _8882 ^ _8883;
  wire _8885 = _8881 ^ _8884;
  wire _8886 = r1751 ^ r1758;
  wire _8887 = r1808 ^ r1936;
  wire _8888 = _8886 ^ _8887;
  wire _8889 = r1951 ^ r2000;
  wire _8890 = r2004 ^ r2010;
  wire _8891 = _8889 ^ _8890;
  wire _8892 = _8888 ^ _8891;
  wire _8893 = _8885 ^ _8892;
  wire _8894 = _8878 ^ _8893;
  wire _8895 = _8863 | _8894;
  wire _8896 = r32 ^ r70;
  wire _8897 = r141 ^ r229;
  wire _8898 = _8896 ^ _8897;
  wire _8899 = r328 ^ r388;
  wire _8900 = r423 ^ r502;
  wire _8901 = _8899 ^ _8900;
  wire _8902 = _8898 ^ _8901;
  wire _8903 = r509 ^ r630;
  wire _8904 = r689 ^ r766;
  wire _8905 = _8903 ^ _8904;
  wire _8906 = r819 ^ r847;
  wire _8907 = r915 ^ r986;
  wire _8908 = _8906 ^ _8907;
  wire _8909 = _8905 ^ _8908;
  wire _8910 = _8902 ^ _8909;
  wire _8911 = r1044 ^ r1102;
  wire _8912 = r1163 ^ r1196;
  wire _8913 = _8911 ^ _8912;
  wire _8914 = r1236 ^ r1306;
  wire _8915 = r1329 ^ r1422;
  wire _8916 = _8914 ^ _8915;
  wire _8917 = _8913 ^ _8916;
  wire _8918 = r1434 ^ r1588;
  wire _8919 = r1638 ^ r1679;
  wire _8920 = _8918 ^ _8919;
  wire _8921 = r1782 ^ r1854;
  wire _8922 = r1934 ^ r1949;
  wire _8923 = _8921 ^ _8922;
  wire _8924 = _8920 ^ _8923;
  wire _8925 = _8917 ^ _8924;
  wire _8926 = _8910 ^ _8925;
  wire _8927 = r31 ^ r58;
  wire _8928 = r144 ^ r219;
  wire _8929 = _8927 ^ _8928;
  wire _8930 = r239 ^ r368;
  wire _8931 = r444 ^ r450;
  wire _8932 = _8930 ^ _8931;
  wire _8933 = _8929 ^ _8932;
  wire _8934 = r614 ^ r660;
  wire _8935 = r851 ^ r939;
  wire _8936 = _8934 ^ _8935;
  wire _8937 = r972 ^ r1054;
  wire _8938 = r1208 ^ r1273;
  wire _8939 = _8937 ^ _8938;
  wire _8940 = _8936 ^ _8939;
  wire _8941 = _8933 ^ _8940;
  wire _8942 = r1294 ^ r1352;
  wire _8943 = r1401 ^ r1452;
  wire _8944 = _8942 ^ _8943;
  wire _8945 = r1460 ^ r1471;
  wire _8946 = r1622 ^ r1676;
  wire _8947 = _8945 ^ _8946;
  wire _8948 = _8944 ^ _8947;
  wire _8949 = r1768 ^ r1779;
  wire _8950 = r1964 ^ r1991;
  wire _8951 = _8949 ^ _8950;
  wire _8952 = r2007 ^ r2011;
  wire _8953 = r2013 ^ r2025;
  wire _8954 = _8952 ^ _8953;
  wire _8955 = _8951 ^ _8954;
  wire _8956 = _8948 ^ _8955;
  wire _8957 = _8941 ^ _8956;
  wire _8958 = _8926 | _8957;
  wire _8959 = _8895 | _8958;
  wire _8960 = _8832 | _8959;
  wire _8961 = r30 ^ r84;
  wire _8962 = r129 ^ r215;
  wire _8963 = _8961 ^ _8962;
  wire _8964 = r233 ^ r310;
  wire _8965 = r376 ^ r445;
  wire _8966 = _8964 ^ _8965;
  wire _8967 = _8963 ^ _8966;
  wire _8968 = r505 ^ r555;
  wire _8969 = r606 ^ r675;
  wire _8970 = _8968 ^ _8969;
  wire _8971 = r723 ^ r824;
  wire _8972 = r840 ^ r989;
  wire _8973 = _8971 ^ _8972;
  wire _8974 = _8970 ^ _8973;
  wire _8975 = _8967 ^ _8974;
  wire _8976 = r1049 ^ r1084;
  wire _8977 = r1136 ^ r1223;
  wire _8978 = _8976 ^ _8977;
  wire _8979 = r1229 ^ r1316;
  wire _8980 = r1360 ^ r1386;
  wire _8981 = _8979 ^ _8980;
  wire _8982 = _8978 ^ _8981;
  wire _8983 = r1424 ^ r1600;
  wire _8984 = r1708 ^ r1740;
  wire _8985 = _8983 ^ _8984;
  wire _8986 = r1777 ^ r1896;
  wire _8987 = r1924 ^ r1927;
  wire _8988 = _8986 ^ _8987;
  wire _8989 = _8985 ^ _8988;
  wire _8990 = _8982 ^ _8989;
  wire _8991 = _8975 ^ _8990;
  wire _8992 = r29 ^ r90;
  wire _8993 = r163 ^ r182;
  wire _8994 = _8992 ^ _8993;
  wire _8995 = r236 ^ r298;
  wire _8996 = r340 ^ r422;
  wire _8997 = _8995 ^ _8996;
  wire _8998 = _8994 ^ _8997;
  wire _8999 = r449 ^ r557;
  wire _9000 = r569 ^ r648;
  wire _9001 = _8999 ^ _9000;
  wire _9002 = r700 ^ r771;
  wire _9003 = r799 ^ r875;
  wire _9004 = _9002 ^ _9003;
  wire _9005 = _9001 ^ _9004;
  wire _9006 = _8998 ^ _9005;
  wire _9007 = r931 ^ r950;
  wire _9008 = r1055 ^ r1060;
  wire _9009 = _9007 ^ _9008;
  wire _9010 = r1099 ^ r1120;
  wire _9011 = r1190 ^ r1237;
  wire _9012 = _9010 ^ _9011;
  wire _9013 = _9009 ^ _9012;
  wire _9014 = r1308 ^ r1356;
  wire _9015 = r1545 ^ r1560;
  wire _9016 = _9014 ^ _9015;
  wire _9017 = r1591 ^ r1617;
  wire _9018 = r1666 ^ r1791;
  wire _9019 = _9017 ^ _9018;
  wire _9020 = _9016 ^ _9019;
  wire _9021 = _9013 ^ _9020;
  wire _9022 = _9006 ^ _9021;
  wire _9023 = _8991 | _9022;
  wire _9024 = r28 ^ r74;
  wire _9025 = r125 ^ r200;
  wire _9026 = _9024 ^ _9025;
  wire _9027 = r226 ^ r338;
  wire _9028 = r413 ^ r500;
  wire _9029 = _9027 ^ _9028;
  wire _9030 = _9026 ^ _9029;
  wire _9031 = r573 ^ r626;
  wire _9032 = r746 ^ r859;
  wire _9033 = _9031 ^ _9032;
  wire _9034 = r940 ^ r960;
  wire _9035 = r1043 ^ r1203;
  wire _9036 = _9034 ^ _9035;
  wire _9037 = _9033 ^ _9036;
  wire _9038 = _9030 ^ _9037;
  wire _9039 = r1265 ^ r1298;
  wire _9040 = r1331 ^ r1361;
  wire _9041 = _9039 ^ _9040;
  wire _9042 = r1388 ^ r1541;
  wire _9043 = r1605 ^ r1627;
  wire _9044 = _9042 ^ _9043;
  wire _9045 = _9041 ^ _9044;
  wire _9046 = r1766 ^ r1785;
  wire _9047 = r1974 ^ r2003;
  wire _9048 = _9046 ^ _9047;
  wire _9049 = r2009 ^ r2040;
  wire _9050 = r2041 ^ r2047;
  wire _9051 = _9049 ^ _9050;
  wire _9052 = _9048 ^ _9051;
  wire _9053 = _9045 ^ _9052;
  wire _9054 = _9038 ^ _9053;
  wire _9055 = r27 ^ r76;
  wire _9056 = r153 ^ r201;
  wire _9057 = _9055 ^ _9056;
  wire _9058 = r260 ^ r294;
  wire _9059 = r374 ^ r431;
  wire _9060 = _9058 ^ _9059;
  wire _9061 = _9057 ^ _9060;
  wire _9062 = r482 ^ r616;
  wire _9063 = r650 ^ r692;
  wire _9064 = _9062 ^ _9063;
  wire _9065 = r756 ^ r810;
  wire _9066 = r870 ^ r955;
  wire _9067 = _9065 ^ _9066;
  wire _9068 = _9064 ^ _9067;
  wire _9069 = _9061 ^ _9068;
  wire _9070 = r1012 ^ r1075;
  wire _9071 = r1147 ^ r1276;
  wire _9072 = _9070 ^ _9071;
  wire _9073 = r1351 ^ r1396;
  wire _9074 = r1435 ^ r1491;
  wire _9075 = _9073 ^ _9074;
  wire _9076 = _9072 ^ _9075;
  wire _9077 = r1524 ^ r1585;
  wire _9078 = r1697 ^ r1829;
  wire _9079 = _9077 ^ _9078;
  wire _9080 = r1835 ^ r1900;
  wire _9081 = r1947 ^ r1955;
  wire _9082 = _9080 ^ _9081;
  wire _9083 = _9079 ^ _9082;
  wire _9084 = _9076 ^ _9083;
  wire _9085 = _9069 ^ _9084;
  wire _9086 = _9054 | _9085;
  wire _9087 = _9023 | _9086;
  wire _9088 = r26 ^ r100;
  wire _9089 = r137 ^ r181;
  wire _9090 = _9088 ^ _9089;
  wire _9091 = r245 ^ r320;
  wire _9092 = r353 ^ r436;
  wire _9093 = _9091 ^ _9092;
  wire _9094 = _9090 ^ _9093;
  wire _9095 = r488 ^ r517;
  wire _9096 = r572 ^ r662;
  wire _9097 = _9095 ^ _9096;
  wire _9098 = r701 ^ r749;
  wire _9099 = r803 ^ r881;
  wire _9100 = _9098 ^ _9099;
  wire _9101 = _9097 ^ _9100;
  wire _9102 = _9094 ^ _9101;
  wire _9103 = r928 ^ r961;
  wire _9104 = r1018 ^ r1088;
  wire _9105 = _9103 ^ _9104;
  wire _9106 = r1128 ^ r1164;
  wire _9107 = r1211 ^ r1252;
  wire _9108 = _9106 ^ _9107;
  wire _9109 = _9105 ^ _9108;
  wire _9110 = r1291 ^ r1374;
  wire _9111 = r1418 ^ r1432;
  wire _9112 = _9110 ^ _9111;
  wire _9113 = r1583 ^ r1640;
  wire _9114 = r1684 ^ r1792;
  wire _9115 = _9113 ^ _9114;
  wire _9116 = _9112 ^ _9115;
  wire _9117 = _9109 ^ _9116;
  wire _9118 = _9102 ^ _9117;
  wire _9119 = r25 ^ r82;
  wire _9120 = r165 ^ r172;
  wire _9121 = _9119 ^ _9120;
  wire _9122 = r255 ^ r304;
  wire _9123 = r355 ^ r447;
  wire _9124 = _9122 ^ _9123;
  wire _9125 = _9121 ^ _9124;
  wire _9126 = r456 ^ r524;
  wire _9127 = r567 ^ r658;
  wire _9128 = _9126 ^ _9127;
  wire _9129 = r674 ^ r753;
  wire _9130 = r780 ^ r901;
  wire _9131 = _9129 ^ _9130;
  wire _9132 = _9128 ^ _9131;
  wire _9133 = _9125 ^ _9132;
  wire _9134 = r949 ^ r1081;
  wire _9135 = r1139 ^ r1178;
  wire _9136 = _9134 ^ _9135;
  wire _9137 = r1232 ^ r1281;
  wire _9138 = r1288 ^ r1380;
  wire _9139 = _9137 ^ _9138;
  wire _9140 = _9136 ^ _9139;
  wire _9141 = r1419 ^ r1474;
  wire _9142 = r1504 ^ r1593;
  wire _9143 = _9141 ^ _9142;
  wire _9144 = r1701 ^ r1731;
  wire _9145 = r1755 ^ r1865;
  wire _9146 = _9144 ^ _9145;
  wire _9147 = _9143 ^ _9146;
  wire _9148 = _9140 ^ _9147;
  wire _9149 = _9133 ^ _9148;
  wire _9150 = _9118 | _9149;
  wire _9151 = r24 ^ r93;
  wire _9152 = r155 ^ r189;
  wire _9153 = _9151 ^ _9152;
  wire _9154 = r267 ^ r330;
  wire _9155 = r341 ^ r435;
  wire _9156 = _9154 ^ _9155;
  wire _9157 = _9153 ^ _9156;
  wire _9158 = r454 ^ r556;
  wire _9159 = r603 ^ r623;
  wire _9160 = _9158 ^ _9159;
  wire _9161 = r688 ^ r744;
  wire _9162 = r790 ^ r842;
  wire _9163 = _9161 ^ _9162;
  wire _9164 = _9160 ^ _9163;
  wire _9165 = _9157 ^ _9164;
  wire _9166 = r887 ^ r934;
  wire _9167 = r975 ^ r1005;
  wire _9168 = _9166 ^ _9167;
  wire _9169 = r1148 ^ r1192;
  wire _9170 = r1254 ^ r1333;
  wire _9171 = _9169 ^ _9170;
  wire _9172 = _9168 ^ _9171;
  wire _9173 = r1364 ^ r1507;
  wire _9174 = r1589 ^ r1643;
  wire _9175 = _9173 ^ _9174;
  wire _9176 = r1659 ^ r1752;
  wire _9177 = r1764 ^ r1866;
  wire _9178 = _9176 ^ _9177;
  wire _9179 = _9175 ^ _9178;
  wire _9180 = _9172 ^ _9179;
  wire _9181 = _9165 ^ _9180;
  wire _9182 = r23 ^ r101;
  wire _9183 = r142 ^ r193;
  wire _9184 = _9182 ^ _9183;
  wire _9185 = r240 ^ r322;
  wire _9186 = r375 ^ r429;
  wire _9187 = _9185 ^ _9186;
  wire _9188 = _9184 ^ _9187;
  wire _9189 = r486 ^ r514;
  wire _9190 = r610 ^ r643;
  wire _9191 = _9189 ^ _9190;
  wire _9192 = r716 ^ r722;
  wire _9193 = r724 ^ r784;
  wire _9194 = _9192 ^ _9193;
  wire _9195 = _9191 ^ _9194;
  wire _9196 = _9188 ^ _9195;
  wire _9197 = r884 ^ r903;
  wire _9198 = r981 ^ r1028;
  wire _9199 = _9197 ^ _9198;
  wire _9200 = r1068 ^ r1121;
  wire _9201 = r1188 ^ r1267;
  wire _9202 = _9200 ^ _9201;
  wire _9203 = _9199 ^ _9202;
  wire _9204 = r1296 ^ r1334;
  wire _9205 = r1366 ^ r1476;
  wire _9206 = _9204 ^ _9205;
  wire _9207 = r1551 ^ r1611;
  wire _9208 = r1687 ^ r1793;
  wire _9209 = _9207 ^ _9208;
  wire _9210 = _9206 ^ _9209;
  wire _9211 = _9203 ^ _9210;
  wire _9212 = _9196 ^ _9211;
  wire _9213 = _9181 | _9212;
  wire _9214 = _9150 | _9213;
  wire _9215 = _9087 | _9214;
  wire _9216 = _8960 | _9215;
  wire _9217 = _8705 | _9216;
  wire _9218 = r22 ^ r75;
  wire _9219 = r161 ^ r224;
  wire _9220 = _9218 ^ _9219;
  wire _9221 = r228 ^ r308;
  wire _9222 = r337 ^ r410;
  wire _9223 = _9221 ^ _9222;
  wire _9224 = _9220 ^ _9223;
  wire _9225 = r468 ^ r542;
  wire _9226 = r578 ^ r644;
  wire _9227 = _9225 ^ _9226;
  wire _9228 = r695 ^ r763;
  wire _9229 = r787 ^ r845;
  wire _9230 = _9228 ^ _9229;
  wire _9231 = _9227 ^ _9230;
  wire _9232 = _9224 ^ _9231;
  wire _9233 = r916 ^ r964;
  wire _9234 = r1010 ^ r1061;
  wire _9235 = _9233 ^ _9234;
  wire _9236 = r1135 ^ r1168;
  wire _9237 = r1206 ^ r1263;
  wire _9238 = _9236 ^ _9237;
  wire _9239 = _9235 ^ _9238;
  wire _9240 = r1324 ^ r1405;
  wire _9241 = r1473 ^ r1487;
  wire _9242 = _9240 ^ _9241;
  wire _9243 = r1619 ^ r1658;
  wire _9244 = r1713 ^ r1794;
  wire _9245 = _9243 ^ _9244;
  wire _9246 = _9242 ^ _9245;
  wire _9247 = _9239 ^ _9246;
  wire _9248 = _9232 ^ _9247;
  wire _9249 = r21 ^ r89;
  wire _9250 = r134 ^ r192;
  wire _9251 = _9249 ^ _9250;
  wire _9252 = r269 ^ r327;
  wire _9253 = r365 ^ r418;
  wire _9254 = _9252 ^ _9253;
  wire _9255 = _9251 ^ _9254;
  wire _9256 = r471 ^ r519;
  wire _9257 = r577 ^ r622;
  wire _9258 = _9256 ^ _9257;
  wire _9259 = r717 ^ r774;
  wire _9260 = r778 ^ r913;
  wire _9261 = _9259 ^ _9260;
  wire _9262 = _9258 ^ _9261;
  wire _9263 = _9255 ^ _9262;
  wire _9264 = r966 ^ r1021;
  wire _9265 = r1065 ^ r1110;
  wire _9266 = _9264 ^ _9265;
  wire _9267 = r1173 ^ r1227;
  wire _9268 = r1283 ^ r1372;
  wire _9269 = _9267 ^ _9268;
  wire _9270 = _9266 ^ _9269;
  wire _9271 = r1410 ^ r1441;
  wire _9272 = r1479 ^ r1510;
  wire _9273 = _9271 ^ _9272;
  wire _9274 = r1614 ^ r1654;
  wire _9275 = r1994 ^ r1998;
  wire _9276 = _9274 ^ _9275;
  wire _9277 = _9273 ^ _9276;
  wire _9278 = _9270 ^ _9277;
  wire _9279 = _9263 ^ _9278;
  wire _9280 = _9248 | _9279;
  wire _9281 = r20 ^ r60;
  wire _9282 = r131 ^ r187;
  wire _9283 = _9281 ^ _9282;
  wire _9284 = r231 ^ r350;
  wire _9285 = r440 ^ r457;
  wire _9286 = _9284 ^ _9285;
  wire _9287 = _9283 ^ _9286;
  wire _9288 = r544 ^ r608;
  wire _9289 = r676 ^ r730;
  wire _9290 = _9288 ^ _9289;
  wire _9291 = r811 ^ r872;
  wire _9292 = r992 ^ r1107;
  wire _9293 = _9291 ^ _9292;
  wire _9294 = _9290 ^ _9293;
  wire _9295 = _9287 ^ _9294;
  wire _9296 = r1142 ^ r1174;
  wire _9297 = r1247 ^ r1328;
  wire _9298 = _9296 ^ _9297;
  wire _9299 = r1483 ^ r1552;
  wire _9300 = r1558 ^ r1563;
  wire _9301 = _9299 ^ _9300;
  wire _9302 = _9298 ^ _9301;
  wire _9303 = r1620 ^ r1712;
  wire _9304 = r1783 ^ r1820;
  wire _9305 = _9303 ^ _9304;
  wire _9306 = r1850 ^ r1886;
  wire _9307 = r1972 ^ r1977;
  wire _9308 = _9306 ^ _9307;
  wire _9309 = _9305 ^ _9308;
  wire _9310 = _9302 ^ _9309;
  wire _9311 = _9295 ^ _9310;
  wire _9312 = r19 ^ r96;
  wire _9313 = r147 ^ r223;
  wire _9314 = _9312 ^ _9313;
  wire _9315 = r249 ^ r377;
  wire _9316 = r439 ^ r487;
  wire _9317 = _9315 ^ _9316;
  wire _9318 = _9314 ^ _9317;
  wire _9319 = r558 ^ r590;
  wire _9320 = r629 ^ r673;
  wire _9321 = _9319 ^ _9320;
  wire _9322 = r757 ^ r796;
  wire _9323 = r867 ^ r896;
  wire _9324 = _9322 ^ _9323;
  wire _9325 = _9321 ^ _9324;
  wire _9326 = _9318 ^ _9325;
  wire _9327 = r973 ^ r1004;
  wire _9328 = r1089 ^ r1205;
  wire _9329 = _9327 ^ _9328;
  wire _9330 = r1248 ^ r1336;
  wire _9331 = r1409 ^ r1450;
  wire _9332 = _9330 ^ _9331;
  wire _9333 = _9329 ^ _9332;
  wire _9334 = r1465 ^ r1494;
  wire _9335 = r1512 ^ r1529;
  wire _9336 = _9334 ^ _9335;
  wire _9337 = r1568 ^ r1610;
  wire _9338 = r1767 ^ r1867;
  wire _9339 = _9337 ^ _9338;
  wire _9340 = _9336 ^ _9339;
  wire _9341 = _9333 ^ _9340;
  wire _9342 = _9326 ^ _9341;
  wire _9343 = _9311 | _9342;
  wire _9344 = _9280 | _9343;
  wire _9345 = r18 ^ r62;
  wire _9346 = r139 ^ r177;
  wire _9347 = _9345 ^ _9346;
  wire _9348 = r257 ^ r313;
  wire _9349 = r367 ^ r416;
  wire _9350 = _9348 ^ _9349;
  wire _9351 = _9347 ^ _9350;
  wire _9352 = r453 ^ r554;
  wire _9353 = r592 ^ r633;
  wire _9354 = _9352 ^ _9353;
  wire _9355 = r690 ^ r745;
  wire _9356 = r806 ^ r873;
  wire _9357 = _9355 ^ _9356;
  wire _9358 = _9354 ^ _9357;
  wire _9359 = _9351 ^ _9358;
  wire _9360 = r897 ^ r985;
  wire _9361 = r1017 ^ r1074;
  wire _9362 = _9360 ^ _9361;
  wire _9363 = r1122 ^ r1197;
  wire _9364 = r1226 ^ r1321;
  wire _9365 = _9363 ^ _9364;
  wire _9366 = _9362 ^ _9365;
  wire _9367 = r1365 ^ r1403;
  wire _9368 = r1575 ^ r1594;
  wire _9369 = _9367 ^ _9368;
  wire _9370 = r1630 ^ r1663;
  wire _9371 = r1705 ^ r1795;
  wire _9372 = _9370 ^ _9371;
  wire _9373 = _9369 ^ _9372;
  wire _9374 = _9366 ^ _9373;
  wire _9375 = _9359 ^ _9374;
  wire _9376 = r17 ^ r77;
  wire _9377 = r113 ^ r197;
  wire _9378 = _9376 ^ _9377;
  wire _9379 = r306 ^ r354;
  wire _9380 = r397 ^ r479;
  wire _9381 = _9379 ^ _9380;
  wire _9382 = _9378 ^ _9381;
  wire _9383 = r516 ^ r579;
  wire _9384 = r668 ^ r712;
  wire _9385 = _9383 ^ _9384;
  wire _9386 = r732 ^ r818;
  wire _9387 = r864 ^ r930;
  wire _9388 = _9386 ^ _9387;
  wire _9389 = _9385 ^ _9388;
  wire _9390 = _9382 ^ _9389;
  wire _9391 = r993 ^ r1045;
  wire _9392 = r1085 ^ r1119;
  wire _9393 = _9391 ^ _9392;
  wire _9394 = r1214 ^ r1274;
  wire _9395 = r1302 ^ r1379;
  wire _9396 = _9394 ^ _9395;
  wire _9397 = _9393 ^ _9396;
  wire _9398 = r1448 ^ r1548;
  wire _9399 = r1567 ^ r1582;
  wire _9400 = _9398 ^ _9399;
  wire _9401 = r1636 ^ r1662;
  wire _9402 = r1696 ^ r1796;
  wire _9403 = _9401 ^ _9402;
  wire _9404 = _9400 ^ _9403;
  wire _9405 = _9397 ^ _9404;
  wire _9406 = _9390 ^ _9405;
  wire _9407 = _9375 | _9406;
  wire _9408 = r16 ^ r73;
  wire _9409 = r123 ^ r196;
  wire _9410 = _9408 ^ _9409;
  wire _9411 = r258 ^ r284;
  wire _9412 = r373 ^ r400;
  wire _9413 = _9411 ^ _9412;
  wire _9414 = _9410 ^ _9413;
  wire _9415 = r465 ^ r537;
  wire _9416 = r609 ^ r632;
  wire _9417 = _9415 ^ _9416;
  wire _9418 = r713 ^ r748;
  wire _9419 = r791 ^ r831;
  wire _9420 = _9418 ^ _9419;
  wire _9421 = _9417 ^ _9420;
  wire _9422 = _9414 ^ _9421;
  wire _9423 = r922 ^ r965;
  wire _9424 = r1024 ^ r1094;
  wire _9425 = _9423 ^ _9424;
  wire _9426 = r1138 ^ r1217;
  wire _9427 = r1235 ^ r1287;
  wire _9428 = _9426 ^ _9427;
  wire _9429 = _9425 ^ _9428;
  wire _9430 = r1353 ^ r1393;
  wire _9431 = r1555 ^ r1562;
  wire _9432 = _9430 ^ _9431;
  wire _9433 = r1624 ^ r1686;
  wire _9434 = r1689 ^ r1797;
  wire _9435 = _9433 ^ _9434;
  wire _9436 = _9432 ^ _9435;
  wire _9437 = _9429 ^ _9436;
  wire _9438 = _9422 ^ _9437;
  wire _9439 = r15 ^ r92;
  wire _9440 = r117 ^ r175;
  wire _9441 = _9439 ^ _9440;
  wire _9442 = r346 ^ r441;
  wire _9443 = r489 ^ r538;
  wire _9444 = _9442 ^ _9443;
  wire _9445 = _9441 ^ _9444;
  wire _9446 = r576 ^ r628;
  wire _9447 = r768 ^ r837;
  wire _9448 = _9446 ^ _9447;
  wire _9449 = r938 ^ r1047;
  wire _9450 = r1160 ^ r1169;
  wire _9451 = _9449 ^ _9450;
  wire _9452 = _9448 ^ _9451;
  wire _9453 = _9445 ^ _9452;
  wire _9454 = r1299 ^ r1415;
  wire _9455 = r1439 ^ r1519;
  wire _9456 = _9454 ^ _9455;
  wire _9457 = r1535 ^ r1670;
  wire _9458 = r1699 ^ r1737;
  wire _9459 = _9457 ^ _9458;
  wire _9460 = _9456 ^ _9459;
  wire _9461 = r1756 ^ r1826;
  wire _9462 = r1843 ^ r1931;
  wire _9463 = _9461 ^ _9462;
  wire _9464 = r1975 ^ r1982;
  wire _9465 = r1987 ^ r1989;
  wire _9466 = _9464 ^ _9465;
  wire _9467 = _9463 ^ _9466;
  wire _9468 = _9460 ^ _9467;
  wire _9469 = _9453 ^ _9468;
  wire _9470 = _9438 | _9469;
  wire _9471 = _9407 | _9470;
  wire _9472 = _9344 | _9471;
  wire _9473 = r14 ^ r55;
  wire _9474 = r121 ^ r208;
  wire _9475 = _9473 ^ _9474;
  wire _9476 = r286 ^ r343;
  wire _9477 = r417 ^ r481;
  wire _9478 = _9476 ^ _9477;
  wire _9479 = _9475 ^ _9478;
  wire _9480 = r515 ^ r665;
  wire _9481 = r681 ^ r820;
  wire _9482 = _9480 ^ _9481;
  wire _9483 = r951 ^ r1109;
  wire _9484 = r1161 ^ r1216;
  wire _9485 = _9483 ^ _9484;
  wire _9486 = _9482 ^ _9485;
  wire _9487 = _9479 ^ _9486;
  wire _9488 = r1307 ^ r1413;
  wire _9489 = r1469 ^ r1525;
  wire _9490 = _9488 ^ _9489;
  wire _9491 = r1577 ^ r1646;
  wire _9492 = r1671 ^ r1832;
  wire _9493 = _9491 ^ _9492;
  wire _9494 = _9490 ^ _9493;
  wire _9495 = r1838 ^ r1880;
  wire _9496 = r1882 ^ r1897;
  wire _9497 = _9495 ^ _9496;
  wire _9498 = r1902 ^ r1933;
  wire _9499 = r1950 ^ r1956;
  wire _9500 = _9498 ^ _9499;
  wire _9501 = _9497 ^ _9500;
  wire _9502 = _9494 ^ _9501;
  wire _9503 = _9487 ^ _9502;
  wire _9504 = r13 ^ r56;
  wire _9505 = r111 ^ r211;
  wire _9506 = _9504 ^ _9505;
  wire _9507 = r277 ^ r290;
  wire _9508 = r358 ^ r438;
  wire _9509 = _9507 ^ _9508;
  wire _9510 = _9506 ^ _9509;
  wire _9511 = r469 ^ r508;
  wire _9512 = r587 ^ r620;
  wire _9513 = _9511 ^ _9512;
  wire _9514 = r699 ^ r772;
  wire _9515 = r782 ^ r878;
  wire _9516 = _9514 ^ _9515;
  wire _9517 = _9513 ^ _9516;
  wire _9518 = _9510 ^ _9517;
  wire _9519 = r988 ^ r1058;
  wire _9520 = r1096 ^ r1137;
  wire _9521 = _9519 ^ _9520;
  wire _9522 = r1165 ^ r1239;
  wire _9523 = r1284 ^ r1367;
  wire _9524 = _9522 ^ _9523;
  wire _9525 = _9521 ^ _9524;
  wire _9526 = r1502 ^ r1629;
  wire _9527 = r1734 ^ r1744;
  wire _9528 = _9526 ^ _9527;
  wire _9529 = r1763 ^ r1781;
  wire _9530 = r1784 ^ r1868;
  wire _9531 = _9529 ^ _9530;
  wire _9532 = _9528 ^ _9531;
  wire _9533 = _9525 ^ _9532;
  wire _9534 = _9518 ^ _9533;
  wire _9535 = _9503 | _9534;
  wire _9536 = r12 ^ r91;
  wire _9537 = r148 ^ r198;
  wire _9538 = _9536 ^ _9537;
  wire _9539 = r262 ^ r282;
  wire _9540 = r351 ^ r408;
  wire _9541 = _9539 ^ _9540;
  wire _9542 = _9538 ^ _9541;
  wire _9543 = r485 ^ r523;
  wire _9544 = r611 ^ r639;
  wire _9545 = _9543 ^ _9544;
  wire _9546 = r704 ^ r776;
  wire _9547 = r800 ^ r849;
  wire _9548 = _9546 ^ _9547;
  wire _9549 = _9545 ^ _9548;
  wire _9550 = _9542 ^ _9549;
  wire _9551 = r942 ^ r953;
  wire _9552 = r1020 ^ r1129;
  wire _9553 = _9551 ^ _9552;
  wire _9554 = r1194 ^ r1224;
  wire _9555 = r1234 ^ r1323;
  wire _9556 = _9554 ^ _9555;
  wire _9557 = _9553 ^ _9556;
  wire _9558 = r1495 ^ r1508;
  wire _9559 = r1572 ^ r1602;
  wire _9560 = _9558 ^ _9559;
  wire _9561 = r1639 ^ r1772;
  wire _9562 = r1776 ^ r1869;
  wire _9563 = _9561 ^ _9562;
  wire _9564 = _9560 ^ _9563;
  wire _9565 = _9557 ^ _9564;
  wire _9566 = _9550 ^ _9565;
  wire _9567 = r83 ^ r130;
  wire _9568 = r176 ^ r264;
  wire _9569 = _9567 ^ _9568;
  wire _9570 = r314 ^ r385;
  wire _9571 = r393 ^ r462;
  wire _9572 = _9570 ^ _9571;
  wire _9573 = _9569 ^ _9572;
  wire _9574 = r527 ^ r637;
  wire _9575 = r767 ^ r808;
  wire _9576 = _9574 ^ _9575;
  wire _9577 = r885 ^ r936;
  wire _9578 = r967 ^ r1040;
  wire _9579 = _9577 ^ _9578;
  wire _9580 = _9576 ^ _9579;
  wire _9581 = _9573 ^ _9580;
  wire _9582 = r1079 ^ r1146;
  wire _9583 = r1201 ^ r1271;
  wire _9584 = _9582 ^ _9583;
  wire _9585 = r1382 ^ r1451;
  wire _9586 = r1467 ^ r1477;
  wire _9587 = _9585 ^ _9586;
  wire _9588 = _9584 ^ _9587;
  wire _9589 = r1498 ^ r1538;
  wire _9590 = r1647 ^ r1733;
  wire _9591 = _9589 ^ _9590;
  wire _9592 = r1746 ^ r1883;
  wire _9593 = r1889 ^ r1912;
  wire _9594 = _9592 ^ _9593;
  wire _9595 = _9591 ^ _9594;
  wire _9596 = _9588 ^ _9595;
  wire _9597 = _9581 ^ _9596;
  wire _9598 = _9566 | _9597;
  wire _9599 = _9535 | _9598;
  wire _9600 = r11 ^ r99;
  wire _9601 = r143 ^ r195;
  wire _9602 = _9600 ^ _9601;
  wire _9603 = r299 ^ r335;
  wire _9604 = r419 ^ r459;
  wire _9605 = _9603 ^ _9604;
  wire _9606 = _9602 ^ _9605;
  wire _9607 = r591 ^ r618;
  wire _9608 = r703 ^ r735;
  wire _9609 = _9607 ^ _9608;
  wire _9610 = r804 ^ r841;
  wire _9611 = r920 ^ r1041;
  wire _9612 = _9610 ^ _9611;
  wire _9613 = _9609 ^ _9612;
  wire _9614 = _9606 ^ _9613;
  wire _9615 = r1087 ^ r1151;
  wire _9616 = r1326 ^ r1348;
  wire _9617 = _9615 ^ _9616;
  wire _9618 = r1426 ^ r1497;
  wire _9619 = r1518 ^ r1522;
  wire _9620 = _9618 ^ _9619;
  wire _9621 = _9617 ^ _9620;
  wire _9622 = r1557 ^ r1587;
  wire _9623 = r1625 ^ r1680;
  wire _9624 = _9622 ^ _9623;
  wire _9625 = r1774 ^ r1831;
  wire _9626 = r1859 ^ r1894;
  wire _9627 = _9625 ^ _9626;
  wire _9628 = _9624 ^ _9627;
  wire _9629 = _9621 ^ _9628;
  wire _9630 = _9614 ^ _9629;
  wire _9631 = r10 ^ r103;
  wire _9632 = r154 ^ r220;
  wire _9633 = _9631 ^ _9632;
  wire _9634 = r270 ^ r309;
  wire _9635 = r389 ^ r409;
  wire _9636 = _9634 ^ _9635;
  wire _9637 = _9633 ^ _9636;
  wire _9638 = r474 ^ r526;
  wire _9639 = r697 ^ r741;
  wire _9640 = _9638 ^ _9639;
  wire _9641 = r809 ^ r850;
  wire _9642 = r983 ^ r1019;
  wire _9643 = _9641 ^ _9642;
  wire _9644 = _9640 ^ _9643;
  wire _9645 = _9637 ^ _9644;
  wire _9646 = r1082 ^ r1243;
  wire _9647 = r1349 ^ r1428;
  wire _9648 = _9646 ^ _9647;
  wire _9649 = r1514 ^ r1553;
  wire _9650 = r1691 ^ r1773;
  wire _9651 = _9649 ^ _9650;
  wire _9652 = _9648 ^ _9651;
  wire _9653 = r1812 ^ r1847;
  wire _9654 = r1855 ^ r1856;
  wire _9655 = _9653 ^ _9654;
  wire _9656 = r1903 ^ r1904;
  wire _9657 = r1916 ^ r1920;
  wire _9658 = _9656 ^ _9657;
  wire _9659 = _9655 ^ _9658;
  wire _9660 = _9652 ^ _9659;
  wire _9661 = _9645 ^ _9660;
  wire _9662 = _9630 | _9661;
  wire _9663 = r9 ^ r110;
  wire _9664 = r124 ^ r206;
  wire _9665 = _9663 ^ _9664;
  wire _9666 = r227 ^ r321;
  wire _9667 = r398 ^ r521;
  wire _9668 = _9666 ^ _9667;
  wire _9669 = _9665 ^ _9668;
  wire _9670 = r583 ^ r679;
  wire _9671 = r725 ^ r877;
  wire _9672 = _9670 ^ _9671;
  wire _9673 = r892 ^ r946;
  wire _9674 = r1011 ^ r1150;
  wire _9675 = _9673 ^ _9674;
  wire _9676 = _9672 ^ _9675;
  wire _9677 = _9669 ^ _9676;
  wire _9678 = r1199 ^ r1381;
  wire _9679 = r1412 ^ r1443;
  wire _9680 = _9678 ^ _9679;
  wire _9681 = r1573 ^ r1590;
  wire _9682 = r1649 ^ r1759;
  wire _9683 = _9681 ^ _9682;
  wire _9684 = _9680 ^ _9683;
  wire _9685 = r1769 ^ r1816;
  wire _9686 = r1818 ^ r1821;
  wire _9687 = _9685 ^ _9686;
  wire _9688 = r1823 ^ r1885;
  wire _9689 = r1914 ^ r1917;
  wire _9690 = _9688 ^ _9689;
  wire _9691 = _9687 ^ _9690;
  wire _9692 = _9684 ^ _9691;
  wire _9693 = _9677 ^ _9692;
  wire _9694 = r8 ^ r102;
  wire _9695 = r112 ^ r178;
  wire _9696 = _9694 ^ _9695;
  wire _9697 = r235 ^ r293;
  wire _9698 = r382 ^ r415;
  wire _9699 = _9697 ^ _9698;
  wire _9700 = _9696 ^ _9699;
  wire _9701 = r497 ^ r506;
  wire _9702 = r581 ^ r640;
  wire _9703 = _9701 ^ _9702;
  wire _9704 = r686 ^ r727;
  wire _9705 = r823 ^ r836;
  wire _9706 = _9704 ^ _9705;
  wire _9707 = _9703 ^ _9706;
  wire _9708 = _9700 ^ _9707;
  wire _9709 = r890 ^ r947;
  wire _9710 = r1003 ^ r1027;
  wire _9711 = _9709 ^ _9710;
  wire _9712 = r1078 ^ r1144;
  wire _9713 = r1181 ^ r1373;
  wire _9714 = _9712 ^ _9713;
  wire _9715 = _9711 ^ _9714;
  wire _9716 = r1468 ^ r1520;
  wire _9717 = r1546 ^ r1592;
  wire _9718 = _9716 ^ _9717;
  wire _9719 = r1642 ^ r1681;
  wire _9720 = r1762 ^ r1870;
  wire _9721 = _9719 ^ _9720;
  wire _9722 = _9718 ^ _9721;
  wire _9723 = _9715 ^ _9722;
  wire _9724 = _9708 ^ _9723;
  wire _9725 = _9693 | _9724;
  wire _9726 = _9662 | _9725;
  wire _9727 = _9599 | _9726;
  wire _9728 = _9472 | _9727;
  wire _9729 = r7 ^ r97;
  wire _9730 = r157 ^ r222;
  wire _9731 = _9729 ^ _9730;
  wire _9732 = r263 ^ r283;
  wire _9733 = r359 ^ r446;
  wire _9734 = _9732 ^ _9733;
  wire _9735 = _9731 ^ _9734;
  wire _9736 = r451 ^ r512;
  wire _9737 = r595 ^ r619;
  wire _9738 = _9736 ^ _9737;
  wire _9739 = r709 ^ r751;
  wire _9740 = r828 ^ r865;
  wire _9741 = _9739 ^ _9740;
  wire _9742 = _9738 ^ _9741;
  wire _9743 = _9735 ^ _9742;
  wire _9744 = r925 ^ r982;
  wire _9745 = r1031 ^ r1098;
  wire _9746 = _9744 ^ _9745;
  wire _9747 = r1126 ^ r1167;
  wire _9748 = r1184 ^ r1256;
  wire _9749 = _9747 ^ _9748;
  wire _9750 = _9746 ^ _9749;
  wire _9751 = r1301 ^ r1423;
  wire _9752 = r1571 ^ r1586;
  wire _9753 = _9751 ^ _9752;
  wire _9754 = r1613 ^ r1716;
  wire _9755 = r1809 ^ r1871;
  wire _9756 = _9754 ^ _9755;
  wire _9757 = _9753 ^ _9756;
  wire _9758 = _9750 ^ _9757;
  wire _9759 = _9743 ^ _9758;
  wire _9760 = r6 ^ r80;
  wire _9761 = r115 ^ r209;
  wire _9762 = _9760 ^ _9761;
  wire _9763 = r276 ^ r323;
  wire _9764 = r342 ^ r443;
  wire _9765 = _9763 ^ _9764;
  wire _9766 = _9762 ^ _9765;
  wire _9767 = r501 ^ r533;
  wire _9768 = r588 ^ r636;
  wire _9769 = _9767 ^ _9768;
  wire _9770 = r707 ^ r733;
  wire _9771 = r813 ^ r844;
  wire _9772 = _9770 ^ _9771;
  wire _9773 = _9769 ^ _9772;
  wire _9774 = _9766 ^ _9773;
  wire _9775 = r906 ^ r974;
  wire _9776 = r1104 ^ r1112;
  wire _9777 = _9775 ^ _9776;
  wire _9778 = r1133 ^ r1170;
  wire _9779 = r1258 ^ r1292;
  wire _9780 = _9778 ^ _9779;
  wire _9781 = _9777 ^ _9780;
  wire _9782 = r1338 ^ r1436;
  wire _9783 = r1505 ^ r1604;
  wire _9784 = _9782 ^ _9783;
  wire _9785 = r1626 ^ r1685;
  wire _9786 = r1702 ^ r1798;
  wire _9787 = _9785 ^ _9786;
  wire _9788 = _9784 ^ _9787;
  wire _9789 = _9781 ^ _9788;
  wire _9790 = _9774 ^ _9789;
  wire _9791 = _9759 | _9790;
  wire _9792 = r5 ^ r87;
  wire _9793 = r136 ^ r174;
  wire _9794 = _9792 ^ _9793;
  wire _9795 = r402 ^ r448;
  wire _9796 = r531 ^ r564;
  wire _9797 = _9795 ^ _9796;
  wire _9798 = _9794 ^ _9797;
  wire _9799 = r663 ^ r684;
  wire _9800 = r815 ^ r909;
  wire _9801 = _9799 ^ _9800;
  wire _9802 = r1030 ^ r1156;
  wire _9803 = r1200 ^ r1244;
  wire _9804 = _9802 ^ _9803;
  wire _9805 = _9801 ^ _9804;
  wire _9806 = _9798 ^ _9805;
  wire _9807 = r1312 ^ r1387;
  wire _9808 = r1462 ^ r1536;
  wire _9809 = _9807 ^ _9808;
  wire _9810 = r1623 ^ r1667;
  wire _9811 = r1732 ^ r1861;
  wire _9812 = _9810 ^ _9811;
  wire _9813 = _9809 ^ _9812;
  wire _9814 = r1876 ^ r1878;
  wire _9815 = r1887 ^ r1890;
  wire _9816 = _9814 ^ _9815;
  wire _9817 = r1942 ^ r1944;
  wire _9818 = r2016 ^ r2026;
  wire _9819 = _9817 ^ _9818;
  wire _9820 = _9816 ^ _9819;
  wire _9821 = _9813 ^ _9820;
  wire _9822 = _9806 ^ _9821;
  wire _9823 = r4 ^ r107;
  wire _9824 = r145 ^ r202;
  wire _9825 = _9823 ^ _9824;
  wire _9826 = r230 ^ r302;
  wire _9827 = r366 ^ r395;
  wire _9828 = _9826 ^ _9827;
  wire _9829 = _9825 ^ _9828;
  wire _9830 = r494 ^ r510;
  wire _9831 = r574 ^ r649;
  wire _9832 = _9830 ^ _9831;
  wire _9833 = r719 ^ r752;
  wire _9834 = r785 ^ r879;
  wire _9835 = _9833 ^ _9834;
  wire _9836 = _9832 ^ _9835;
  wire _9837 = _9829 ^ _9836;
  wire _9838 = r893 ^ r996;
  wire _9839 = r1025 ^ r1091;
  wire _9840 = _9838 ^ _9839;
  wire _9841 = r1154 ^ r1318;
  wire _9842 = r1470 ^ r1521;
  wire _9843 = _9841 ^ _9842;
  wire _9844 = _9840 ^ _9843;
  wire _9845 = r1537 ^ r1637;
  wire _9846 = r1665 ^ r1745;
  wire _9847 = _9845 ^ _9846;
  wire _9848 = r1748 ^ r1923;
  wire _9849 = r1932 ^ r1940;
  wire _9850 = _9848 ^ _9849;
  wire _9851 = _9847 ^ _9850;
  wire _9852 = _9844 ^ _9851;
  wire _9853 = _9837 ^ _9852;
  wire _9854 = _9822 | _9853;
  wire _9855 = _9791 | _9854;
  wire _9856 = r140 ^ r199;
  wire _9857 = r251 ^ r311;
  wire _9858 = _9856 ^ _9857;
  wire _9859 = r336 ^ r426;
  wire _9860 = r475 ^ r547;
  wire _9861 = _9859 ^ _9860;
  wire _9862 = _9858 ^ _9861;
  wire _9863 = r568 ^ r669;
  wire _9864 = r726 ^ r821;
  wire _9865 = _9863 ^ _9864;
  wire _9866 = r876 ^ r926;
  wire _9867 = r1008 ^ r1063;
  wire _9868 = _9866 ^ _9867;
  wire _9869 = _9865 ^ _9868;
  wire _9870 = _9862 ^ _9869;
  wire _9871 = r1131 ^ r1241;
  wire _9872 = r1280 ^ r1392;
  wire _9873 = _9871 ^ _9872;
  wire _9874 = r1438 ^ r1503;
  wire _9875 = r1597 ^ r1674;
  wire _9876 = _9874 ^ _9875;
  wire _9877 = _9873 ^ _9876;
  wire _9878 = r1703 ^ r1741;
  wire _9879 = r1930 ^ r1946;
  wire _9880 = _9878 ^ _9879;
  wire _9881 = r1966 ^ r1979;
  wire _9882 = r2018 ^ r2024;
  wire _9883 = _9881 ^ _9882;
  wire _9884 = _9880 ^ _9883;
  wire _9885 = _9877 ^ _9884;
  wire _9886 = _9870 ^ _9885;
  wire _9887 = r3 ^ r86;
  wire _9888 = r146 ^ r214;
  wire _9889 = _9887 ^ _9888;
  wire _9890 = r265 ^ r307;
  wire _9891 = r384 ^ r437;
  wire _9892 = _9890 ^ _9891;
  wire _9893 = _9889 ^ _9892;
  wire _9894 = r458 ^ r550;
  wire _9895 = r571 ^ r664;
  wire _9896 = _9894 ^ _9895;
  wire _9897 = r710 ^ r740;
  wire _9898 = r779 ^ r839;
  wire _9899 = _9897 ^ _9898;
  wire _9900 = _9896 ^ _9899;
  wire _9901 = _9893 ^ _9900;
  wire _9902 = r889 ^ r995;
  wire _9903 = r1015 ^ r1097;
  wire _9904 = _9902 ^ _9903;
  wire _9905 = r1177 ^ r1268;
  wire _9906 = r1304 ^ r1370;
  wire _9907 = _9905 ^ _9906;
  wire _9908 = _9904 ^ _9907;
  wire _9909 = r1420 ^ r1427;
  wire _9910 = r1481 ^ r1513;
  wire _9911 = _9909 ^ _9910;
  wire _9912 = r1715 ^ r1730;
  wire _9913 = r1742 ^ r1872;
  wire _9914 = _9912 ^ _9913;
  wire _9915 = _9911 ^ _9914;
  wire _9916 = _9908 ^ _9915;
  wire _9917 = _9901 ^ _9916;
  wire _9918 = _9886 | _9917;
  wire _9919 = r2 ^ r65;
  wire _9920 = r135 ^ r261;
  wire _9921 = _9919 ^ _9920;
  wire _9922 = r312 ^ r369;
  wire _9923 = r430 ^ r470;
  wire _9924 = _9922 ^ _9923;
  wire _9925 = _9921 ^ _9924;
  wire _9926 = r534 ^ r561;
  wire _9927 = r653 ^ r685;
  wire _9928 = _9926 ^ _9927;
  wire _9929 = r786 ^ r861;
  wire _9930 = r917 ^ r990;
  wire _9931 = _9929 ^ _9930;
  wire _9932 = _9928 ^ _9931;
  wire _9933 = _9925 ^ _9932;
  wire _9934 = r1036 ^ r1202;
  wire _9935 = r1219 ^ r1253;
  wire _9936 = _9934 ^ _9935;
  wire _9937 = r1417 ^ r1506;
  wire _9938 = r1527 ^ r1694;
  wire _9939 = _9937 ^ _9938;
  wire _9940 = _9936 ^ _9939;
  wire _9941 = r1819 ^ r1828;
  wire _9942 = r1860 ^ r1879;
  wire _9943 = _9941 ^ _9942;
  wire _9944 = r1909 ^ r1937;
  wire _9945 = r1957 ^ r1967;
  wire _9946 = _9944 ^ _9945;
  wire _9947 = _9943 ^ _9946;
  wire _9948 = _9940 ^ _9947;
  wire _9949 = _9933 ^ _9948;
  wire _9950 = r1 ^ r68;
  wire _9951 = r160 ^ r225;
  wire _9952 = _9950 ^ _9951;
  wire _9953 = r301 ^ r387;
  wire _9954 = r434 ^ r480;
  wire _9955 = _9953 ^ _9954;
  wire _9956 = _9952 ^ _9955;
  wire _9957 = r511 ^ r596;
  wire _9958 = r617 ^ r706;
  wire _9959 = _9957 ^ _9958;
  wire _9960 = r747 ^ r814;
  wire _9961 = r862 ^ r902;
  wire _9962 = _9960 ^ _9961;
  wire _9963 = _9959 ^ _9962;
  wire _9964 = _9956 ^ _9963;
  wire _9965 = r971 ^ r1034;
  wire _9966 = r1064 ^ r1157;
  wire _9967 = _9965 ^ _9966;
  wire _9968 = r1193 ^ r1221;
  wire _9969 = r1310 ^ r1344;
  wire _9970 = _9968 ^ _9969;
  wire _9971 = _9967 ^ _9970;
  wire _9972 = r1466 ^ r1523;
  wire _9973 = r1660 ^ r1750;
  wire _9974 = _9972 ^ _9973;
  wire _9975 = r1760 ^ r1804;
  wire _9976 = r1899 ^ r1913;
  wire _9977 = _9975 ^ _9976;
  wire _9978 = _9974 ^ _9977;
  wire _9979 = _9971 ^ _9978;
  wire _9980 = _9964 ^ _9979;
  wire _9981 = _9949 | _9980;
  wire _9982 = _9918 | _9981;
  wire _9983 = _9855 | _9982;
  wire _9984 = r0 ^ r108;
  wire _9985 = r167 ^ r246;
  wire _9986 = _9984 ^ _9985;
  wire _9987 = r326 ^ r348;
  wire _9988 = r452 ^ r530;
  wire _9989 = _9987 ^ _9988;
  wire _9990 = _9986 ^ _9989;
  wire _9991 = r580 ^ r645;
  wire _9992 = r770 ^ r827;
  wire _9993 = _9991 ^ _9992;
  wire _9994 = r838 ^ r927;
  wire _9995 = r979 ^ r1090;
  wire _9996 = _9994 ^ _9995;
  wire _9997 = _9993 ^ _9996;
  wire _9998 = _9990 ^ _9997;
  wire _9999 = r1132 ^ r1182;
  wire _10000 = r1270 ^ r1322;
  wire _10001 = _9999 ^ _10000;
  wire _10002 = r1342 ^ r1425;
  wire _10003 = r1446 ^ r1482;
  wire _10004 = _10002 ^ _10003;
  wire _10005 = _10001 ^ _10004;
  wire _10006 = r1645 ^ r1655;
  wire _10007 = r1698 ^ r1729;
  wire _10008 = _10006 ^ _10007;
  wire _10009 = r1925 ^ r1969;
  wire _10010 = r2021 ^ r2027;
  wire _10011 = _10009 ^ _10010;
  wire _10012 = _10008 ^ _10011;
  wire _10013 = _10005 ^ _10012;
  wire _10014 = _9998 ^ _10013;
  wire _10015 = r150 ^ r188;
  wire _10016 = r247 ^ r356;
  wire _10017 = _10015 ^ _10016;
  wire _10018 = r403 ^ r496;
  wire _10019 = r642 ^ r728;
  wire _10020 = _10018 ^ _10019;
  wire _10021 = _10017 ^ _10020;
  wire _10022 = r886 ^ r919;
  wire _10023 = r1001 ^ r1050;
  wire _10024 = _10022 ^ _10023;
  wire _10025 = r1103 ^ r1278;
  wire _10026 = r1376 ^ r1400;
  wire _10027 = _10025 ^ _10026;
  wire _10028 = _10024 ^ _10027;
  wire _10029 = _10021 ^ _10028;
  wire _10030 = r1489 ^ r1528;
  wire _10031 = r1596 ^ r1710;
  wire _10032 = _10030 ^ _10031;
  wire _10033 = r1723 ^ r1814;
  wire _10034 = r1830 ^ r1881;
  wire _10035 = _10033 ^ _10034;
  wire _10036 = _10032 ^ _10035;
  wire _10037 = r1919 ^ r1953;
  wire _10038 = r1973 ^ r1983;
  wire _10039 = _10037 ^ _10038;
  wire _10040 = r2022 ^ r2034;
  wire _10041 = r2038 ^ r2044;
  wire _10042 = _10040 ^ _10041;
  wire _10043 = _10039 ^ _10042;
  wire _10044 = _10036 ^ _10043;
  wire _10045 = _10029 ^ _10044;
  wire _10046 = _10014 | _10045;
  wire _10047 = r191 ^ r278;
  wire _10048 = r316 ^ r352;
  wire _10049 = _10047 ^ _10048;
  wire _10050 = r442 ^ r483;
  wire _10051 = r543 ^ r602;
  wire _10052 = _10050 ^ _10051;
  wire _10053 = _10049 ^ _10052;
  wire _10054 = r656 ^ r687;
  wire _10055 = r781 ^ r848;
  wire _10056 = _10054 ^ _10055;
  wire _10057 = r907 ^ r1053;
  wire _10058 = r1123 ^ r1357;
  wire _10059 = _10057 ^ _10058;
  wire _10060 = _10056 ^ _10059;
  wire _10061 = _10053 ^ _10060;
  wire _10062 = r1389 ^ r1411;
  wire _10063 = r1461 ^ r1556;
  wire _10064 = _10062 ^ _10063;
  wire _10065 = r1648 ^ r1651;
  wire _10066 = r1717 ^ r1749;
  wire _10067 = _10065 ^ _10066;
  wire _10068 = _10064 ^ _10067;
  wire _10069 = r1836 ^ r1853;
  wire _10070 = r1907 ^ r1926;
  wire _10071 = _10069 ^ _10070;
  wire _10072 = r1928 ^ r1938;
  wire _10073 = r1958 ^ r1968;
  wire _10074 = _10072 ^ _10073;
  wire _10075 = _10071 ^ _10074;
  wire _10076 = _10068 ^ _10075;
  wire _10077 = _10061 ^ _10076;
  wire _10078 = r78 ^ r119;
  wire _10079 = r183 ^ r271;
  wire _10080 = _10078 ^ _10079;
  wire _10081 = r318 ^ r357;
  wire _10082 = r399 ^ r499;
  wire _10083 = _10081 ^ _10082;
  wire _10084 = _10080 ^ _10083;
  wire _10085 = r513 ^ r575;
  wire _10086 = r651 ^ r678;
  wire _10087 = _10085 ^ _10086;
  wire _10088 = r743 ^ r802;
  wire _10089 = r853 ^ r924;
  wire _10090 = _10088 ^ _10089;
  wire _10091 = _10087 ^ _10090;
  wire _10092 = _10084 ^ _10091;
  wire _10093 = r977 ^ r1037;
  wire _10094 = r1111 ^ r1172;
  wire _10095 = _10093 ^ _10094;
  wire _10096 = r1249 ^ r1317;
  wire _10097 = r1359 ^ r1404;
  wire _10098 = _10096 ^ _10097;
  wire _10099 = _10095 ^ _10098;
  wire _10100 = r1447 ^ r1457;
  wire _10101 = r1488 ^ r1511;
  wire _10102 = _10100 ^ _10101;
  wire _10103 = r1675 ^ r1714;
  wire _10104 = r1722 ^ r1799;
  wire _10105 = _10103 ^ _10104;
  wire _10106 = _10102 ^ _10105;
  wire _10107 = _10099 ^ _10106;
  wire _10108 = _10092 ^ _10107;
  wire _10109 = _10077 | _10108;
  wire _10110 = _10046 | _10109;
  wire _10111 = r61 ^ r158;
  wire _10112 = r234 ^ r288;
  wire _10113 = _10111 ^ _10112;
  wire _10114 = r347 ^ r560;
  wire _10115 = r563 ^ r625;
  wire _10116 = _10114 ^ _10115;
  wire _10117 = _10113 ^ _10116;
  wire _10118 = r720 ^ r764;
  wire _10119 = r816 ^ r898;
  wire _10120 = _10118 ^ _10119;
  wire _10121 = r956 ^ r1014;
  wire _10122 = r1080 ^ r1134;
  wire _10123 = _10121 ^ _10122;
  wire _10124 = _10120 ^ _10123;
  wire _10125 = _10117 ^ _10124;
  wire _10126 = r1186 ^ r1220;
  wire _10127 = r1246 ^ r1293;
  wire _10128 = _10126 ^ _10127;
  wire _10129 = r1345 ^ r1408;
  wire _10130 = r1501 ^ r1569;
  wire _10131 = _10129 ^ _10130;
  wire _10132 = _10128 ^ _10131;
  wire _10133 = r1664 ^ r1721;
  wire _10134 = r1727 ^ r1754;
  wire _10135 = _10133 ^ _10134;
  wire _10136 = r1961 ^ r2014;
  wire _10137 = r2035 ^ r2039;
  wire _10138 = _10136 ^ _10137;
  wire _10139 = _10135 ^ _10138;
  wire _10140 = _10132 ^ _10139;
  wire _10141 = _10125 ^ _10140;
  wire _10142 = r88 ^ r238;
  wire _10143 = r324 ^ r372;
  wire _10144 = _10142 ^ _10143;
  wire _10145 = r472 ^ r548;
  wire _10146 = r604 ^ r634;
  wire _10147 = _10145 ^ _10146;
  wire _10148 = _10144 ^ _10147;
  wire _10149 = r683 ^ r765;
  wire _10150 = r812 ^ r852;
  wire _10151 = _10149 ^ _10150;
  wire _10152 = r895 ^ r959;
  wire _10153 = r1092 ^ r1125;
  wire _10154 = _10152 ^ _10153;
  wire _10155 = _10151 ^ _10154;
  wire _10156 = _10148 ^ _10155;
  wire _10157 = r1179 ^ r1261;
  wire _10158 = r1325 ^ r1332;
  wire _10159 = _10157 ^ _10158;
  wire _10160 = r1377 ^ r1397;
  wire _10161 = r1719 ^ r1775;
  wire _10162 = _10160 ^ _10161;
  wire _10163 = _10159 ^ _10162;
  wire _10164 = r1811 ^ r1839;
  wire _10165 = r1939 ^ r1952;
  wire _10166 = _10164 ^ _10165;
  wire _10167 = r1960 ^ r1999;
  wire _10168 = r2001 ^ r2012;
  wire _10169 = _10167 ^ _10168;
  wire _10170 = _10166 ^ _10169;
  wire _10171 = _10163 ^ _10170;
  wire _10172 = _10156 ^ _10171;
  wire _10173 = _10141 | _10172;
  wire _10174 = r120 ^ r210;
  wire _10175 = r279 ^ r379;
  wire _10176 = _10174 ^ _10175;
  wire _10177 = r425 ^ r467;
  wire _10178 = r566 ^ r742;
  wire _10179 = _10177 ^ _10178;
  wire _10180 = _10176 ^ _10179;
  wire _10181 = r846 ^ r911;
  wire _10182 = r1002 ^ r1006;
  wire _10183 = _10181 ^ _10182;
  wire _10184 = r1059 ^ r1210;
  wire _10185 = r1295 ^ r1341;
  wire _10186 = _10184 ^ _10185;
  wire _10187 = _10183 ^ _10186;
  wire _10188 = _10180 ^ _10187;
  wire _10189 = r1540 ^ r1566;
  wire _10190 = r1598 ^ r1634;
  wire _10191 = _10189 ^ _10190;
  wire _10192 = r1720 ^ r1805;
  wire _10193 = r1837 ^ r1877;
  wire _10194 = _10192 ^ _10193;
  wire _10195 = _10191 ^ _10194;
  wire _10196 = r1935 ^ r1976;
  wire _10197 = r1980 ^ r2005;
  wire _10198 = _10196 ^ _10197;
  wire _10199 = r2008 ^ r2036;
  wire _10200 = r2037 ^ r2045;
  wire _10201 = _10199 ^ _10200;
  wire _10202 = _10198 ^ _10201;
  wire _10203 = _10195 ^ _10202;
  wire _10204 = _10188 ^ _10203;
  wire _10205 = r52 ^ r66;
  wire _10206 = r151 ^ r221;
  wire _10207 = _10205 ^ _10206;
  wire _10208 = r237 ^ r289;
  wire _10209 = r361 ^ r411;
  wire _10210 = _10208 ^ _10209;
  wire _10211 = _10207 ^ _10210;
  wire _10212 = r473 ^ r539;
  wire _10213 = r585 ^ r631;
  wire _10214 = _10212 ^ _10213;
  wire _10215 = r711 ^ r734;
  wire _10216 = r797 ^ r883;
  wire _10217 = _10215 ^ _10216;
  wire _10218 = _10214 ^ _10217;
  wire _10219 = _10211 ^ _10218;
  wire _10220 = r904 ^ r978;
  wire _10221 = r1046 ^ r1106;
  wire _10222 = _10220 ^ _10221;
  wire _10223 = r1130 ^ r1231;
  wire _10224 = r1305 ^ r1368;
  wire _10225 = _10223 ^ _10224;
  wire _10226 = _10222 ^ _10225;
  wire _10227 = r1416 ^ r1475;
  wire _10228 = r1485 ^ r1515;
  wire _10229 = _10227 ^ _10228;
  wire _10230 = r1595 ^ r1661;
  wire _10231 = r1695 ^ r1800;
  wire _10232 = _10230 ^ _10231;
  wire _10233 = _10229 ^ _10232;
  wire _10234 = _10226 ^ _10233;
  wire _10235 = _10219 ^ _10234;
  wire _10236 = _10204 | _10235;
  wire _10237 = _10173 | _10236;
  wire _10238 = _10110 | _10237;
  wire _10239 = _9983 | _10238;
  wire _10240 = _9728 | _10239;
  wire _10241 = _9217 | _10240;
  wire _10242 = r53 ^ r126;
  wire _10243 = r196 ^ r295;
  wire _10244 = _10242 ^ _10243;
  wire _10245 = r338 ^ r439;
  wire _10246 = r454 ^ r531;
  wire _10247 = _10245 ^ _10246;
  wire _10248 = _10244 ^ _10247;
  wire _10249 = r577 ^ r637;
  wire _10250 = r707 ^ r759;
  wire _10251 = _10249 ^ _10250;
  wire _10252 = r792 ^ r856;
  wire _10253 = r890 ^ r1034;
  wire _10254 = _10252 ^ _10253;
  wire _10255 = _10251 ^ _10254;
  wire _10256 = _10248 ^ _10255;
  wire _10257 = r1070 ^ r1154;
  wire _10258 = r1342 ^ r1413;
  wire _10259 = _10257 ^ _10258;
  wire _10260 = r1453 ^ r1484;
  wire _10261 = r1572 ^ r1579;
  wire _10262 = _10260 ^ _10261;
  wire _10263 = _10259 ^ _10262;
  wire _10264 = r1662 ^ r1725;
  wire _10265 = r1741 ^ r1761;
  wire _10266 = _10264 ^ _10265;
  wire _10267 = r1816 ^ r1836;
  wire _10268 = r1856 ^ r1895;
  wire _10269 = _10267 ^ _10268;
  wire _10270 = _10266 ^ _10269;
  wire _10271 = _10263 ^ _10270;
  wire _10272 = _10256 ^ _10271;
  wire _10273 = r51 ^ r65;
  wire _10274 = r150 ^ r220;
  wire _10275 = _10273 ^ _10274;
  wire _10276 = r236 ^ r288;
  wire _10277 = r360 ^ r410;
  wire _10278 = _10276 ^ _10277;
  wire _10279 = _10275 ^ _10278;
  wire _10280 = r472 ^ r538;
  wire _10281 = r584 ^ r630;
  wire _10282 = _10280 ^ _10281;
  wire _10283 = r733 ^ r882;
  wire _10284 = r903 ^ r977;
  wire _10285 = _10283 ^ _10284;
  wire _10286 = _10282 ^ _10285;
  wire _10287 = _10279 ^ _10286;
  wire _10288 = r1045 ^ r1105;
  wire _10289 = r1217 ^ r1230;
  wire _10290 = _10288 ^ _10289;
  wire _10291 = r1304 ^ r1367;
  wire _10292 = r1474 ^ r1558;
  wire _10293 = _10291 ^ _10292;
  wire _10294 = _10290 ^ _10293;
  wire _10295 = r1594 ^ r1660;
  wire _10296 = r1759 ^ r1831;
  wire _10297 = _10295 ^ _10296;
  wire _10298 = r1929 ^ r1992;
  wire _10299 = r2003 ^ r2013;
  wire _10300 = _10298 ^ _10299;
  wire _10301 = _10297 ^ _10300;
  wire _10302 = _10294 ^ _10301;
  wire _10303 = _10287 ^ _10302;
  wire _10304 = _10272 | _10303;
  wire _10305 = r50 ^ r84;
  wire _10306 = r165 ^ r231;
  wire _10307 = _10305 ^ _10306;
  wire _10308 = r316 ^ r362;
  wire _10309 = r427 ^ r462;
  wire _10310 = _10308 ^ _10309;
  wire _10311 = _10307 ^ _10310;
  wire _10312 = r535 ^ r592;
  wire _10313 = r623 ^ r749;
  wire _10314 = _10312 ^ _10313;
  wire _10315 = r797 ^ r834;
  wire _10316 = r932 ^ r998;
  wire _10317 = _10315 ^ _10316;
  wire _10318 = _10314 ^ _10317;
  wire _10319 = _10311 ^ _10318;
  wire _10320 = r1015 ^ r1060;
  wire _10321 = r1075 ^ r1161;
  wire _10322 = _10320 ^ _10321;
  wire _10323 = r1302 ^ r1353;
  wire _10324 = r1463 ^ r1492;
  wire _10325 = _10323 ^ _10324;
  wire _10326 = _10322 ^ _10325;
  wire _10327 = r1537 ^ r1756;
  wire _10328 = r1813 ^ r1868;
  wire _10329 = _10327 ^ _10328;
  wire _10330 = r1878 ^ r1911;
  wire _10331 = r1953 ^ r1969;
  wire _10332 = _10330 ^ _10331;
  wire _10333 = _10329 ^ _10332;
  wire _10334 = _10326 ^ _10333;
  wire _10335 = _10319 ^ _10334;
  wire _10336 = r56 ^ r136;
  wire _10337 = r184 ^ r268;
  wire _10338 = _10336 ^ _10337;
  wire _10339 = r330 ^ r390;
  wire _10340 = r392 ^ r484;
  wire _10341 = _10339 ^ _10340;
  wire _10342 = _10338 ^ _10341;
  wire _10343 = r552 ^ r588;
  wire _10344 = r656 ^ r717;
  wire _10345 = _10343 ^ _10344;
  wire _10346 = r754 ^ r828;
  wire _10347 = r967 ^ r1007;
  wire _10348 = _10346 ^ _10347;
  wire _10349 = _10345 ^ _10348;
  wire _10350 = _10342 ^ _10349;
  wire _10351 = r1076 ^ r1158;
  wire _10352 = r1221 ^ r1234;
  wire _10353 = _10351 ^ _10352;
  wire _10354 = r1319 ^ r1546;
  wire _10355 = r1573 ^ r1583;
  wire _10356 = _10354 ^ _10355;
  wire _10357 = _10353 ^ _10356;
  wire _10358 = r1631 ^ r1701;
  wire _10359 = r1783 ^ r1832;
  wire _10360 = _10358 ^ _10359;
  wire _10361 = r1833 ^ r1846;
  wire _10362 = r1860 ^ r1896;
  wire _10363 = _10361 ^ _10362;
  wire _10364 = _10360 ^ _10363;
  wire _10365 = _10357 ^ _10364;
  wire _10366 = _10350 ^ _10365;
  wire _10367 = _10335 | _10366;
  wire _10368 = _10304 | _10367;
  wire _10369 = r49 ^ r109;
  wire _10370 = r113 ^ r223;
  wire _10371 = _10369 ^ _10370;
  wire _10372 = r273 ^ r302;
  wire _10373 = r369 ^ r400;
  wire _10374 = _10372 ^ _10373;
  wire _10375 = _10371 ^ _10374;
  wire _10376 = r490 ^ r544;
  wire _10377 = r593 ^ r640;
  wire _10378 = _10376 ^ _10377;
  wire _10379 = r693 ^ r821;
  wire _10380 = r855 ^ r936;
  wire _10381 = _10379 ^ _10380;
  wire _10382 = _10378 ^ _10381;
  wire _10383 = _10375 ^ _10382;
  wire _10384 = r951 ^ r1050;
  wire _10385 = r1104 ^ r1116;
  wire _10386 = _10384 ^ _10385;
  wire _10387 = r1169 ^ r1206;
  wire _10388 = r1237 ^ r1288;
  wire _10389 = _10387 ^ _10388;
  wire _10390 = _10386 ^ _10389;
  wire _10391 = r1369 ^ r1411;
  wire _10392 = r1427 ^ r1499;
  wire _10393 = _10391 ^ _10392;
  wire _10394 = r1614 ^ r1653;
  wire _10395 = r1704 ^ r1801;
  wire _10396 = _10394 ^ _10395;
  wire _10397 = _10393 ^ _10396;
  wire _10398 = _10390 ^ _10397;
  wire _10399 = _10383 ^ _10398;
  wire _10400 = r48 ^ r70;
  wire _10401 = r137 ^ r185;
  wire _10402 = _10400 ^ _10401;
  wire _10403 = r242 ^ r284;
  wire _10404 = r382 ^ r395;
  wire _10405 = _10403 ^ _10404;
  wire _10406 = _10402 ^ _10405;
  wire _10407 = r476 ^ r518;
  wire _10408 = r583 ^ r653;
  wire _10409 = _10407 ^ _10408;
  wire _10410 = r704 ^ r753;
  wire _10411 = r784 ^ r832;
  wire _10412 = _10410 ^ _10411;
  wire _10413 = _10409 ^ _10412;
  wire _10414 = _10406 ^ _10413;
  wire _10415 = r940 ^ r979;
  wire _10416 = r1012 ^ r1097;
  wire _10417 = _10415 ^ _10416;
  wire _10418 = r1186 ^ r1227;
  wire _10419 = r1289 ^ r1357;
  wire _10420 = _10418 ^ _10419;
  wire _10421 = _10417 ^ _10420;
  wire _10422 = r1398 ^ r1436;
  wire _10423 = r1462 ^ r1512;
  wire _10424 = _10422 ^ _10423;
  wire _10425 = r1554 ^ r1617;
  wire _10426 = r1718 ^ r1802;
  wire _10427 = _10425 ^ _10426;
  wire _10428 = _10424 ^ _10427;
  wire _10429 = _10421 ^ _10428;
  wire _10430 = _10414 ^ _10429;
  wire _10431 = _10399 | _10430;
  wire _10432 = r47 ^ r62;
  wire _10433 = r203 ^ r241;
  wire _10434 = _10432 ^ _10433;
  wire _10435 = r304 ^ r527;
  wire _10436 = r606 ^ r663;
  wire _10437 = _10435 ^ _10436;
  wire _10438 = _10434 ^ _10437;
  wire _10439 = r697 ^ r722;
  wire _10440 = r748 ^ r788;
  wire _10441 = _10439 ^ _10440;
  wire _10442 = r867 ^ r969;
  wire _10443 = r1041 ^ r1061;
  wire _10444 = _10442 ^ _10443;
  wire _10445 = _10441 ^ _10444;
  wire _10446 = _10438 ^ _10445;
  wire _10447 = r1140 ^ r1170;
  wire _10448 = r1261 ^ r1318;
  wire _10449 = _10447 ^ _10448;
  wire _10450 = r1374 ^ r1485;
  wire _10451 = r1548 ^ r1569;
  wire _10452 = _10450 ^ _10451;
  wire _10453 = _10449 ^ _10452;
  wire _10454 = r1671 ^ r1764;
  wire _10455 = r1827 ^ r1909;
  wire _10456 = _10454 ^ _10455;
  wire _10457 = r1922 ^ r1926;
  wire _10458 = r1972 ^ r1981;
  wire _10459 = _10457 ^ _10458;
  wire _10460 = _10456 ^ _10459;
  wire _10461 = _10453 ^ _10460;
  wire _10462 = _10446 ^ _10461;
  wire _10463 = r46 ^ r94;
  wire _10464 = r148 ^ r211;
  wire _10465 = _10463 ^ _10464;
  wire _10466 = r272 ^ r318;
  wire _10467 = r361 ^ r446;
  wire _10468 = _10466 ^ _10467;
  wire _10469 = _10465 ^ _10468;
  wire _10470 = r502 ^ r521;
  wire _10471 = r612 ^ r634;
  wire _10472 = _10470 ^ _10471;
  wire _10473 = r701 ^ r777;
  wire _10474 = r870 ^ r911;
  wire _10475 = _10473 ^ _10474;
  wire _10476 = _10472 ^ _10475;
  wire _10477 = _10469 ^ _10476;
  wire _10478 = r956 ^ r1038;
  wire _10479 = r1066 ^ r1151;
  wire _10480 = _10478 ^ _10479;
  wire _10481 = r1182 ^ r1244;
  wire _10482 = r1310 ^ r1349;
  wire _10483 = _10481 ^ _10482;
  wire _10484 = _10480 ^ _10483;
  wire _10485 = r1401 ^ r1456;
  wire _10486 = r1479 ^ r1500;
  wire _10487 = _10485 ^ _10486;
  wire _10488 = r1632 ^ r1699;
  wire _10489 = r1730 ^ r1873;
  wire _10490 = _10488 ^ _10489;
  wire _10491 = _10487 ^ _10490;
  wire _10492 = _10484 ^ _10491;
  wire _10493 = _10477 ^ _10492;
  wire _10494 = _10462 | _10493;
  wire _10495 = _10431 | _10494;
  wire _10496 = _10368 | _10495;
  wire _10497 = r45 ^ r103;
  wire _10498 = r168 ^ r314;
  wire _10499 = _10497 ^ _10498;
  wire _10500 = r377 ^ r413;
  wire _10501 = r483 ^ r524;
  wire _10502 = _10500 ^ _10501;
  wire _10503 = _10499 ^ _10502;
  wire _10504 = r597 ^ r690;
  wire _10505 = r737 ^ r787;
  wire _10506 = _10504 ^ _10505;
  wire _10507 = r857 ^ r893;
  wire _10508 = r975 ^ r1055;
  wire _10509 = _10507 ^ _10508;
  wire _10510 = _10506 ^ _10509;
  wire _10511 = _10503 ^ _10510;
  wire _10512 = r1144 ^ r1328;
  wire _10513 = r1346 ^ r1421;
  wire _10514 = _10512 ^ _10513;
  wire _10515 = r1439 ^ r1486;
  wire _10516 = r1491 ^ r1509;
  wire _10517 = _10515 ^ _10516;
  wire _10518 = _10514 ^ _10517;
  wire _10519 = r1672 ^ r1688;
  wire _10520 = r1742 ^ r1796;
  wire _10521 = _10519 ^ _10520;
  wire _10522 = r1814 ^ r1936;
  wire _10523 = r1946 ^ r1957;
  wire _10524 = _10522 ^ _10523;
  wire _10525 = _10521 ^ _10524;
  wire _10526 = _10518 ^ _10525;
  wire _10527 = _10511 ^ _10526;
  wire _10528 = r44 ^ r97;
  wire _10529 = r131 ^ r212;
  wire _10530 = _10528 ^ _10529;
  wire _10531 = r255 ^ r280;
  wire _10532 = r348 ^ r420;
  wire _10533 = _10531 ^ _10532;
  wire _10534 = _10530 ^ _10533;
  wire _10535 = r494 ^ r516;
  wire _10536 = r599 ^ r665;
  wire _10537 = _10535 ^ _10536;
  wire _10538 = r671 ^ r760;
  wire _10539 = r782 ^ r833;
  wire _10540 = _10538 ^ _10539;
  wire _10541 = _10537 ^ _10540;
  wire _10542 = _10534 ^ _10541;
  wire _10543 = r907 ^ r947;
  wire _10544 = r1047 ^ r1065;
  wire _10545 = _10543 ^ _10544;
  wire _10546 = r1148 ^ r1268;
  wire _10547 = r1278 ^ r1361;
  wire _10548 = _10546 ^ _10547;
  wire _10549 = _10545 ^ _10548;
  wire _10550 = r1515 ^ r1530;
  wire _10551 = r1538 ^ r1560;
  wire _10552 = _10550 ^ _10551;
  wire _10553 = r1607 ^ r1626;
  wire _10554 = r1667 ^ r1803;
  wire _10555 = _10553 ^ _10554;
  wire _10556 = _10552 ^ _10555;
  wire _10557 = _10549 ^ _10556;
  wire _10558 = _10542 ^ _10557;
  wire _10559 = _10527 | _10558;
  wire _10560 = r43 ^ r101;
  wire _10561 = r132 ^ r202;
  wire _10562 = _10560 ^ _10561;
  wire _10563 = r243 ^ r385;
  wire _10564 = r404 ^ r503;
  wire _10565 = _10563 ^ _10564;
  wire _10566 = _10562 ^ _10565;
  wire _10567 = r553 ^ r569;
  wire _10568 = r626 ^ r710;
  wire _10569 = _10567 ^ _10568;
  wire _10570 = r758 ^ r819;
  wire _10571 = r917 ^ r944;
  wire _10572 = _10570 ^ _10571;
  wire _10573 = _10569 ^ _10572;
  wire _10574 = _10566 ^ _10573;
  wire _10575 = r1022 ^ r1138;
  wire _10576 = r1208 ^ r1240;
  wire _10577 = _10575 ^ _10576;
  wire _10578 = r1384 ^ r1425;
  wire _10579 = r1483 ^ r1508;
  wire _10580 = _10578 ^ _10579;
  wire _10581 = _10577 ^ _10580;
  wire _10582 = r1532 ^ r1684;
  wire _10583 = r1747 ^ r1795;
  wire _10584 = _10582 ^ _10583;
  wire _10585 = r1823 ^ r1865;
  wire _10586 = r1867 ^ r1897;
  wire _10587 = _10585 ^ _10586;
  wire _10588 = _10584 ^ _10587;
  wire _10589 = _10581 ^ _10588;
  wire _10590 = _10574 ^ _10589;
  wire _10591 = r42 ^ r92;
  wire _10592 = r167 ^ r172;
  wire _10593 = _10591 ^ _10592;
  wire _10594 = r350 ^ r406;
  wire _10595 = r534 ^ r604;
  wire _10596 = _10594 ^ _10595;
  wire _10597 = _10593 ^ _10596;
  wire _10598 = r646 ^ r720;
  wire _10599 = r736 ^ r826;
  wire _10600 = _10598 ^ _10599;
  wire _10601 = r879 ^ r943;
  wire _10602 = r961 ^ r1031;
  wire _10603 = _10601 ^ _10602;
  wire _10604 = _10600 ^ _10603;
  wire _10605 = _10597 ^ _10604;
  wire _10606 = r1117 ^ r1194;
  wire _10607 = r1229 ^ r1428;
  wire _10608 = _10606 ^ _10607;
  wire _10609 = r1449 ^ r1477;
  wire _10610 = r1529 ^ r1533;
  wire _10611 = _10609 ^ _10610;
  wire _10612 = _10608 ^ _10611;
  wire _10613 = r1634 ^ r1650;
  wire _10614 = r1706 ^ r1753;
  wire _10615 = _10613 ^ _10614;
  wire _10616 = r1862 ^ r1963;
  wire _10617 = r1991 ^ r1993;
  wire _10618 = _10616 ^ _10617;
  wire _10619 = _10615 ^ _10618;
  wire _10620 = _10612 ^ _10619;
  wire _10621 = _10605 ^ _10620;
  wire _10622 = _10590 | _10621;
  wire _10623 = _10559 | _10622;
  wire _10624 = r41 ^ r71;
  wire _10625 = r158 ^ r179;
  wire _10626 = _10624 ^ _10625;
  wire _10627 = r240 ^ r363;
  wire _10628 = r431 ^ r489;
  wire _10629 = _10627 ^ _10628;
  wire _10630 = _10626 ^ _10629;
  wire _10631 = r548 ^ r561;
  wire _10632 = r772 ^ r793;
  wire _10633 = _10631 ^ _10632;
  wire _10634 = r865 ^ r931;
  wire _10635 = r953 ^ r1025;
  wire _10636 = _10634 ^ _10635;
  wire _10637 = _10633 ^ _10636;
  wire _10638 = _10630 ^ _10637;
  wire _10639 = r1157 ^ r1211;
  wire _10640 = r1271 ^ r1326;
  wire _10641 = _10639 ^ _10640;
  wire _10642 = r1338 ^ r1389;
  wire _10643 = r1420 ^ r1600;
  wire _10644 = _10642 ^ _10643;
  wire _10645 = _10641 ^ _10644;
  wire _10646 = r1627 ^ r1676;
  wire _10647 = r1724 ^ r1782;
  wire _10648 = _10646 ^ _10647;
  wire _10649 = r1885 ^ r1925;
  wire _10650 = r2022 ^ r2029;
  wire _10651 = _10649 ^ _10650;
  wire _10652 = _10648 ^ _10651;
  wire _10653 = _10645 ^ _10652;
  wire _10654 = _10638 ^ _10653;
  wire _10655 = r108 ^ r117;
  wire _10656 = r215 ^ r265;
  wire _10657 = _10655 ^ _10656;
  wire _10658 = r324 ^ r359;
  wire _10659 = r411 ^ r651;
  wire _10660 = _10658 ^ _10659;
  wire _10661 = _10657 ^ _10660;
  wire _10662 = r774 ^ r835;
  wire _10663 = r920 ^ r986;
  wire _10664 = _10662 ^ _10663;
  wire _10665 = r1071 ^ r1175;
  wire _10666 = r1232 ^ r1308;
  wire _10667 = _10665 ^ _10666;
  wire _10668 = _10664 ^ _10667;
  wire _10669 = _10661 ^ _10668;
  wire _10670 = r1429 ^ r1448;
  wire _10671 = r1458 ^ r1551;
  wire _10672 = _10670 ^ _10671;
  wire _10673 = r1615 ^ r1726;
  wire _10674 = r1776 ^ r1810;
  wire _10675 = _10673 ^ _10674;
  wire _10676 = _10672 ^ _10675;
  wire _10677 = r1820 ^ r1888;
  wire _10678 = r1961 ^ r1980;
  wire _10679 = _10677 ^ _10678;
  wire _10680 = r2018 ^ r2019;
  wire _10681 = r2020 ^ r2034;
  wire _10682 = _10680 ^ _10681;
  wire _10683 = _10679 ^ _10682;
  wire _10684 = _10676 ^ _10683;
  wire _10685 = _10669 ^ _10684;
  wire _10686 = _10654 | _10685;
  wire _10687 = r40 ^ r66;
  wire _10688 = r217 ^ r286;
  wire _10689 = _10687 ^ _10688;
  wire _10690 = r380 ^ r497;
  wire _10691 = r528 ^ r598;
  wire _10692 = _10690 ^ _10691;
  wire _10693 = _10689 ^ _10692;
  wire _10694 = r654 ^ r692;
  wire _10695 = r761 ^ r824;
  wire _10696 = _10694 ^ _10695;
  wire _10697 = r881 ^ r934;
  wire _10698 = r996 ^ r1020;
  wire _10699 = _10697 ^ _10698;
  wire _10700 = _10696 ^ _10699;
  wire _10701 = _10693 ^ _10700;
  wire _10702 = r1069 ^ r1123;
  wire _10703 = r1184 ^ r1250;
  wire _10704 = _10702 ^ _10703;
  wire _10705 = r1314 ^ r1336;
  wire _10706 = r1394 ^ r1443;
  wire _10707 = _10705 ^ _10706;
  wire _10708 = _10704 ^ _10707;
  wire _10709 = r1630 ^ r1712;
  wire _10710 = r1755 ^ r1852;
  wire _10711 = _10709 ^ _10710;
  wire _10712 = r1913 ^ r1997;
  wire _10713 = r2021 ^ r2026;
  wire _10714 = _10712 ^ _10713;
  wire _10715 = _10711 ^ _10714;
  wire _10716 = _10708 ^ _10715;
  wire _10717 = _10701 ^ _10716;
  wire _10718 = r39 ^ r78;
  wire _10719 = r170 ^ r189;
  wire _10720 = _10718 ^ _10719;
  wire _10721 = r274 ^ r291;
  wire _10722 = r343 ^ r432;
  wire _10723 = _10721 ^ _10722;
  wire _10724 = _10720 ^ _10723;
  wire _10725 = r465 ^ r517;
  wire _10726 = r611 ^ r645;
  wire _10727 = _10725 ^ _10726;
  wire _10728 = r679 ^ r804;
  wire _10729 = r868 ^ r899;
  wire _10730 = _10728 ^ _10729;
  wire _10731 = _10727 ^ _10730;
  wire _10732 = _10724 ^ _10731;
  wire _10733 = r990 ^ r1056;
  wire _10734 = r1099 ^ r1152;
  wire _10735 = _10733 ^ _10734;
  wire _10736 = r1179 ^ r1258;
  wire _10737 = r1276 ^ r1285;
  wire _10738 = _10736 ^ _10737;
  wire _10739 = _10735 ^ _10738;
  wire _10740 = r1382 ^ r1441;
  wire _10741 = r1541 ^ r1578;
  wire _10742 = _10740 ^ _10741;
  wire _10743 = r1682 ^ r1845;
  wire _10744 = r1872 ^ r1898;
  wire _10745 = _10743 ^ _10744;
  wire _10746 = _10742 ^ _10745;
  wire _10747 = _10739 ^ _10746;
  wire _10748 = _10732 ^ _10747;
  wire _10749 = _10717 | _10748;
  wire _10750 = _10686 | _10749;
  wire _10751 = _10623 | _10750;
  wire _10752 = _10496 | _10751;
  wire _10753 = r38 ^ r104;
  wire _10754 = r121 ^ r267;
  wire _10755 = _10753 ^ _10754;
  wire _10756 = r332 ^ r344;
  wire _10757 = r405 ^ r477;
  wire _10758 = _10756 ^ _10757;
  wire _10759 = _10755 ^ _10758;
  wire _10760 = r506 ^ r585;
  wire _10761 = r695 ^ r757;
  wire _10762 = _10760 ^ _10761;
  wire _10763 = r806 ^ r831;
  wire _10764 = r909 ^ r993;
  wire _10765 = _10763 ^ _10764;
  wire _10766 = _10762 ^ _10765;
  wire _10767 = _10759 ^ _10766;
  wire _10768 = r1037 ^ r1082;
  wire _10769 = r1139 ^ r1185;
  wire _10770 = _10768 ^ _10769;
  wire _10771 = r1329 ^ r1362;
  wire _10772 = r1471 ^ r1543;
  wire _10773 = _10771 ^ _10772;
  wire _10774 = _10770 ^ _10773;
  wire _10775 = r1605 ^ r1651;
  wire _10776 = r1692 ^ r1740;
  wire _10777 = _10775 ^ _10776;
  wire _10778 = r1850 ^ r1935;
  wire _10779 = r1951 ^ r1970;
  wire _10780 = _10778 ^ _10779;
  wire _10781 = _10777 ^ _10780;
  wire _10782 = _10774 ^ _10781;
  wire _10783 = _10767 ^ _10782;
  wire _10784 = r37 ^ r93;
  wire _10785 = r115 ^ r183;
  wire _10786 = _10784 ^ _10785;
  wire _10787 = r253 ^ r290;
  wire _10788 = r379 ^ r419;
  wire _10789 = _10787 ^ _10788;
  wire _10790 = _10786 ^ _10789;
  wire _10791 = r475 ^ r519;
  wire _10792 = r564 ^ r714;
  wire _10793 = _10791 ^ _10792;
  wire _10794 = r728 ^ r794;
  wire _10795 = r862 ^ r904;
  wire _10796 = _10794 ^ _10795;
  wire _10797 = _10793 ^ _10796;
  wire _10798 = _10790 ^ _10797;
  wire _10799 = r983 ^ r1051;
  wire _10800 = r1085 ^ r1126;
  wire _10801 = _10799 ^ _10800;
  wire _10802 = r1259 ^ r1345;
  wire _10803 = r1405 ^ r1432;
  wire _10804 = _10802 ^ _10803;
  wire _10805 = _10801 ^ _10804;
  wire _10806 = r1454 ^ r1590;
  wire _10807 = r1620 ^ r1656;
  wire _10808 = _10806 ^ _10807;
  wire _10809 = r1705 ^ r1927;
  wire _10810 = r1947 ^ r1958;
  wire _10811 = _10809 ^ _10810;
  wire _10812 = _10808 ^ _10811;
  wire _10813 = _10805 ^ _10812;
  wire _10814 = _10798 ^ _10813;
  wire _10815 = _10783 | _10814;
  wire _10816 = r36 ^ r80;
  wire _10817 = r155 ^ r190;
  wire _10818 = _10816 ^ _10817;
  wire _10819 = r370 ^ r492;
  wire _10820 = r540 ^ r587;
  wire _10821 = _10819 ^ _10820;
  wire _10822 = _10818 ^ _10821;
  wire _10823 = r658 ^ r669;
  wire _10824 = r825 ^ r859;
  wire _10825 = _10823 ^ _10824;
  wire _10826 = r962 ^ r1006;
  wire _10827 = r1072 ^ r1142;
  wire _10828 = _10826 ^ _10827;
  wire _10829 = _10825 ^ _10828;
  wire _10830 = _10822 ^ _10829;
  wire _10831 = r1197 ^ r1249;
  wire _10832 = r1434 ^ r1452;
  wire _10833 = _10831 ^ _10832;
  wire _10834 = r1549 ^ r1613;
  wire _10835 = r1677 ^ r1717;
  wire _10836 = _10834 ^ _10835;
  wire _10837 = _10833 ^ _10836;
  wire _10838 = r1732 ^ r1770;
  wire _10839 = r1797 ^ r1819;
  wire _10840 = _10838 ^ _10839;
  wire _10841 = r1822 ^ r1870;
  wire _10842 = r1933 ^ r1941;
  wire _10843 = _10841 ^ _10842;
  wire _10844 = _10840 ^ _10843;
  wire _10845 = _10837 ^ _10844;
  wire _10846 = _10830 ^ _10845;
  wire _10847 = r35 ^ r96;
  wire _10848 = r163 ^ r216;
  wire _10849 = _10847 ^ _10848;
  wire _10850 = r247 ^ r322;
  wire _10851 = r389 ^ r426;
  wire _10852 = _10850 ^ _10851;
  wire _10853 = _10849 ^ _10852;
  wire _10854 = r459 ^ r550;
  wire _10855 = r600 ^ r660;
  wire _10856 = _10854 ^ _10855;
  wire _10857 = r718 ^ r738;
  wire _10858 = r791 ^ r873;
  wire _10859 = _10857 ^ _10858;
  wire _10860 = _10856 ^ _10859;
  wire _10861 = _10853 ^ _10860;
  wire _10862 = r898 ^ r1002;
  wire _10863 = r1032 ^ r1100;
  wire _10864 = _10862 ^ _10863;
  wire _10865 = r1163 ^ r1203;
  wire _10866 = r1274 ^ r1281;
  wire _10867 = _10865 ^ _10866;
  wire _10868 = _10864 ^ _10867;
  wire _10869 = r1299 ^ r1368;
  wire _10870 = r1397 ^ r1563;
  wire _10871 = _10869 ^ _10870;
  wire _10872 = r1580 ^ r1640;
  wire _10873 = r1649 ^ r1804;
  wire _10874 = _10872 ^ _10873;
  wire _10875 = _10871 ^ _10874;
  wire _10876 = _10868 ^ _10875;
  wire _10877 = _10861 ^ _10876;
  wire _10878 = _10846 | _10877;
  wire _10879 = _10815 | _10878;
  wire _10880 = r34 ^ r58;
  wire _10881 = r127 ^ r178;
  wire _10882 = _10880 ^ _10881;
  wire _10883 = r245 ^ r334;
  wire _10884 = r393 ^ r460;
  wire _10885 = _10883 ^ _10884;
  wire _10886 = _10882 ^ _10885;
  wire _10887 = r545 ^ r596;
  wire _10888 = r629 ^ r670;
  wire _10889 = _10887 ^ _10888;
  wire _10890 = r730 ^ r816;
  wire _10891 = r922 ^ r957;
  wire _10892 = _10890 ^ _10891;
  wire _10893 = _10889 ^ _10892;
  wire _10894 = _10886 ^ _10893;
  wire _10895 = r1021 ^ r1112;
  wire _10896 = r1188 ^ r1339;
  wire _10897 = _10895 ^ _10896;
  wire _10898 = r1406 ^ r1489;
  wire _10899 = r1524 ^ r1606;
  wire _10900 = _10898 ^ _10899;
  wire _10901 = _10897 ^ _10900;
  wire _10902 = r1693 ^ r1765;
  wire _10903 = r1788 ^ r1828;
  wire _10904 = _10902 ^ _10903;
  wire _10905 = r1887 ^ r1974;
  wire _10906 = r1978 ^ r1982;
  wire _10907 = _10905 ^ _10906;
  wire _10908 = _10904 ^ _10907;
  wire _10909 = _10901 ^ _10908;
  wire _10910 = _10894 ^ _10909;
  wire _10911 = r33 ^ r68;
  wire _10912 = r125 ^ r204;
  wire _10913 = _10911 ^ _10912;
  wire _10914 = r258 ^ r296;
  wire _10915 = r491 ^ r551;
  wire _10916 = _10914 ^ _10915;
  wire _10917 = _10913 ^ _10916;
  wire _10918 = r614 ^ r666;
  wire _10919 = r842 ^ r928;
  wire _10920 = _10918 ^ _10919;
  wire _10921 = r968 ^ r1008;
  wire _10922 = r1092 ^ r1165;
  wire _10923 = _10921 ^ _10922;
  wire _10924 = _10920 ^ _10923;
  wire _10925 = _10917 ^ _10924;
  wire _10926 = r1190 ^ r1263;
  wire _10927 = r1313 ^ r1475;
  wire _10928 = _10926 ^ _10927;
  wire _10929 = r1496 ^ r1542;
  wire _10930 = r1577 ^ r1727;
  wire _10931 = _10929 ^ _10930;
  wire _10932 = _10928 ^ _10931;
  wire _10933 = r1767 ^ r1824;
  wire _10934 = r1864 ^ r1879;
  wire _10935 = _10933 ^ _10934;
  wire _10936 = r1943 ^ r1976;
  wire _10937 = r1977 ^ r1983;
  wire _10938 = _10936 ^ _10937;
  wire _10939 = _10935 ^ _10938;
  wire _10940 = _10932 ^ _10939;
  wire _10941 = _10925 ^ _10940;
  wire _10942 = _10910 | _10941;
  wire _10943 = r32 ^ r63;
  wire _10944 = r161 ^ r251;
  wire _10945 = _10943 ^ _10944;
  wire _10946 = r294 ^ r403;
  wire _10947 = r539 ^ r581;
  wire _10948 = _10946 ^ _10947;
  wire _10949 = _10945 ^ _10948;
  wire _10950 = r624 ^ r681;
  wire _10951 = r735 ^ r853;
  wire _10952 = _10950 ^ _10951;
  wire _10953 = r913 ^ r997;
  wire _10954 = r1024 ^ r1115;
  wire _10955 = _10953 ^ _10954;
  wire _10956 = _10952 ^ _10955;
  wire _10957 = _10949 ^ _10956;
  wire _10958 = r1214 ^ r1265;
  wire _10959 = r1284 ^ r1370;
  wire _10960 = _10958 ^ _10959;
  wire _10961 = r1455 ^ r1564;
  wire _10962 = r1598 ^ r1647;
  wire _10963 = _10961 ^ _10962;
  wire _10964 = _10960 ^ _10963;
  wire _10965 = r1711 ^ r1769;
  wire _10966 = r1773 ^ r1798;
  wire _10967 = _10965 ^ _10966;
  wire _10968 = r1815 ^ r1840;
  wire _10969 = r1853 ^ r1899;
  wire _10970 = _10968 ^ _10969;
  wire _10971 = _10967 ^ _10970;
  wire _10972 = _10964 ^ _10971;
  wire _10973 = _10957 ^ _10972;
  wire _10974 = r31 ^ r69;
  wire _10975 = r140 ^ r206;
  wire _10976 = _10974 ^ _10975;
  wire _10977 = r228 ^ r327;
  wire _10978 = r387 ^ r422;
  wire _10979 = _10977 ^ _10978;
  wire _10980 = _10976 ^ _10979;
  wire _10981 = r501 ^ r508;
  wire _10982 = r582 ^ r688;
  wire _10983 = _10981 ^ _10982;
  wire _10984 = r765 ^ r818;
  wire _10985 = r846 ^ r985;
  wire _10986 = _10984 ^ _10985;
  wire _10987 = _10983 ^ _10986;
  wire _10988 = _10980 ^ _10987;
  wire _10989 = r1043 ^ r1101;
  wire _10990 = r1162 ^ r1195;
  wire _10991 = _10989 ^ _10990;
  wire _10992 = r1235 ^ r1282;
  wire _10993 = r1305 ^ r1433;
  wire _10994 = _10992 ^ _10993;
  wire _10995 = _10991 ^ _10994;
  wire _10996 = r1535 ^ r1637;
  wire _10997 = r1678 ^ r1691;
  wire _10998 = _10996 ^ _10997;
  wire _10999 = r1799 ^ r1825;
  wire _11000 = r1841 ^ r1900;
  wire _11001 = _10999 ^ _11000;
  wire _11002 = _10998 ^ _11001;
  wire _11003 = _10995 ^ _11002;
  wire _11004 = _10988 ^ _11003;
  wire _11005 = _10973 | _11004;
  wire _11006 = _10942 | _11005;
  wire _11007 = _10879 | _11006;
  wire _11008 = r30 ^ r57;
  wire _11009 = r143 ^ r218;
  wire _11010 = _11008 ^ _11009;
  wire _11011 = r238 ^ r307;
  wire _11012 = r367 ^ r443;
  wire _11013 = _11011 ^ _11012;
  wire _11014 = _11010 ^ _11013;
  wire _11015 = r449 ^ r514;
  wire _11016 = r613 ^ r659;
  wire _11017 = _11015 ^ _11016;
  wire _11018 = r673 ^ r763;
  wire _11019 = r805 ^ r850;
  wire _11020 = _11018 ^ _11019;
  wire _11021 = _11017 ^ _11020;
  wire _11022 = _11014 ^ _11021;
  wire _11023 = r938 ^ r971;
  wire _11024 = r1053 ^ r1094;
  wire _11025 = _11023 ^ _11024;
  wire _11026 = r1129 ^ r1207;
  wire _11027 = r1272 ^ r1293;
  wire _11028 = _11026 ^ _11027;
  wire _11029 = _11025 ^ _11028;
  wire _11030 = r1351 ^ r1400;
  wire _11031 = r1451 ^ r1459;
  wire _11032 = _11030 ^ _11031;
  wire _11033 = r1470 ^ r1621;
  wire _11034 = r1675 ^ r1805;
  wire _11035 = _11033 ^ _11034;
  wire _11036 = _11032 ^ _11035;
  wire _11037 = _11029 ^ _11036;
  wire _11038 = _11022 ^ _11037;
  wire _11039 = r29 ^ r83;
  wire _11040 = r128 ^ r232;
  wire _11041 = _11039 ^ _11040;
  wire _11042 = r309 ^ r375;
  wire _11043 = r444 ^ r505;
  wire _11044 = _11042 ^ _11043;
  wire _11045 = _11041 ^ _11044;
  wire _11046 = r554 ^ r605;
  wire _11047 = r674 ^ r776;
  wire _11048 = _11046 ^ _11047;
  wire _11049 = r823 ^ r839;
  wire _11050 = r921 ^ r988;
  wire _11051 = _11049 ^ _11050;
  wire _11052 = _11048 ^ _11051;
  wire _11053 = _11045 ^ _11052;
  wire _11054 = r1048 ^ r1083;
  wire _11055 = r1135 ^ r1222;
  wire _11056 = _11054 ^ _11055;
  wire _11057 = r1228 ^ r1315;
  wire _11058 = r1359 ^ r1385;
  wire _11059 = _11057 ^ _11058;
  wire _11060 = _11056 ^ _11059;
  wire _11061 = r1423 ^ r1493;
  wire _11062 = r1737 ^ r1835;
  wire _11063 = _11061 ^ _11062;
  wire _11064 = r1966 ^ r1994;
  wire _11065 = r2004 ^ r2014;
  wire _11066 = _11064 ^ _11065;
  wire _11067 = _11063 ^ _11066;
  wire _11068 = _11060 ^ _11067;
  wire _11069 = _11053 ^ _11068;
  wire _11070 = _11038 | _11069;
  wire _11071 = r28 ^ r89;
  wire _11072 = r162 ^ r181;
  wire _11073 = _11071 ^ _11072;
  wire _11074 = r235 ^ r297;
  wire _11075 = r339 ^ r421;
  wire _11076 = _11074 ^ _11075;
  wire _11077 = _11073 ^ _11076;
  wire _11078 = r448 ^ r556;
  wire _11079 = r568 ^ r647;
  wire _11080 = _11078 ^ _11079;
  wire _11081 = r699 ^ r770;
  wire _11082 = r798 ^ r874;
  wire _11083 = _11081 ^ _11082;
  wire _11084 = _11080 ^ _11083;
  wire _11085 = _11077 ^ _11084;
  wire _11086 = r949 ^ r1054;
  wire _11087 = r1059 ^ r1098;
  wire _11088 = _11086 ^ _11087;
  wire _11089 = r1119 ^ r1189;
  wire _11090 = r1236 ^ r1307;
  wire _11091 = _11089 ^ _11090;
  wire _11092 = _11088 ^ _11091;
  wire _11093 = r1355 ^ r1457;
  wire _11094 = r1544 ^ r1616;
  wire _11095 = _11093 ^ _11094;
  wire _11096 = r1665 ^ r1746;
  wire _11097 = r1789 ^ r1874;
  wire _11098 = _11096 ^ _11097;
  wire _11099 = _11095 ^ _11098;
  wire _11100 = _11092 ^ _11099;
  wire _11101 = _11085 ^ _11100;
  wire _11102 = r27 ^ r73;
  wire _11103 = r124 ^ r199;
  wire _11104 = _11102 ^ _11103;
  wire _11105 = r225 ^ r328;
  wire _11106 = r337 ^ r412;
  wire _11107 = _11105 ^ _11106;
  wire _11108 = _11104 ^ _11107;
  wire _11109 = r499 ^ r523;
  wire _11110 = r572 ^ r625;
  wire _11111 = _11109 ^ _11110;
  wire _11112 = r680 ^ r745;
  wire _11113 = r796 ^ r858;
  wire _11114 = _11112 ^ _11113;
  wire _11115 = _11111 ^ _11114;
  wire _11116 = _11108 ^ _11115;
  wire _11117 = r939 ^ r959;
  wire _11118 = r1042 ^ r1077;
  wire _11119 = _11117 ^ _11118;
  wire _11120 = r1121 ^ r1202;
  wire _11121 = r1264 ^ r1297;
  wire _11122 = _11120 ^ _11121;
  wire _11123 = _11119 ^ _11122;
  wire _11124 = r1330 ^ r1360;
  wire _11125 = r1387 ^ r1540;
  wire _11126 = _11124 ^ _11125;
  wire _11127 = r1604 ^ r1666;
  wire _11128 = r1710 ^ r1806;
  wire _11129 = _11127 ^ _11128;
  wire _11130 = _11126 ^ _11129;
  wire _11131 = _11123 ^ _11130;
  wire _11132 = _11116 ^ _11131;
  wire _11133 = _11101 | _11132;
  wire _11134 = _11070 | _11133;
  wire _11135 = r26 ^ r75;
  wire _11136 = r152 ^ r200;
  wire _11137 = _11135 ^ _11136;
  wire _11138 = r259 ^ r293;
  wire _11139 = r373 ^ r430;
  wire _11140 = _11138 ^ _11139;
  wire _11141 = _11137 ^ _11140;
  wire _11142 = r481 ^ r507;
  wire _11143 = r616 ^ r649;
  wire _11144 = _11142 ^ _11143;
  wire _11145 = r691 ^ r755;
  wire _11146 = r809 ^ r869;
  wire _11147 = _11145 ^ _11146;
  wire _11148 = _11144 ^ _11147;
  wire _11149 = _11141 ^ _11148;
  wire _11150 = r914 ^ r954;
  wire _11151 = r1011 ^ r1074;
  wire _11152 = _11150 ^ _11151;
  wire _11153 = r1146 ^ r1176;
  wire _11154 = r1224 ^ r1312;
  wire _11155 = _11153 ^ _11154;
  wire _11156 = _11152 ^ _11155;
  wire _11157 = r1350 ^ r1490;
  wire _11158 = r1523 ^ r1584;
  wire _11159 = _11157 ^ _11158;
  wire _11160 = r1696 ^ r1752;
  wire _11161 = r1908 ^ r1918;
  wire _11162 = _11160 ^ _11161;
  wire _11163 = _11159 ^ _11162;
  wire _11164 = _11156 ^ _11163;
  wire _11165 = _11149 ^ _11164;
  wire _11166 = r25 ^ r99;
  wire _11167 = r180 ^ r244;
  wire _11168 = _11166 ^ _11167;
  wire _11169 = r319 ^ r352;
  wire _11170 = r435 ^ r487;
  wire _11171 = _11169 ^ _11170;
  wire _11172 = _11168 ^ _11171;
  wire _11173 = r571 ^ r661;
  wire _11174 = r700 ^ r802;
  wire _11175 = _11173 ^ _11174;
  wire _11176 = r880 ^ r927;
  wire _11177 = r960 ^ r1017;
  wire _11178 = _11176 ^ _11177;
  wire _11179 = _11175 ^ _11178;
  wire _11180 = _11172 ^ _11179;
  wire _11181 = r1113 ^ r1127;
  wire _11182 = r1210 ^ r1251;
  wire _11183 = _11181 ^ _11182;
  wire _11184 = r1290 ^ r1373;
  wire _11185 = r1417 ^ r1431;
  wire _11186 = _11184 ^ _11185;
  wire _11187 = _11183 ^ _11186;
  wire _11188 = r1582 ^ r1639;
  wire _11189 = r1683 ^ r1728;
  wire _11190 = _11188 ^ _11189;
  wire _11191 = r1818 ^ r1842;
  wire _11192 = r1863 ^ r1901;
  wire _11193 = _11191 ^ _11192;
  wire _11194 = _11190 ^ _11193;
  wire _11195 = _11187 ^ _11194;
  wire _11196 = _11180 ^ _11195;
  wire _11197 = _11165 | _11196;
  wire _11198 = r24 ^ r81;
  wire _11199 = r164 ^ r171;
  wire _11200 = _11198 ^ _11199;
  wire _11201 = r254 ^ r303;
  wire _11202 = r447 ^ r455;
  wire _11203 = _11201 ^ _11202;
  wire _11204 = _11200 ^ _11203;
  wire _11205 = r566 ^ r657;
  wire _11206 = r752 ^ r854;
  wire _11207 = _11205 ^ _11206;
  wire _11208 = r900 ^ r948;
  wire _11209 = r1058 ^ r1080;
  wire _11210 = _11208 ^ _11209;
  wire _11211 = _11207 ^ _11210;
  wire _11212 = _11204 ^ _11211;
  wire _11213 = r1177 ^ r1231;
  wire _11214 = r1280 ^ r1287;
  wire _11215 = _11213 ^ _11214;
  wire _11216 = r1379 ^ r1418;
  wire _11217 = r1473 ^ r1592;
  wire _11218 = _11216 ^ _11217;
  wire _11219 = _11215 ^ _11218;
  wire _11220 = r1655 ^ r1700;
  wire _11221 = r1839 ^ r1942;
  wire _11222 = _11220 ^ _11221;
  wire _11223 = r1964 ^ r1987;
  wire _11224 = r2043 ^ r2047;
  wire _11225 = _11223 ^ _11224;
  wire _11226 = _11222 ^ _11225;
  wire _11227 = _11219 ^ _11226;
  wire _11228 = _11212 ^ _11227;
  wire _11229 = r23 ^ r154;
  wire _11230 = r188 ^ r266;
  wire _11231 = _11229 ^ _11230;
  wire _11232 = r329 ^ r340;
  wire _11233 = r434 ^ r453;
  wire _11234 = _11232 ^ _11233;
  wire _11235 = _11231 ^ _11234;
  wire _11236 = r555 ^ r622;
  wire _11237 = r687 ^ r743;
  wire _11238 = _11236 ^ _11237;
  wire _11239 = r789 ^ r830;
  wire _11240 = r841 ^ r933;
  wire _11241 = _11239 ^ _11240;
  wire _11242 = _11238 ^ _11241;
  wire _11243 = _11235 ^ _11242;
  wire _11244 = r974 ^ r1004;
  wire _11245 = r1109 ^ r1147;
  wire _11246 = _11244 ^ _11245;
  wire _11247 = r1191 ^ r1253;
  wire _11248 = r1301 ^ r1395;
  wire _11249 = _11247 ^ _11248;
  wire _11250 = _11246 ^ _11249;
  wire _11251 = r1642 ^ r1658;
  wire _11252 = r1703 ^ r1869;
  wire _11253 = _11251 ^ _11252;
  wire _11254 = r1883 ^ r1996;
  wire _11255 = r2012 ^ r2027;
  wire _11256 = _11254 ^ _11255;
  wire _11257 = _11253 ^ _11256;
  wire _11258 = _11250 ^ _11257;
  wire _11259 = _11243 ^ _11258;
  wire _11260 = _11228 | _11259;
  wire _11261 = _11197 | _11260;
  wire _11262 = _11134 | _11261;
  wire _11263 = _11007 | _11262;
  wire _11264 = _10752 | _11263;
  wire _11265 = r22 ^ r100;
  wire _11266 = r141 ^ r192;
  wire _11267 = _11265 ^ _11266;
  wire _11268 = r239 ^ r321;
  wire _11269 = r374 ^ r428;
  wire _11270 = _11268 ^ _11269;
  wire _11271 = _11267 ^ _11270;
  wire _11272 = r485 ^ r513;
  wire _11273 = r609 ^ r642;
  wire _11274 = _11272 ^ _11273;
  wire _11275 = r715 ^ r723;
  wire _11276 = r783 ^ r883;
  wire _11277 = _11275 ^ _11276;
  wire _11278 = _11274 ^ _11277;
  wire _11279 = _11271 ^ _11278;
  wire _11280 = r902 ^ r1027;
  wire _11281 = r1067 ^ r1120;
  wire _11282 = _11280 ^ _11281;
  wire _11283 = r1187 ^ r1266;
  wire _11284 = r1295 ^ r1333;
  wire _11285 = _11283 ^ _11284;
  wire _11286 = _11282 ^ _11285;
  wire _11287 = r1365 ^ r1550;
  wire _11288 = r1610 ^ r1687;
  wire _11289 = _11287 ^ _11288;
  wire _11290 = r1754 ^ r1784;
  wire _11291 = r1843 ^ r1902;
  wire _11292 = _11290 ^ _11291;
  wire _11293 = _11289 ^ _11292;
  wire _11294 = _11286 ^ _11293;
  wire _11295 = _11279 ^ _11294;
  wire _11296 = r21 ^ r74;
  wire _11297 = r160 ^ r224;
  wire _11298 = _11296 ^ _11297;
  wire _11299 = r227 ^ r336;
  wire _11300 = r409 ^ r467;
  wire _11301 = _11299 ^ _11300;
  wire _11302 = _11298 ^ _11301;
  wire _11303 = r541 ^ r643;
  wire _11304 = r694 ^ r762;
  wire _11305 = _11303 ^ _11304;
  wire _11306 = r786 ^ r844;
  wire _11307 = r915 ^ r1009;
  wire _11308 = _11306 ^ _11307;
  wire _11309 = _11305 ^ _11308;
  wire _11310 = _11302 ^ _11309;
  wire _11311 = r1134 ^ r1205;
  wire _11312 = r1262 ^ r1323;
  wire _11313 = _11311 ^ _11312;
  wire _11314 = r1404 ^ r1472;
  wire _11315 = r1576 ^ r1618;
  wire _11316 = _11314 ^ _11315;
  wire _11317 = _11313 ^ _11316;
  wire _11318 = r1780 ^ r1791;
  wire _11319 = r1871 ^ r1881;
  wire _11320 = _11318 ^ _11319;
  wire _11321 = r1890 ^ r1894;
  wire _11322 = r2011 ^ r2028;
  wire _11323 = _11321 ^ _11322;
  wire _11324 = _11320 ^ _11323;
  wire _11325 = _11317 ^ _11324;
  wire _11326 = _11310 ^ _11325;
  wire _11327 = _11295 | _11326;
  wire _11328 = r20 ^ r88;
  wire _11329 = r133 ^ r191;
  wire _11330 = _11328 ^ _11329;
  wire _11331 = r326 ^ r364;
  wire _11332 = r417 ^ r470;
  wire _11333 = _11331 ^ _11332;
  wire _11334 = _11330 ^ _11333;
  wire _11335 = r576 ^ r621;
  wire _11336 = r773 ^ r864;
  wire _11337 = _11335 ^ _11336;
  wire _11338 = r912 ^ r965;
  wire _11339 = r1064 ^ r1108;
  wire _11340 = _11338 ^ _11339;
  wire _11341 = _11337 ^ _11340;
  wire _11342 = _11334 ^ _11341;
  wire _11343 = r1172 ^ r1226;
  wire _11344 = r1371 ^ r1409;
  wire _11345 = _11343 ^ _11344;
  wire _11346 = r1440 ^ r1478;
  wire _11347 = r1531 ^ r1707;
  wire _11348 = _11346 ^ _11347;
  wire _11349 = _11345 ^ _11348;
  wire _11350 = r1738 ^ r1817;
  wire _11351 = r1877 ^ r1892;
  wire _11352 = _11350 ^ _11351;
  wire _11353 = r1921 ^ r1973;
  wire _11354 = r2002 ^ r2015;
  wire _11355 = _11353 ^ _11354;
  wire _11356 = _11352 ^ _11355;
  wire _11357 = _11349 ^ _11356;
  wire _11358 = _11342 ^ _11357;
  wire _11359 = r19 ^ r59;
  wire _11360 = r130 ^ r186;
  wire _11361 = _11359 ^ _11360;
  wire _11362 = r230 ^ r300;
  wire _11363 = r349 ^ r456;
  wire _11364 = _11362 ^ _11363;
  wire _11365 = _11361 ^ _11364;
  wire _11366 = r543 ^ r667;
  wire _11367 = r675 ^ r729;
  wire _11368 = _11366 ^ _11367;
  wire _11369 = r810 ^ r871;
  wire _11370 = r930 ^ r1028;
  wire _11371 = _11369 ^ _11370;
  wire _11372 = _11368 ^ _11371;
  wire _11373 = _11365 ^ _11372;
  wire _11374 = r1106 ^ r1141;
  wire _11375 = r1173 ^ r1246;
  wire _11376 = _11374 ^ _11375;
  wire _11377 = r1327 ^ r1383;
  wire _11378 = r1482 ^ r1552;
  wire _11379 = _11377 ^ _11378;
  wire _11380 = _11376 ^ _11379;
  wire _11381 = r1557 ^ r1619;
  wire _11382 = r1681 ^ r1847;
  wire _11383 = _11381 ^ _11382;
  wire _11384 = r1990 ^ r2000;
  wire _11385 = r2001 ^ r2016;
  wire _11386 = _11384 ^ _11385;
  wire _11387 = _11383 ^ _11386;
  wire _11388 = _11380 ^ _11387;
  wire _11389 = _11373 ^ _11388;
  wire _11390 = _11358 | _11389;
  wire _11391 = _11327 | _11390;
  wire _11392 = r18 ^ r95;
  wire _11393 = r146 ^ r222;
  wire _11394 = _11392 ^ _11393;
  wire _11395 = r299 ^ r376;
  wire _11396 = r438 ^ r486;
  wire _11397 = _11395 ^ _11396;
  wire _11398 = _11394 ^ _11397;
  wire _11399 = r557 ^ r589;
  wire _11400 = r672 ^ r756;
  wire _11401 = _11399 ^ _11400;
  wire _11402 = r795 ^ r895;
  wire _11403 = r972 ^ r1088;
  wire _11404 = _11402 ^ _11403;
  wire _11405 = _11401 ^ _11404;
  wire _11406 = _11398 ^ _11405;
  wire _11407 = r1204 ^ r1247;
  wire _11408 = r1408 ^ r1464;
  wire _11409 = _11407 ^ _11408;
  wire _11410 = r1495 ^ r1504;
  wire _11411 = r1511 ^ r1528;
  wire _11412 = _11410 ^ _11411;
  wire _11413 = _11409 ^ _11412;
  wire _11414 = r1567 ^ r1609;
  wire _11415 = r1736 ^ r1794;
  wire _11416 = _11414 ^ _11415;
  wire _11417 = r1893 ^ r1931;
  wire _11418 = r2005 ^ r2006;
  wire _11419 = _11417 ^ _11418;
  wire _11420 = _11416 ^ _11419;
  wire _11421 = _11413 ^ _11420;
  wire _11422 = _11406 ^ _11421;
  wire _11423 = r17 ^ r61;
  wire _11424 = r138 ^ r176;
  wire _11425 = _11423 ^ _11424;
  wire _11426 = r256 ^ r312;
  wire _11427 = r366 ^ r415;
  wire _11428 = _11426 ^ _11427;
  wire _11429 = _11425 ^ _11428;
  wire _11430 = r452 ^ r632;
  wire _11431 = r872 ^ r896;
  wire _11432 = _11430 ^ _11431;
  wire _11433 = r984 ^ r1016;
  wire _11434 = r1073 ^ r1196;
  wire _11435 = _11433 ^ _11434;
  wire _11436 = _11432 ^ _11435;
  wire _11437 = _11429 ^ _11436;
  wire _11438 = r1225 ^ r1320;
  wire _11439 = r1364 ^ r1402;
  wire _11440 = _11438 ^ _11439;
  wire _11441 = r1444 ^ r1575;
  wire _11442 = r1593 ^ r1760;
  wire _11443 = _11441 ^ _11442;
  wire _11444 = _11440 ^ _11443;
  wire _11445 = r1792 ^ r1830;
  wire _11446 = r1876 ^ r1962;
  wire _11447 = _11445 ^ _11446;
  wire _11448 = r1975 ^ r2025;
  wire _11449 = r2032 ^ r2041;
  wire _11450 = _11448 ^ _11449;
  wire _11451 = _11447 ^ _11450;
  wire _11452 = _11444 ^ _11451;
  wire _11453 = _11437 ^ _11452;
  wire _11454 = _11422 | _11453;
  wire _11455 = r16 ^ r76;
  wire _11456 = r112 ^ r252;
  wire _11457 = _11455 ^ _11456;
  wire _11458 = r305 ^ r353;
  wire _11459 = r396 ^ r478;
  wire _11460 = _11458 ^ _11459;
  wire _11461 = _11457 ^ _11460;
  wire _11462 = r515 ^ r578;
  wire _11463 = r668 ^ r711;
  wire _11464 = _11462 ^ _11463;
  wire _11465 = r731 ^ r817;
  wire _11466 = r863 ^ r929;
  wire _11467 = _11465 ^ _11466;
  wire _11468 = _11464 ^ _11467;
  wire _11469 = _11461 ^ _11468;
  wire _11470 = r992 ^ r1044;
  wire _11471 = r1084 ^ r1118;
  wire _11472 = _11470 ^ _11471;
  wire _11473 = r1213 ^ r1273;
  wire _11474 = r1378 ^ r1447;
  wire _11475 = _11473 ^ _11474;
  wire _11476 = _11472 ^ _11475;
  wire _11477 = r1566 ^ r1581;
  wire _11478 = r1733 ^ r1812;
  wire _11479 = _11477 ^ _11478;
  wire _11480 = r1866 ^ r1932;
  wire _11481 = r1944 ^ r1959;
  wire _11482 = _11480 ^ _11481;
  wire _11483 = _11479 ^ _11482;
  wire _11484 = _11476 ^ _11483;
  wire _11485 = _11469 ^ _11484;
  wire _11486 = r15 ^ r72;
  wire _11487 = r122 ^ r195;
  wire _11488 = _11486 ^ _11487;
  wire _11489 = r257 ^ r283;
  wire _11490 = r372 ^ r399;
  wire _11491 = _11489 ^ _11490;
  wire _11492 = _11488 ^ _11491;
  wire _11493 = r464 ^ r536;
  wire _11494 = r608 ^ r631;
  wire _11495 = _11493 ^ _11494;
  wire _11496 = r712 ^ r747;
  wire _11497 = r790 ^ r886;
  wire _11498 = _11496 ^ _11497;
  wire _11499 = _11495 ^ _11498;
  wire _11500 = _11492 ^ _11499;
  wire _11501 = r964 ^ r1023;
  wire _11502 = r1093 ^ r1137;
  wire _11503 = _11501 ^ _11502;
  wire _11504 = r1216 ^ r1286;
  wire _11505 = r1352 ^ r1561;
  wire _11506 = _11504 ^ _11505;
  wire _11507 = _11503 ^ _11506;
  wire _11508 = r1591 ^ r1623;
  wire _11509 = r1685 ^ r1743;
  wire _11510 = _11508 ^ _11509;
  wire _11511 = r1771 ^ r1834;
  wire _11512 = r1920 ^ r1924;
  wire _11513 = _11511 ^ _11512;
  wire _11514 = _11510 ^ _11513;
  wire _11515 = _11507 ^ _11514;
  wire _11516 = _11500 ^ _11515;
  wire _11517 = _11485 | _11516;
  wire _11518 = _11454 | _11517;
  wire _11519 = _11391 | _11518;
  wire _11520 = r14 ^ r91;
  wire _11521 = r116 ^ r174;
  wire _11522 = _11520 ^ _11521;
  wire _11523 = r248 ^ r292;
  wire _11524 = r345 ^ r440;
  wire _11525 = _11523 ^ _11524;
  wire _11526 = _11522 ^ _11525;
  wire _11527 = r488 ^ r537;
  wire _11528 = r575 ^ r627;
  wire _11529 = _11527 ^ _11528;
  wire _11530 = r689 ^ r767;
  wire _11531 = r779 ^ r836;
  wire _11532 = _11530 ^ _11531;
  wire _11533 = _11529 ^ _11532;
  wire _11534 = _11526 ^ _11533;
  wire _11535 = r937 ^ r980;
  wire _11536 = r1046 ^ r1068;
  wire _11537 = _11535 ^ _11536;
  wire _11538 = r1159 ^ r1168;
  wire _11539 = r1239 ^ r1298;
  wire _11540 = _11538 ^ _11539;
  wire _11541 = _11537 ^ _11540;
  wire _11542 = r1414 ^ r1438;
  wire _11543 = r1519 ^ r1534;
  wire _11544 = _11542 ^ _11543;
  wire _11545 = r1599 ^ r1625;
  wire _11546 = r1698 ^ r1807;
  wire _11547 = _11545 ^ _11546;
  wire _11548 = _11544 ^ _11547;
  wire _11549 = _11541 ^ _11548;
  wire _11550 = _11534 ^ _11549;
  wire _11551 = r13 ^ r54;
  wire _11552 = r120 ^ r207;
  wire _11553 = _11551 ^ _11552;
  wire _11554 = r271 ^ r285;
  wire _11555 = r342 ^ r391;
  wire _11556 = _11554 ^ _11555;
  wire _11557 = _11553 ^ _11556;
  wire _11558 = r416 ^ r480;
  wire _11559 = r601 ^ r664;
  wire _11560 = _11558 ^ _11559;
  wire _11561 = r775 ^ r876;
  wire _11562 = r942 ^ r950;
  wire _11563 = _11561 ^ _11562;
  wire _11564 = _11560 ^ _11563;
  wire _11565 = _11557 ^ _11564;
  wire _11566 = r1005 ^ r1160;
  wire _11567 = r1215 ^ r1306;
  wire _11568 = _11566 ^ _11567;
  wire _11569 = r1354 ^ r1412;
  wire _11570 = r1468 ^ r1487;
  wire _11571 = _11569 ^ _11570;
  wire _11572 = _11568 ^ _11571;
  wire _11573 = r1506 ^ r1525;
  wire _11574 = r1645 ^ r1774;
  wire _11575 = _11573 ^ _11574;
  wire _11576 = r1811 ^ r1915;
  wire _11577 = r2007 ^ r2009;
  wire _11578 = _11576 ^ _11577;
  wire _11579 = _11575 ^ _11578;
  wire _11580 = _11572 ^ _11579;
  wire _11581 = _11565 ^ _11580;
  wire _11582 = _11550 | _11581;
  wire _11583 = r12 ^ r55;
  wire _11584 = r169 ^ r210;
  wire _11585 = _11583 ^ _11584;
  wire _11586 = r276 ^ r289;
  wire _11587 = r357 ^ r468;
  wire _11588 = _11586 ^ _11587;
  wire _11589 = _11585 ^ _11588;
  wire _11590 = r586 ^ r619;
  wire _11591 = r698 ^ r771;
  wire _11592 = _11590 ^ _11591;
  wire _11593 = r781 ^ r877;
  wire _11594 = r987 ^ r1057;
  wire _11595 = _11593 ^ _11594;
  wire _11596 = _11592 ^ _11595;
  wire _11597 = _11589 ^ _11596;
  wire _11598 = r1095 ^ r1136;
  wire _11599 = r1164 ^ r1212;
  wire _11600 = _11598 ^ _11599;
  wire _11601 = r1238 ^ r1283;
  wire _11602 = r1366 ^ r1392;
  wire _11603 = _11601 ^ _11602;
  wire _11604 = _11600 ^ _11603;
  wire _11605 = r1466 ^ r1502;
  wire _11606 = r1663 ^ r1731;
  wire _11607 = _11605 ^ _11606;
  wire _11608 = r1739 ^ r1829;
  wire _11609 = r1995 ^ r1999;
  wire _11610 = _11608 ^ _11609;
  wire _11611 = _11607 ^ _11610;
  wire _11612 = _11604 ^ _11611;
  wire _11613 = _11597 ^ _11612;
  wire _11614 = r90 ^ r147;
  wire _11615 = r197 ^ r261;
  wire _11616 = _11614 ^ _11615;
  wire _11617 = r281 ^ r407;
  wire _11618 = r522 ^ r610;
  wire _11619 = _11617 ^ _11618;
  wire _11620 = _11616 ^ _11619;
  wire _11621 = r638 ^ r703;
  wire _11622 = r848 ^ r941;
  wire _11623 = _11621 ^ _11622;
  wire _11624 = r952 ^ r1019;
  wire _11625 = r1111 ^ r1128;
  wire _11626 = _11624 ^ _11625;
  wire _11627 = _11623 ^ _11626;
  wire _11628 = _11620 ^ _11627;
  wire _11629 = r1193 ^ r1223;
  wire _11630 = r1233 ^ r1322;
  wire _11631 = _11629 ^ _11630;
  wire _11632 = r1363 ^ r1571;
  wire _11633 = r1601 ^ r1638;
  wire _11634 = _11632 ^ _11633;
  wire _11635 = _11631 ^ _11634;
  wire _11636 = r1686 ^ r1785;
  wire _11637 = r1821 ^ r1858;
  wire _11638 = _11636 ^ _11637;
  wire _11639 = r1889 ^ r1945;
  wire _11640 = r1956 ^ r1965;
  wire _11641 = _11639 ^ _11640;
  wire _11642 = _11638 ^ _11641;
  wire _11643 = _11635 ^ _11642;
  wire _11644 = _11628 ^ _11643;
  wire _11645 = _11613 | _11644;
  wire _11646 = _11582 | _11645;
  wire _11647 = r11 ^ r82;
  wire _11648 = r129 ^ r175;
  wire _11649 = _11647 ^ _11648;
  wire _11650 = r263 ^ r313;
  wire _11651 = r384 ^ r461;
  wire _11652 = _11650 ^ _11651;
  wire _11653 = _11649 ^ _11652;
  wire _11654 = r526 ^ r602;
  wire _11655 = r636 ^ r766;
  wire _11656 = _11654 ^ _11655;
  wire _11657 = r807 ^ r884;
  wire _11658 = r935 ^ r966;
  wire _11659 = _11657 ^ _11658;
  wire _11660 = _11656 ^ _11659;
  wire _11661 = _11653 ^ _11660;
  wire _11662 = r1039 ^ r1078;
  wire _11663 = r1145 ^ r1200;
  wire _11664 = _11662 ^ _11663;
  wire _11665 = r1270 ^ r1309;
  wire _11666 = r1381 ^ r1450;
  wire _11667 = _11665 ^ _11666;
  wire _11668 = _11664 ^ _11667;
  wire _11669 = r1498 ^ r1646;
  wire _11670 = r1661 ^ r1763;
  wire _11671 = _11669 ^ _11670;
  wire _11672 = r1786 ^ r1967;
  wire _11673 = r2035 ^ r2042;
  wire _11674 = _11672 ^ _11673;
  wire _11675 = _11671 ^ _11674;
  wire _11676 = _11668 ^ _11675;
  wire _11677 = _11661 ^ _11676;
  wire _11678 = r10 ^ r98;
  wire _11679 = r142 ^ r194;
  wire _11680 = _11678 ^ _11679;
  wire _11681 = r234 ^ r298;
  wire _11682 = r418 ^ r458;
  wire _11683 = _11681 ^ _11682;
  wire _11684 = _11680 ^ _11683;
  wire _11685 = r590 ^ r617;
  wire _11686 = r702 ^ r734;
  wire _11687 = _11685 ^ _11686;
  wire _11688 = r803 ^ r840;
  wire _11689 = r919 ^ r963;
  wire _11690 = _11688 ^ _11689;
  wire _11691 = _11687 ^ _11690;
  wire _11692 = _11684 ^ _11691;
  wire _11693 = r1040 ^ r1086;
  wire _11694 = r1150 ^ r1325;
  wire _11695 = _11693 ^ _11694;
  wire _11696 = r1347 ^ r1390;
  wire _11697 = r1415 ^ r1497;
  wire _11698 = _11696 ^ _11697;
  wire _11699 = _11695 ^ _11698;
  wire _11700 = r1517 ^ r1521;
  wire _11701 = r1556 ^ r1586;
  wire _11702 = _11700 ^ _11701;
  wire _11703 = r1624 ^ r1679;
  wire _11704 = r1768 ^ r1875;
  wire _11705 = _11703 ^ _11704;
  wire _11706 = _11702 ^ _11705;
  wire _11707 = _11699 ^ _11706;
  wire _11708 = _11692 ^ _11707;
  wire _11709 = _11677 | _11708;
  wire _11710 = r9 ^ r102;
  wire _11711 = r153 ^ r219;
  wire _11712 = _11710 ^ _11711;
  wire _11713 = r269 ^ r308;
  wire _11714 = r388 ^ r473;
  wire _11715 = _11713 ^ _11714;
  wire _11716 = _11712 ^ _11715;
  wire _11717 = r525 ^ r607;
  wire _11718 = r652 ^ r696;
  wire _11719 = _11717 ^ _11718;
  wire _11720 = r740 ^ r808;
  wire _11721 = r849 ^ r926;
  wire _11722 = _11720 ^ _11721;
  wire _11723 = _11719 ^ _11722;
  wire _11724 = _11716 ^ _11723;
  wire _11725 = r982 ^ r1018;
  wire _11726 = r1081 ^ r1242;
  wire _11727 = _11725 ^ _11726;
  wire _11728 = r1277 ^ r1292;
  wire _11729 = r1348 ^ r1514;
  wire _11730 = _11728 ^ _11729;
  wire _11731 = _11727 ^ _11730;
  wire _11732 = r1635 ^ r1668;
  wire _11733 = r1690 ^ r1744;
  wire _11734 = _11732 ^ _11733;
  wire _11735 = r1748 ^ r1986;
  wire _11736 = r2031 ^ r2039;
  wire _11737 = _11735 ^ _11736;
  wire _11738 = _11734 ^ _11737;
  wire _11739 = _11731 ^ _11738;
  wire _11740 = _11724 ^ _11739;
  wire _11741 = r8 ^ r110;
  wire _11742 = r123 ^ r205;
  wire _11743 = _11741 ^ _11742;
  wire _11744 = r226 ^ r320;
  wire _11745 = r333 ^ r397;
  wire _11746 = _11744 ^ _11745;
  wire _11747 = _11743 ^ _11746;
  wire _11748 = r466 ^ r520;
  wire _11749 = r678 ^ r799;
  wire _11750 = _11748 ^ _11749;
  wire _11751 = r891 ^ r945;
  wire _11752 = r1010 ^ r1087;
  wire _11753 = _11751 ^ _11752;
  wire _11754 = _11750 ^ _11753;
  wire _11755 = _11747 ^ _11754;
  wire _11756 = r1149 ^ r1241;
  wire _11757 = r1300 ^ r1380;
  wire _11758 = _11756 ^ _11757;
  wire _11759 = r1494 ^ r1589;
  wire _11760 = r1611 ^ r1694;
  wire _11761 = _11759 ^ _11760;
  wire _11762 = _11758 ^ _11761;
  wire _11763 = r1734 ^ r1735;
  wire _11764 = r1749 ^ r1800;
  wire _11765 = _11763 ^ _11764;
  wire _11766 = r1857 ^ r1919;
  wire _11767 = r1934 ^ r1950;
  wire _11768 = _11766 ^ _11767;
  wire _11769 = _11765 ^ _11768;
  wire _11770 = _11762 ^ _11769;
  wire _11771 = _11755 ^ _11770;
  wire _11772 = _11740 | _11771;
  wire _11773 = _11709 | _11772;
  wire _11774 = _11646 | _11773;
  wire _11775 = _11519 | _11774;
  wire _11776 = r7 ^ r177;
  wire _11777 = r381 ^ r414;
  wire _11778 = _11776 ^ _11777;
  wire _11779 = r496 ^ r560;
  wire _11780 = r580 ^ r639;
  wire _11781 = _11779 ^ _11780;
  wire _11782 = _11778 ^ _11781;
  wire _11783 = r685 ^ r726;
  wire _11784 = r822 ^ r889;
  wire _11785 = _11783 ^ _11784;
  wire _11786 = r946 ^ r1026;
  wire _11787 = r1143 ^ r1180;
  wire _11788 = _11786 ^ _11787;
  wire _11789 = _11785 ^ _11788;
  wire _11790 = _11782 ^ _11789;
  wire _11791 = r1296 ^ r1372;
  wire _11792 = r1467 ^ r1545;
  wire _11793 = _11791 ^ _11792;
  wire _11794 = r1641 ^ r1714;
  wire _11795 = r1787 ^ r1837;
  wire _11796 = _11794 ^ _11795;
  wire _11797 = _11793 ^ _11796;
  wire _11798 = r1859 ^ r1907;
  wire _11799 = r1916 ^ r1940;
  wire _11800 = _11798 ^ _11799;
  wire _11801 = r1952 ^ r1989;
  wire _11802 = r2040 ^ r2046;
  wire _11803 = _11801 ^ _11802;
  wire _11804 = _11800 ^ _11803;
  wire _11805 = _11797 ^ _11804;
  wire _11806 = _11790 ^ _11805;
  wire _11807 = r6 ^ r156;
  wire _11808 = r221 ^ r262;
  wire _11809 = _11807 ^ _11808;
  wire _11810 = r358 ^ r445;
  wire _11811 = r450 ^ r511;
  wire _11812 = _11810 ^ _11811;
  wire _11813 = _11809 ^ _11812;
  wire _11814 = r594 ^ r618;
  wire _11815 = r708 ^ r750;
  wire _11816 = _11814 ^ _11815;
  wire _11817 = r827 ^ r924;
  wire _11818 = r981 ^ r1030;
  wire _11819 = _11817 ^ _11818;
  wire _11820 = _11816 ^ _11819;
  wire _11821 = _11813 ^ _11820;
  wire _11822 = r1125 ^ r1166;
  wire _11823 = r1183 ^ r1255;
  wire _11824 = _11822 ^ _11823;
  wire _11825 = r1335 ^ r1422;
  wire _11826 = r1570 ^ r1585;
  wire _11827 = _11825 ^ _11826;
  wire _11828 = _11824 ^ _11827;
  wire _11829 = r1612 ^ r1670;
  wire _11830 = r1715 ^ r1917;
  wire _11831 = _11829 ^ _11830;
  wire _11832 = r1998 ^ r2008;
  wire _11833 = r2017 ^ r2030;
  wire _11834 = _11832 ^ _11833;
  wire _11835 = _11831 ^ _11834;
  wire _11836 = _11828 ^ _11835;
  wire _11837 = _11821 ^ _11836;
  wire _11838 = _11806 | _11837;
  wire _11839 = r5 ^ r114;
  wire _11840 = r208 ^ r275;
  wire _11841 = _11839 ^ _11840;
  wire _11842 = r341 ^ r442;
  wire _11843 = r500 ^ r532;
  wire _11844 = _11842 ^ _11843;
  wire _11845 = _11841 ^ _11844;
  wire _11846 = r635 ^ r706;
  wire _11847 = r732 ^ r812;
  wire _11848 = _11846 ^ _11847;
  wire _11849 = r843 ^ r905;
  wire _11850 = r973 ^ r1103;
  wire _11851 = _11849 ^ _11850;
  wire _11852 = _11848 ^ _11851;
  wire _11853 = _11845 ^ _11852;
  wire _11854 = r1110 ^ r1132;
  wire _11855 = r1257 ^ r1291;
  wire _11856 = _11854 ^ _11855;
  wire _11857 = r1393 ^ r1435;
  wire _11858 = r1505 ^ r1518;
  wire _11859 = _11857 ^ _11858;
  wire _11860 = _11856 ^ _11859;
  wire _11861 = r1603 ^ r1745;
  wire _11862 = r1757 ^ r1778;
  wire _11863 = _11861 ^ _11862;
  wire _11864 = r1826 ^ r1910;
  wire _11865 = r2033 ^ r2036;
  wire _11866 = _11864 ^ _11865;
  wire _11867 = _11863 ^ _11866;
  wire _11868 = _11860 ^ _11867;
  wire _11869 = _11853 ^ _11868;
  wire _11870 = r4 ^ r135;
  wire _11871 = r173 ^ r249;
  wire _11872 = _11870 ^ _11871;
  wire _11873 = r354 ^ r401;
  wire _11874 = r504 ^ r530;
  wire _11875 = _11873 ^ _11874;
  wire _11876 = _11872 ^ _11875;
  wire _11877 = r563 ^ r662;
  wire _11878 = r683 ^ r744;
  wire _11879 = _11877 ^ _11878;
  wire _11880 = r814 ^ r866;
  wire _11881 = r908 ^ r991;
  wire _11882 = _11880 ^ _11881;
  wire _11883 = _11879 ^ _11882;
  wire _11884 = _11876 ^ _11883;
  wire _11885 = r1029 ^ r1155;
  wire _11886 = r1167 ^ r1199;
  wire _11887 = _11885 ^ _11886;
  wire _11888 = r1243 ^ r1311;
  wire _11889 = r1386 ^ r1461;
  wire _11890 = _11888 ^ _11889;
  wire _11891 = _11887 ^ _11890;
  wire _11892 = r1536 ^ r1547;
  wire _11893 = r1622 ^ r1689;
  wire _11894 = _11892 ^ _11893;
  wire _11895 = r1766 ^ r1988;
  wire _11896 = r2038 ^ r2045;
  wire _11897 = _11895 ^ _11896;
  wire _11898 = _11894 ^ _11897;
  wire _11899 = _11891 ^ _11898;
  wire _11900 = _11884 ^ _11899;
  wire _11901 = _11869 | _11900;
  wire _11902 = _11838 | _11901;
  wire _11903 = r106 ^ r144;
  wire _11904 = r201 ^ r229;
  wire _11905 = _11903 ^ _11904;
  wire _11906 = r301 ^ r365;
  wire _11907 = r394 ^ r493;
  wire _11908 = _11906 ^ _11907;
  wire _11909 = _11905 ^ _11908;
  wire _11910 = r573 ^ r648;
  wire _11911 = r751 ^ r878;
  wire _11912 = _11910 ^ _11911;
  wire _11913 = r887 ^ r892;
  wire _11914 = r995 ^ r1090;
  wire _11915 = _11913 ^ _11914;
  wire _11916 = _11912 ^ _11915;
  wire _11917 = _11909 ^ _11916;
  wire _11918 = r1317 ^ r1337;
  wire _11919 = r1469 ^ r1516;
  wire _11920 = _11918 ^ _11919;
  wire _11921 = r1520 ^ r1595;
  wire _11922 = r1664 ^ r1772;
  wire _11923 = _11921 ^ _11922;
  wire _11924 = _11920 ^ _11923;
  wire _11925 = r1793 ^ r1937;
  wire _11926 = r1985 ^ r2010;
  wire _11927 = _11925 ^ _11926;
  wire _11928 = r2023 ^ r2024;
  wire _11929 = r2037 ^ r2044;
  wire _11930 = _11928 ^ _11929;
  wire _11931 = _11927 ^ _11930;
  wire _11932 = _11924 ^ _11931;
  wire _11933 = _11917 ^ _11932;
  wire _11934 = r3 ^ r139;
  wire _11935 = r250 ^ r310;
  wire _11936 = _11934 ^ _11935;
  wire _11937 = r335 ^ r425;
  wire _11938 = r474 ^ r546;
  wire _11939 = _11937 ^ _11938;
  wire _11940 = _11936 ^ _11939;
  wire _11941 = r567 ^ r620;
  wire _11942 = r721 ^ r725;
  wire _11943 = _11941 ^ _11942;
  wire _11944 = r820 ^ r875;
  wire _11945 = r925 ^ r1062;
  wire _11946 = _11944 ^ _11945;
  wire _11947 = _11943 ^ _11946;
  wire _11948 = _11940 ^ _11947;
  wire _11949 = r1130 ^ r1192;
  wire _11950 = r1279 ^ r1303;
  wire _11951 = _11949 ^ _11950;
  wire _11952 = r1391 ^ r1437;
  wire _11953 = r1503 ^ r1596;
  wire _11954 = _11952 ^ _11953;
  wire _11955 = _11951 ^ _11954;
  wire _11956 = r1608 ^ r1673;
  wire _11957 = r1702 ^ r1884;
  wire _11958 = _11956 ^ _11957;
  wire _11959 = r1906 ^ r1938;
  wire _11960 = r1949 ^ r1960;
  wire _11961 = _11959 ^ _11960;
  wire _11962 = _11958 ^ _11961;
  wire _11963 = _11955 ^ _11962;
  wire _11964 = _11948 ^ _11963;
  wire _11965 = _11933 | _11964;
  wire _11966 = r2 ^ r85;
  wire _11967 = r145 ^ r213;
  wire _11968 = _11966 ^ _11967;
  wire _11969 = r264 ^ r306;
  wire _11970 = r383 ^ r436;
  wire _11971 = _11969 ^ _11970;
  wire _11972 = _11968 ^ _11971;
  wire _11973 = r457 ^ r549;
  wire _11974 = r570 ^ r709;
  wire _11975 = _11973 ^ _11974;
  wire _11976 = r739 ^ r778;
  wire _11977 = r838 ^ r888;
  wire _11978 = _11976 ^ _11977;
  wire _11979 = _11975 ^ _11978;
  wire _11980 = _11972 ^ _11979;
  wire _11981 = r994 ^ r1014;
  wire _11982 = r1096 ^ r1267;
  wire _11983 = _11981 ^ _11982;
  wire _11984 = r1332 ^ r1419;
  wire _11985 = r1426 ^ r1480;
  wire _11986 = _11984 ^ _11985;
  wire _11987 = _11983 ^ _11986;
  wire _11988 = r1669 ^ r1762;
  wire _11989 = r1790 ^ r1844;
  wire _11990 = _11988 ^ _11989;
  wire _11991 = r1891 ^ r1930;
  wire _11992 = r1955 ^ r1968;
  wire _11993 = _11991 ^ _11992;
  wire _11994 = _11990 ^ _11993;
  wire _11995 = _11987 ^ _11994;
  wire _11996 = _11980 ^ _11995;
  wire _11997 = r1 ^ r64;
  wire _11998 = r134 ^ r260;
  wire _11999 = _11997 ^ _11998;
  wire _12000 = r311 ^ r368;
  wire _12001 = r429 ^ r469;
  wire _12002 = _12000 ^ _12001;
  wire _12003 = _11999 ^ _12002;
  wire _12004 = r533 ^ r615;
  wire _12005 = r684 ^ r768;
  wire _12006 = _12004 ^ _12005;
  wire _12007 = r785 ^ r860;
  wire _12008 = r916 ^ r989;
  wire _12009 = _12007 ^ _12008;
  wire _12010 = _12006 ^ _12009;
  wire _12011 = _12003 ^ _12010;
  wire _12012 = r1035 ^ r1107;
  wire _12013 = r1114 ^ r1201;
  wire _12014 = _12012 ^ _12013;
  wire _12015 = r1218 ^ r1252;
  wire _12016 = r1377 ^ r1416;
  wire _12017 = _12015 ^ _12016;
  wire _12018 = _12014 ^ _12017;
  wire _12019 = r1442 ^ r1526;
  wire _12020 = r1602 ^ r1636;
  wire _12021 = _12019 ^ _12020;
  wire _12022 = r1652 ^ r1848;
  wire _12023 = r1854 ^ r1903;
  wire _12024 = _12022 ^ _12023;
  wire _12025 = _12021 ^ _12024;
  wire _12026 = _12018 ^ _12025;
  wire _12027 = _12011 ^ _12026;
  wire _12028 = _11996 | _12027;
  wire _12029 = _11965 | _12028;
  wire _12030 = _11902 | _12029;
  wire _12031 = r0 ^ r67;
  wire _12032 = r159 ^ r278;
  wire _12033 = _12031 ^ _12032;
  wire _12034 = r386 ^ r433;
  wire _12035 = r479 ^ r510;
  wire _12036 = _12034 ^ _12035;
  wire _12037 = _12033 ^ _12036;
  wire _12038 = r595 ^ r705;
  wire _12039 = r746 ^ r813;
  wire _12040 = _12038 ^ _12039;
  wire _12041 = r861 ^ r901;
  wire _12042 = r970 ^ r1063;
  wire _12043 = _12041 ^ _12042;
  wire _12044 = _12040 ^ _12043;
  wire _12045 = _12037 ^ _12044;
  wire _12046 = r1156 ^ r1220;
  wire _12047 = r1334 ^ r1343;
  wire _12048 = _12046 ^ _12047;
  wire _12049 = r1465 ^ r1522;
  wire _12050 = r1539 ^ r1629;
  wire _12051 = _12049 ^ _12050;
  wire _12052 = _12048 ^ _12051;
  wire _12053 = r1659 ^ r1838;
  wire _12054 = r1886 ^ r1912;
  wire _12055 = _12053 ^ _12054;
  wire _12056 = r1939 ^ r1948;
  wire _12057 = r1954 ^ r1971;
  wire _12058 = _12056 ^ _12057;
  wire _12059 = _12055 ^ _12058;
  wire _12060 = _12052 ^ _12059;
  wire _12061 = _12045 ^ _12060;
  wire _12062 = r107 ^ r166;
  wire _12063 = r193 ^ r325;
  wire _12064 = _12062 ^ _12063;
  wire _12065 = r347 ^ r423;
  wire _12066 = r451 ^ r529;
  wire _12067 = _12065 ^ _12066;
  wire _12068 = _12064 ^ _12067;
  wire _12069 = r579 ^ r644;
  wire _12070 = r676 ^ r769;
  wire _12071 = _12069 ^ _12070;
  wire _12072 = r837 ^ r978;
  wire _12073 = r1013 ^ r1131;
  wire _12074 = _12072 ^ _12073;
  wire _12075 = _12071 ^ _12074;
  wire _12076 = _12068 ^ _12075;
  wire _12077 = r1181 ^ r1269;
  wire _12078 = r1321 ^ r1341;
  wire _12079 = _12077 ^ _12078;
  wire _12080 = r1424 ^ r1445;
  wire _12081 = r1481 ^ r1574;
  wire _12082 = _12080 ^ _12081;
  wire _12083 = _12079 ^ _12082;
  wire _12084 = r1644 ^ r1654;
  wire _12085 = r1697 ^ r1723;
  wire _12086 = _12084 ^ _12085;
  wire _12087 = r1758 ^ r1851;
  wire _12088 = r1861 ^ r1904;
  wire _12089 = _12087 ^ _12088;
  wire _12090 = _12086 ^ _12089;
  wire _12091 = _12083 ^ _12090;
  wire _12092 = _12076 ^ _12091;
  wire _12093 = _12061 | _12092;
  wire _12094 = r86 ^ r149;
  wire _12095 = r187 ^ r246;
  wire _12096 = _12094 ^ _12095;
  wire _12097 = r331 ^ r355;
  wire _12098 = r402 ^ r495;
  wire _12099 = _12097 ^ _12098;
  wire _12100 = _12096 ^ _12099;
  wire _12101 = r558 ^ r591;
  wire _12102 = r641 ^ r716;
  wire _12103 = _12101 ^ _12102;
  wire _12104 = r727 ^ r800;
  wire _12105 = r885 ^ r918;
  wire _12106 = _12104 ^ _12105;
  wire _12107 = _12103 ^ _12106;
  wire _12108 = _12100 ^ _12107;
  wire _12109 = r1000 ^ r1049;
  wire _12110 = r1102 ^ r1153;
  wire _12111 = _12109 ^ _12110;
  wire _12112 = r1198 ^ r1256;
  wire _12113 = r1375 ^ r1399;
  wire _12114 = _12112 ^ _12113;
  wire _12115 = _12111 ^ _12114;
  wire _12116 = r1430 ^ r1488;
  wire _12117 = r1527 ^ r1553;
  wire _12118 = _12116 ^ _12117;
  wire _12119 = r1657 ^ r1709;
  wire _12120 = r1923 ^ r1928;
  wire _12121 = _12119 ^ _12120;
  wire _12122 = _12118 ^ _12121;
  wire _12123 = _12115 ^ _12122;
  wire _12124 = _12108 ^ _12123;
  wire _12125 = r105 ^ r151;
  wire _12126 = r277 ^ r315;
  wire _12127 = _12125 ^ _12126;
  wire _12128 = r351 ^ r441;
  wire _12129 = r482 ^ r542;
  wire _12130 = _12128 ^ _12129;
  wire _12131 = _12127 ^ _12130;
  wire _12132 = r655 ^ r686;
  wire _12133 = r724 ^ r780;
  wire _12134 = _12132 ^ _12133;
  wire _12135 = r847 ^ r906;
  wire _12136 = r999 ^ r1052;
  wire _12137 = _12135 ^ _12136;
  wire _12138 = _12134 ^ _12137;
  wire _12139 = _12131 ^ _12138;
  wire _12140 = r1079 ^ r1122;
  wire _12141 = r1174 ^ r1275;
  wire _12142 = _12140 ^ _12141;
  wire _12143 = r1356 ^ r1388;
  wire _12144 = r1410 ^ r1460;
  wire _12145 = _12143 ^ _12144;
  wire _12146 = _12142 ^ _12145;
  wire _12147 = r1555 ^ r1648;
  wire _12148 = r1716 ^ r1722;
  wire _12149 = _12147 ^ _12148;
  wire _12150 = r1777 ^ r1880;
  wire _12151 = r1979 ^ r1984;
  wire _12152 = _12150 ^ _12151;
  wire _12153 = _12149 ^ _12152;
  wire _12154 = _12146 ^ _12153;
  wire _12155 = _12139 ^ _12154;
  wire _12156 = _12124 | _12155;
  wire _12157 = _12093 | _12156;
  wire _12158 = r77 ^ r118;
  wire _12159 = r182 ^ r270;
  wire _12160 = _12158 ^ _12159;
  wire _12161 = r317 ^ r356;
  wire _12162 = r398 ^ r498;
  wire _12163 = _12161 ^ _12162;
  wire _12164 = _12160 ^ _12163;
  wire _12165 = r512 ^ r574;
  wire _12166 = r650 ^ r677;
  wire _12167 = _12165 ^ _12166;
  wire _12168 = r742 ^ r801;
  wire _12169 = r852 ^ r923;
  wire _12170 = _12168 ^ _12169;
  wire _12171 = _12167 ^ _12170;
  wire _12172 = _12164 ^ _12171;
  wire _12173 = r976 ^ r1036;
  wire _12174 = r1171 ^ r1248;
  wire _12175 = _12173 ^ _12174;
  wire _12176 = r1316 ^ r1358;
  wire _12177 = r1403 ^ r1446;
  wire _12178 = _12176 ^ _12177;
  wire _12179 = _12175 ^ _12178;
  wire _12180 = r1507 ^ r1510;
  wire _12181 = r1559 ^ r1587;
  wire _12182 = _12180 ^ _12181;
  wire _12183 = r1674 ^ r1713;
  wire _12184 = r1721 ^ r1808;
  wire _12185 = _12183 ^ _12184;
  wire _12186 = _12182 ^ _12185;
  wire _12187 = _12179 ^ _12186;
  wire _12188 = _12172 ^ _12187;
  wire _12189 = r60 ^ r157;
  wire _12190 = r214 ^ r233;
  wire _12191 = _12189 ^ _12190;
  wire _12192 = r287 ^ r346;
  wire _12193 = r408 ^ r463;
  wire _12194 = _12192 ^ _12193;
  wire _12195 = _12191 ^ _12194;
  wire _12196 = r559 ^ r562;
  wire _12197 = r719 ^ r815;
  wire _12198 = _12196 ^ _12197;
  wire _12199 = r897 ^ r955;
  wire _12200 = r1133 ^ r1219;
  wire _12201 = _12199 ^ _12200;
  wire _12202 = _12198 ^ _12201;
  wire _12203 = _12195 ^ _12202;
  wire _12204 = r1245 ^ r1344;
  wire _12205 = r1407 ^ r1476;
  wire _12206 = _12204 ^ _12205;
  wire _12207 = r1501 ^ r1568;
  wire _12208 = r1643 ^ r1695;
  wire _12209 = _12207 ^ _12208;
  wire _12210 = _12206 ^ _12209;
  wire _12211 = r1719 ^ r1729;
  wire _12212 = r1751 ^ r1779;
  wire _12213 = _12211 ^ _12212;
  wire _12214 = r1781 ^ r1849;
  wire _12215 = r1855 ^ r1905;
  wire _12216 = _12214 ^ _12215;
  wire _12217 = _12213 ^ _12216;
  wire _12218 = _12210 ^ _12217;
  wire _12219 = _12203 ^ _12218;
  wire _12220 = _12188 | _12219;
  wire _12221 = r87 ^ r111;
  wire _12222 = r198 ^ r237;
  wire _12223 = _12221 ^ _12222;
  wire _12224 = r323 ^ r371;
  wire _12225 = r437 ^ r471;
  wire _12226 = _12224 ^ _12225;
  wire _12227 = _12223 ^ _12226;
  wire _12228 = r547 ^ r603;
  wire _12229 = r633 ^ r682;
  wire _12230 = _12228 ^ _12229;
  wire _12231 = r764 ^ r811;
  wire _12232 = r851 ^ r894;
  wire _12233 = _12231 ^ _12232;
  wire _12234 = _12230 ^ _12233;
  wire _12235 = _12227 ^ _12234;
  wire _12236 = r958 ^ r1033;
  wire _12237 = r1091 ^ r1124;
  wire _12238 = _12236 ^ _12237;
  wire _12239 = r1178 ^ r1260;
  wire _12240 = r1324 ^ r1331;
  wire _12241 = _12239 ^ _12240;
  wire _12242 = _12238 ^ _12241;
  wire _12243 = r1376 ^ r1396;
  wire _12244 = r1562 ^ r1588;
  wire _12245 = _12243 ^ _12244;
  wire _12246 = r1628 ^ r1708;
  wire _12247 = r1720 ^ r1809;
  wire _12248 = _12246 ^ _12247;
  wire _12249 = _12245 ^ _12248;
  wire _12250 = _12242 ^ _12249;
  wire _12251 = _12235 ^ _12250;
  wire _12252 = r52 ^ r79;
  wire _12253 = r119 ^ r209;
  wire _12254 = _12252 ^ _12253;
  wire _12255 = r279 ^ r282;
  wire _12256 = r378 ^ r424;
  wire _12257 = _12255 ^ _12256;
  wire _12258 = _12254 ^ _12257;
  wire _12259 = r509 ^ r565;
  wire _12260 = r628 ^ r713;
  wire _12261 = _12259 ^ _12260;
  wire _12262 = r741 ^ r829;
  wire _12263 = r845 ^ r910;
  wire _12264 = _12262 ^ _12263;
  wire _12265 = _12261 ^ _12264;
  wire _12266 = _12258 ^ _12265;
  wire _12267 = r1001 ^ r1003;
  wire _12268 = r1089 ^ r1209;
  wire _12269 = _12267 ^ _12268;
  wire _12270 = r1254 ^ r1294;
  wire _12271 = r1340 ^ r1513;
  wire _12272 = _12270 ^ _12271;
  wire _12273 = _12269 ^ _12272;
  wire _12274 = r1565 ^ r1597;
  wire _12275 = r1633 ^ r1680;
  wire _12276 = _12274 ^ _12275;
  wire _12277 = r1750 ^ r1775;
  wire _12278 = r1882 ^ r1914;
  wire _12279 = _12277 ^ _12278;
  wire _12280 = _12276 ^ _12279;
  wire _12281 = _12273 ^ _12280;
  wire _12282 = _12266 ^ _12281;
  wire _12283 = _12251 | _12282;
  wire _12284 = _12220 | _12283;
  wire _12285 = _12157 | _12284;
  wire _12286 = _12030 | _12285;
  wire _12287 = _11775 | _12286;
  wire _12288 = _11264 | _12287;
  wire _12289 = _10241 | _12288;
  wire _12290 = _8194 | _12289;
  wire _12291 = ~ _12290;
  wire _12292 = ~ _12291;
  wire _12293 = ~ load;
  wire _12294 = _12293 & _1;
  wire _12295 = _12292 & _12294;
  wire _12296 = _1 & _12295;
  wire _12297 = ~ _12296;
  wire _12298 = _3 & _12297;
  wire _12299 = _0 | _12298;
  wire _12300 = _12299 | _12296;
  wire [3:0] _12301 = 4'd3;
  wire [1:0] _12302 = {_0, _1726} + {_0, _3453};
  wire [1:0] _12303 = {_0, _4256} + {_0, _7485};
  wire [2:0] _12304 = {_0, _12302} + {_0, _12303};
  wire [1:0] _12305 = {_0, _9054} + {_0, _11228};
  wire [3:0] _12306 = {_0, _12304} + {_0, _0, _12305};
  wire _12307 = _12301 < _12306;
  wire _12308 = r2047 ^ _12307;
  wire _12309 = _12298 ? coded_block[2047] : r2047;
  wire _12310 = _12296 ? _12308 : _12309;
  always @ (posedge reset or posedge clock) if (reset) r2047 <= 1'd0; else if (_12300) r2047 <= _12310;
  wire [1:0] _12311 = {_0, _1726} + {_0, _3390};
  wire [1:0] _12312 = {_0, _4958} + {_0, _7132};
  wire [2:0] _12313 = {_0, _12311} + {_0, _12312};
  wire [1:0] _12314 = {_0, _8511} + {_0, _11806};
  wire [3:0] _12315 = {_0, _12313} + {_0, _0, _12314};
  wire _12316 = _12301 < _12315;
  wire _12317 = r2046 ^ _12316;
  wire _12318 = _12298 ? coded_block[2046] : r2046;
  wire _12319 = _12296 ? _12317 : _12318;
  always @ (posedge reset or posedge clock) if (reset) r2046 <= 1'd0; else if (_12300) r2046 <= _12319;
  wire [1:0] _12320 = {_0, _1533} + {_0, _3453};
  wire [1:0] _12321 = {_0, _4958} + {_0, _7262};
  wire [2:0] _12322 = {_0, _12320} + {_0, _12321};
  wire [1:0] _12323 = {_0, _10204} + {_0, _11900};
  wire [3:0] _12324 = {_0, _12322} + {_0, _0, _12323};
  wire _12325 = _12301 < _12324;
  wire _12326 = r2045 ^ _12325;
  wire _12327 = _12298 ? coded_block[2045] : r2045;
  wire _12328 = _12296 ? _12326 : _12327;
  always @ (posedge reset or posedge clock) if (reset) r2045 <= 1'd0; else if (_12300) r2045 <= _12328;
  wire [1:0] _12329 = {_0, _1533} + {_0, _3390};
  wire [1:0] _12330 = {_0, _4256} + {_0, _6589};
  wire [2:0] _12331 = {_0, _12329} + {_0, _12330};
  wire [1:0] _12332 = {_0, _10045} + {_0, _11933};
  wire [3:0] _12333 = {_0, _12331} + {_0, _0, _12332};
  wire _12334 = _12301 < _12333;
  wire _12335 = r2044 ^ _12334;
  wire _12336 = _12298 ? coded_block[2044] : r2044;
  wire _12337 = _12296 ? _12335 : _12336;
  always @ (posedge reset or posedge clock) if (reset) r2044 <= 1'd0; else if (_12300) r2044 <= _12337;
  wire [1:0] _12338 = {_0, _2044} + {_0, _2750};
  wire [1:0] _12339 = {_0, _5373} + {_0, _7357};
  wire [2:0] _12340 = {_0, _12338} + {_0, _12339};
  wire [1:0] _12341 = {_0, _8511} + {_0, _11228};
  wire [3:0] _12342 = {_0, _12340} + {_0, _0, _12341};
  wire _12343 = _12301 < _12342;
  wire _12344 = r2043 ^ _12343;
  wire _12345 = _12298 ? coded_block[2043] : r2043;
  wire _12346 = _12296 ? _12344 : _12345;
  always @ (posedge reset or posedge clock) if (reset) r2043 <= 1'd0; else if (_12300) r2043 <= _12346;
  wire [1:0] _12347 = {_0, _639} + {_0, _3517};
  wire [1:0] _12348 = {_0, _4256} + {_0, _6207};
  wire [2:0] _12349 = {_0, _12347} + {_0, _12348};
  wire [1:0] _12350 = {_0, _8767} + {_0, _11677};
  wire [3:0] _12351 = {_0, _12349} + {_0, _0, _12350};
  wire _12352 = _12301 < _12351;
  wire _12353 = r2042 ^ _12352;
  wire _12354 = _12298 ? coded_block[2042] : r2042;
  wire _12355 = _12296 ? _12353 : _12354;
  always @ (posedge reset or posedge clock) if (reset) r2042 <= 1'd0; else if (_12300) r2042 <= _12355;
  wire [1:0] _12356 = {_0, _639} + {_0, _3167};
  wire [1:0] _12357 = {_0, _4861} + {_0, _7132};
  wire [2:0] _12358 = {_0, _12356} + {_0, _12357};
  wire [1:0] _12359 = {_0, _9054} + {_0, _11453};
  wire [3:0] _12360 = {_0, _12358} + {_0, _0, _12359};
  wire _12361 = _12301 < _12360;
  wire _12362 = r2041 ^ _12361;
  wire _12363 = _12298 ? coded_block[2041] : r2041;
  wire _12364 = _12296 ? _12362 : _12363;
  always @ (posedge reset or posedge clock) if (reset) r2041 <= 1'd0; else if (_12300) r2041 <= _12364;
  wire [1:0] _12365 = {_0, _2044} + {_0, _2847};
  wire [1:0] _12366 = {_0, _6108} + {_0, _6207};
  wire [2:0] _12367 = {_0, _12365} + {_0, _12366};
  wire [1:0] _12368 = {_0, _9054} + {_0, _11806};
  wire [3:0] _12369 = {_0, _12367} + {_0, _0, _12368};
  wire _12370 = _12301 < _12369;
  wire _12371 = r2040 ^ _12370;
  wire _12372 = _12298 ? coded_block[2040] : r2040;
  wire _12373 = _12296 ? _12371 : _12372;
  always @ (posedge reset or posedge clock) if (reset) r2040 <= 1'd0; else if (_12300) r2040 <= _12373;
  wire [1:0] _12374 = {_0, _2044} + {_0, _2302};
  wire [1:0] _12375 = {_0, _4703} + {_0, _7485};
  wire [2:0] _12376 = {_0, _12374} + {_0, _12375};
  wire [1:0] _12377 = {_0, _10141} + {_0, _11740};
  wire [3:0] _12378 = {_0, _12376} + {_0, _0, _12377};
  wire _12379 = _12301 < _12378;
  wire _12380 = r2039 ^ _12379;
  wire _12381 = _12298 ? coded_block[2039] : r2039;
  wire _12382 = _12296 ? _12380 : _12381;
  always @ (posedge reset or posedge clock) if (reset) r2039 <= 1'd0; else if (_12300) r2039 <= _12382;
  wire [1:0] _12383 = {_0, _289} + {_0, _2750};
  wire [1:0] _12384 = {_0, _6108} + {_0, _7837};
  wire [2:0] _12385 = {_0, _12383} + {_0, _12384};
  wire [1:0] _12386 = {_0, _10045} + {_0, _11900};
  wire [3:0] _12387 = {_0, _12385} + {_0, _0, _12386};
  wire _12388 = _12301 < _12387;
  wire _12389 = r2038 ^ _12388;
  wire _12390 = _12298 ? coded_block[2038] : r2038;
  wire _12391 = _12296 ? _12389 : _12390;
  always @ (posedge reset or posedge clock) if (reset) r2038 <= 1'd0; else if (_12300) r2038 <= _12391;
  wire [1:0] _12392 = {_0, _289} + {_0, _2847};
  wire [1:0] _12393 = {_0, _5373} + {_0, _6845};
  wire [2:0] _12394 = {_0, _12392} + {_0, _12393};
  wire [1:0] _12395 = {_0, _10204} + {_0, _11933};
  wire [3:0] _12396 = {_0, _12394} + {_0, _0, _12395};
  wire _12397 = _12301 < _12396;
  wire _12398 = r2037 ^ _12397;
  wire _12399 = _12298 ? coded_block[2037] : r2037;
  wire _12400 = _12296 ? _12398 : _12399;
  always @ (posedge reset or posedge clock) if (reset) r2037 <= 1'd0; else if (_12300) r2037 <= _12400;
  wire [1:0] _12401 = {_0, _545} + {_0, _3167};
  wire [1:0] _12402 = {_0, _5949} + {_0, _6589};
  wire [2:0] _12403 = {_0, _12401} + {_0, _12402};
  wire [1:0] _12404 = {_0, _10204} + {_0, _11869};
  wire [3:0] _12405 = {_0, _12403} + {_0, _0, _12404};
  wire _12406 = _12301 < _12405;
  wire _12407 = r2036 ^ _12406;
  wire _12408 = _12298 ? coded_block[2036] : r2036;
  wire _12409 = _12296 ? _12407 : _12408;
  always @ (posedge reset or posedge clock) if (reset) r2036 <= 1'd0; else if (_12300) r2036 <= _12409;
  wire [1:0] _12410 = {_0, _735} + {_0, _3742};
  wire [1:0] _12411 = {_0, _5373} + {_0, _7132};
  wire [2:0] _12412 = {_0, _12410} + {_0, _12411};
  wire [1:0] _12413 = {_0, _10141} + {_0, _11677};
  wire [3:0] _12414 = {_0, _12412} + {_0, _0, _12413};
  wire _12415 = _12301 < _12414;
  wire _12416 = r2035 ^ _12415;
  wire _12417 = _12298 ? coded_block[2035] : r2035;
  wire _12418 = _12296 ? _12416 : _12417;
  always @ (posedge reset or posedge clock) if (reset) r2035 <= 1'd0; else if (_12300) r2035 <= _12418;
  wire [1:0] _12419 = {_0, _545} + {_0, _2941};
  wire [1:0] _12420 = {_0, _4861} + {_0, _7262};
  wire [2:0] _12421 = {_0, _12419} + {_0, _12420};
  wire [1:0] _12422 = {_0, _10045} + {_0, _10685};
  wire [3:0] _12423 = {_0, _12421} + {_0, _0, _12422};
  wire _12424 = _12301 < _12423;
  wire _12425 = r2034 ^ _12424;
  wire _12426 = _12298 ? coded_block[2034] : r2034;
  wire _12427 = _12296 ? _12425 : _12426;
  always @ (posedge reset or posedge clock) if (reset) r2034 <= 1'd0; else if (_12300) r2034 <= _12427;
  wire [1:0] _12428 = {_0, _1533} + {_0, _2878};
  wire [1:0] _12429 = {_0, _5534} + {_0, _7132};
  wire [2:0] _12430 = {_0, _12428} + {_0, _12429};
  wire [1:0] _12431 = {_0, _8799} + {_0, _11869};
  wire [3:0] _12432 = {_0, _12430} + {_0, _0, _12431};
  wire _12433 = _12301 < _12432;
  wire _12434 = r2033 ^ _12433;
  wire _12435 = _12298 ? coded_block[2033] : r2033;
  wire _12436 = _12296 ? _12434 : _12435;
  always @ (posedge reset or posedge clock) if (reset) r2033 <= 1'd0; else if (_12300) r2033 <= _12436;
  wire [1:0] _12437 = {_0, _735} + {_0, _2557};
  wire [1:0] _12438 = {_0, _4703} + {_0, _6207};
  wire [2:0] _12439 = {_0, _12437} + {_0, _12438};
  wire [1:0] _12440 = {_0, _8511} + {_0, _11453};
  wire [3:0] _12441 = {_0, _12439} + {_0, _0, _12440};
  wire _12442 = _12301 < _12441;
  wire _12443 = r2032 ^ _12442;
  wire _12444 = _12298 ? coded_block[2032] : r2032;
  wire _12445 = _12296 ? _12443 : _12444;
  always @ (posedge reset or posedge clock) if (reset) r2032 <= 1'd0; else if (_12300) r2032 <= _12445;
  wire [1:0] _12446 = {_0, _1726} + {_0, _2494};
  wire [1:0] _12447 = {_0, _4861} + {_0, _7357};
  wire [2:0] _12448 = {_0, _12446} + {_0, _12447};
  wire [1:0] _12449 = {_0, _8767} + {_0, _11740};
  wire [3:0] _12450 = {_0, _12448} + {_0, _0, _12449};
  wire _12451 = _12301 < _12450;
  wire _12452 = r2031 ^ _12451;
  wire _12453 = _12298 ? coded_block[2031] : r2031;
  wire _12454 = _12296 ? _12452 : _12453;
  always @ (posedge reset or posedge clock) if (reset) r2031 <= 1'd0; else if (_12300) r2031 <= _12454;
  wire [1:0] _12455 = {_0, _1184} + {_0, _2302};
  wire [1:0] _12456 = {_0, _5373} + {_0, _7837};
  wire [2:0] _12457 = {_0, _12455} + {_0, _12456};
  wire [1:0] _12458 = {_0, _8352} + {_0, _11837};
  wire [3:0] _12459 = {_0, _12457} + {_0, _0, _12458};
  wire _12460 = _12301 < _12459;
  wire _12461 = r2030 ^ _12460;
  wire _12462 = _12298 ? coded_block[2030] : r2030;
  wire _12463 = _12296 ? _12461 : _12462;
  always @ (posedge reset or posedge clock) if (reset) r2030 <= 1'd0; else if (_12300) r2030 <= _12463;
  wire [1:0] _12464 = {_0, _1057} + {_0, _3517};
  wire [1:0] _12465 = {_0, _4861} + {_0, _6589};
  wire [2:0] _12466 = {_0, _12464} + {_0, _12465};
  wire [1:0] _12467 = {_0, _8799} + {_0, _10654};
  wire [3:0] _12468 = {_0, _12466} + {_0, _0, _12467};
  wire _12469 = _12301 < _12468;
  wire _12470 = r2029 ^ _12469;
  wire _12471 = _12298 ? coded_block[2029] : r2029;
  wire _12472 = _12296 ? _12470 : _12471;
  always @ (posedge reset or posedge clock) if (reset) r2029 <= 1'd0; else if (_12300) r2029 <= _12472;
  wire [1:0] _12473 = {_0, _639} + {_0, _2941};
  wire [1:0] _12474 = {_0, _5949} + {_0, _7485};
  wire [2:0] _12475 = {_0, _12473} + {_0, _12474};
  wire [1:0] _12476 = {_0, _8511} + {_0, _11326};
  wire [3:0] _12477 = {_0, _12475} + {_0, _0, _12476};
  wire _12478 = _12301 < _12477;
  wire _12479 = r2028 ^ _12478;
  wire _12480 = _12298 ? coded_block[2028] : r2028;
  wire _12481 = _12296 ? _12479 : _12480;
  always @ (posedge reset or posedge clock) if (reset) r2028 <= 1'd0; else if (_12300) r2028 <= _12481;
  wire [1:0] _12482 = {_0, _1057} + {_0, _3294};
  wire [1:0] _12483 = {_0, _5534} + {_0, _6207};
  wire [2:0] _12484 = {_0, _12482} + {_0, _12483};
  wire [1:0] _12485 = {_0, _10014} + {_0, _11259};
  wire [3:0] _12486 = {_0, _12484} + {_0, _0, _12485};
  wire _12487 = _12301 < _12486;
  wire _12488 = r2027 ^ _12487;
  wire _12489 = _12298 ? coded_block[2027] : r2027;
  wire _12490 = _12296 ? _12488 : _12489;
  always @ (posedge reset or posedge clock) if (reset) r2027 <= 1'd0; else if (_12300) r2027 <= _12490;
  wire [1:0] _12491 = {_0, _1695} + {_0, _2557};
  wire [1:0] _12492 = {_0, _5310} + {_0, _7262};
  wire [2:0] _12493 = {_0, _12491} + {_0, _12492};
  wire [1:0] _12494 = {_0, _9822} + {_0, _10717};
  wire [3:0] _12495 = {_0, _12493} + {_0, _0, _12494};
  wire _12496 = _12301 < _12495;
  wire _12497 = r2026 ^ _12496;
  wire _12498 = _12298 ? coded_block[2026] : r2026;
  wire _12499 = _12296 ? _12497 : _12498;
  always @ (posedge reset or posedge clock) if (reset) r2026 <= 1'd0; else if (_12300) r2026 <= _12499;
  wire [1:0] _12500 = {_0, _1726} + {_0, _2878};
  wire [1:0] _12501 = {_0, _5470} + {_0, _6589};
  wire [2:0] _12502 = {_0, _12500} + {_0, _12501};
  wire [1:0] _12503 = {_0, _8957} + {_0, _11453};
  wire [3:0] _12504 = {_0, _12502} + {_0, _0, _12503};
  wire _12505 = _12301 < _12504;
  wire _12506 = r2025 ^ _12505;
  wire _12507 = _12298 ? coded_block[2025] : r2025;
  wire _12508 = _12296 ? _12506 : _12507;
  always @ (posedge reset or posedge clock) if (reset) r2025 <= 1'd0; else if (_12300) r2025 <= _12508;
  wire [1:0] _12509 = {_0, _1695} + {_0, _3742};
  wire [1:0] _12510 = {_0, _5790} + {_0, _7837};
  wire [2:0] _12511 = {_0, _12509} + {_0, _12510};
  wire [1:0] _12512 = {_0, _9886} + {_0, _11933};
  wire [3:0] _12513 = {_0, _12511} + {_0, _0, _12512};
  wire _12514 = _12301 < _12513;
  wire _12515 = r2024 ^ _12514;
  wire _12516 = _12298 ? coded_block[2024] : r2024;
  wire _12517 = _12296 ? _12515 : _12516;
  always @ (posedge reset or posedge clock) if (reset) r2024 <= 1'd0; else if (_12300) r2024 <= _12517;
  wire [1:0] _12518 = {_0, _545} + {_0, _3294};
  wire [1:0] _12519 = {_0, _4319} + {_0, _7132};
  wire [2:0] _12520 = {_0, _12518} + {_0, _12519};
  wire [1:0] _12521 = {_0, _8352} + {_0, _11933};
  wire [3:0] _12522 = {_0, _12520} + {_0, _0, _12521};
  wire _12523 = _12301 < _12522;
  wire _12524 = r2023 ^ _12523;
  wire _12525 = _12298 ? coded_block[2023] : r2023;
  wire _12526 = _12296 ? _12524 : _12525;
  always @ (posedge reset or posedge clock) if (reset) r2023 <= 1'd0; else if (_12300) r2023 <= _12526;
  wire [1:0] _12527 = {_0, _1184} + {_0, _2592};
  wire [1:0] _12528 = {_0, _5022} + {_0, _6207};
  wire [2:0] _12529 = {_0, _12527} + {_0, _12528};
  wire [1:0] _12530 = {_0, _10045} + {_0, _10654};
  wire [3:0] _12531 = {_0, _12529} + {_0, _0, _12530};
  wire _12532 = _12301 < _12531;
  wire _12533 = r2022 ^ _12532;
  wire _12534 = _12298 ? coded_block[2022] : r2022;
  wire _12535 = _12296 ? _12533 : _12534;
  always @ (posedge reset or posedge clock) if (reset) r2022 <= 1'd0; else if (_12300) r2022 <= _12535;
  wire [1:0] _12536 = {_0, _1533} + {_0, _2239};
  wire [1:0] _12537 = {_0, _4861} + {_0, _6845};
  wire [2:0] _12538 = {_0, _12536} + {_0, _12537};
  wire [1:0] _12539 = {_0, _10014} + {_0, _10717};
  wire [3:0] _12540 = {_0, _12538} + {_0, _0, _12539};
  wire _12541 = _12301 < _12540;
  wire _12542 = r2021 ^ _12541;
  wire _12543 = _12298 ? coded_block[2021] : r2021;
  wire _12544 = _12296 ? _12542 : _12543;
  always @ (posedge reset or posedge clock) if (reset) r2021 <= 1'd0; else if (_12300) r2021 <= _12544;
  wire [1:0] _12545 = {_0, _1533} + {_0, _2175};
  wire [1:0] _12546 = {_0, _5470} + {_0, _7485};
  wire [2:0] _12547 = {_0, _12545} + {_0, _12546};
  wire [1:0] _12548 = {_0, _8352} + {_0, _10685};
  wire [3:0] _12549 = {_0, _12547} + {_0, _0, _12548};
  wire _12550 = _12301 < _12549;
  wire _12551 = r2020 ^ _12550;
  wire _12552 = _12298 ? coded_block[2020] : r2020;
  wire _12553 = _12296 ? _12551 : _12552;
  always @ (posedge reset or posedge clock) if (reset) r2020 <= 1'd0; else if (_12300) r2020 <= _12553;
  wire [1:0] _12554 = {_0, _289} + {_0, _2144};
  wire [1:0] _12555 = {_0, _5022} + {_0, _7357};
  wire [2:0] _12556 = {_0, _12554} + {_0, _12555};
  wire [1:0] _12557 = {_0, _8799} + {_0, _10685};
  wire [3:0] _12558 = {_0, _12556} + {_0, _0, _12557};
  wire _12559 = _12301 < _12558;
  wire _12560 = r2019 ^ _12559;
  wire _12561 = _12298 ? coded_block[2019] : r2019;
  wire _12562 = _12296 ? _12560 : _12561;
  always @ (posedge reset or posedge clock) if (reset) r2019 <= 1'd0; else if (_12300) r2019 <= _12562;
  wire [1:0] _12563 = {_0, _2013} + {_0, _2302};
  wire [1:0] _12564 = {_0, _5310} + {_0, _6845};
  wire [2:0] _12565 = {_0, _12563} + {_0, _12564};
  wire [1:0] _12566 = {_0, _9886} + {_0, _10685};
  wire [3:0] _12567 = {_0, _12565} + {_0, _0, _12566};
  wire _12568 = _12301 < _12567;
  wire _12569 = r2018 ^ _12568;
  wire _12570 = _12298 ? coded_block[2018] : r2018;
  wire _12571 = _12296 ? _12569 : _12570;
  always @ (posedge reset or posedge clock) if (reset) r2018 <= 1'd0; else if (_12300) r2018 <= _12571;
  wire [1:0] _12572 = {_0, _1917} + {_0, _2494};
  wire [1:0] _12573 = {_0, _4256} + {_0, _7262};
  wire [2:0] _12574 = {_0, _12572} + {_0, _12573};
  wire [1:0] _12575 = {_0, _8799} + {_0, _11837};
  wire [3:0] _12576 = {_0, _12574} + {_0, _0, _12575};
  wire _12577 = _12301 < _12576;
  wire _12578 = r2017 ^ _12577;
  wire _12579 = _12298 ? coded_block[2017] : r2017;
  wire _12580 = _12296 ? _12578 : _12579;
  always @ (posedge reset or posedge clock) if (reset) r2017 <= 1'd0; else if (_12300) r2017 <= _12580;
  wire [1:0] _12581 = {_0, _2013} + {_0, _2750};
  wire [1:0] _12582 = {_0, _5790} + {_0, _6589};
  wire [2:0] _12583 = {_0, _12581} + {_0, _12582};
  wire [1:0] _12584 = {_0, _9822} + {_0, _11389};
  wire [3:0] _12585 = {_0, _12583} + {_0, _0, _12584};
  wire _12586 = _12301 < _12585;
  wire _12587 = r2016 ^ _12586;
  wire _12588 = _12298 ? coded_block[2016] : r2016;
  wire _12589 = _12296 ? _12587 : _12588;
  always @ (posedge reset or posedge clock) if (reset) r2016 <= 1'd0; else if (_12300) r2016 <= _12589;
  wire [1:0] _12590 = {_0, _1917} + {_0, _2239};
  wire [1:0] _12591 = {_0, _4958} + {_0, _6589};
  wire [2:0] _12592 = {_0, _12590} + {_0, _12591};
  wire [1:0] _12593 = {_0, _8352} + {_0, _11358};
  wire [3:0] _12594 = {_0, _12592} + {_0, _0, _12593};
  wire _12595 = _12301 < _12594;
  wire _12596 = r2015 ^ _12595;
  wire _12597 = _12298 ? coded_block[2015] : r2015;
  wire _12598 = _12296 ? _12596 : _12597;
  always @ (posedge reset or posedge clock) if (reset) r2015 <= 1'd0; else if (_12300) r2015 <= _12598;
  wire [1:0] _12599 = {_0, _352} + {_0, _2175};
  wire [1:0] _12600 = {_0, _4319} + {_0, _7837};
  wire [2:0] _12601 = {_0, _12599} + {_0, _12600};
  wire [1:0] _12602 = {_0, _10141} + {_0, _11069};
  wire [3:0] _12603 = {_0, _12601} + {_0, _0, _12602};
  wire _12604 = _12301 < _12603;
  wire _12605 = r2014 ^ _12604;
  wire _12606 = _12298 ? coded_block[2014] : r2014;
  wire _12607 = _12296 ? _12605 : _12606;
  always @ (posedge reset or posedge clock) if (reset) r2014 <= 1'd0; else if (_12300) r2014 <= _12607;
  wire [1:0] _12608 = {_0, _352} + {_0, _2494};
  wire [1:0] _12609 = {_0, _4958} + {_0, _7485};
  wire [2:0] _12610 = {_0, _12608} + {_0, _12609};
  wire [1:0] _12611 = {_0, _8957} + {_0, _10303};
  wire [3:0] _12612 = {_0, _12610} + {_0, _0, _12611};
  wire _12613 = _12301 < _12612;
  wire _12614 = r2013 ^ _12613;
  wire _12615 = _12298 ? coded_block[2013] : r2013;
  wire _12616 = _12296 ? _12614 : _12615;
  always @ (posedge reset or posedge clock) if (reset) r2013 <= 1'd0; else if (_12300) r2013 <= _12616;
  wire [1:0] _12617 = {_0, _1917} + {_0, _3390};
  wire [1:0] _12618 = {_0, _5949} + {_0, _6845};
  wire [2:0] _12619 = {_0, _12617} + {_0, _12618};
  wire [1:0] _12620 = {_0, _10172} + {_0, _11259};
  wire [3:0] _12621 = {_0, _12619} + {_0, _0, _12620};
  wire _12622 = _12301 < _12621;
  wire _12623 = r2012 ^ _12622;
  wire _12624 = _12298 ? coded_block[2012] : r2012;
  wire _12625 = _12296 ? _12623 : _12624;
  always @ (posedge reset or posedge clock) if (reset) r2012 <= 1'd0; else if (_12300) r2012 <= _12625;
  wire [1:0] _12626 = {_0, _2044} + {_0, _2144};
  wire [1:0] _12627 = {_0, _5246} + {_0, _7837};
  wire [2:0] _12628 = {_0, _12626} + {_0, _12627};
  wire [1:0] _12629 = {_0, _8957} + {_0, _11326};
  wire [3:0] _12630 = {_0, _12628} + {_0, _0, _12629};
  wire _12631 = _12301 < _12630;
  wire _12632 = r2011 ^ _12631;
  wire _12633 = _12298 ? coded_block[2011] : r2011;
  wire _12634 = _12296 ? _12632 : _12633;
  always @ (posedge reset or posedge clock) if (reset) r2011 <= 1'd0; else if (_12300) r2011 <= _12634;
  wire [1:0] _12635 = {_0, _2013} + {_0, _2592};
  wire [1:0] _12636 = {_0, _4350} + {_0, _7357};
  wire [2:0] _12637 = {_0, _12635} + {_0, _12636};
  wire [1:0] _12638 = {_0, _8894} + {_0, _11933};
  wire [3:0] _12639 = {_0, _12637} + {_0, _0, _12638};
  wire _12640 = _12301 < _12639;
  wire _12641 = r2010 ^ _12640;
  wire _12642 = _12298 ? coded_block[2010] : r2010;
  wire _12643 = _12296 ? _12641 : _12642;
  always @ (posedge reset or posedge clock) if (reset) r2010 <= 1'd0; else if (_12300) r2010 <= _12643;
  wire [1:0] _12644 = {_0, _352} + {_0, _3870};
  wire [1:0] _12645 = {_0, _5534} + {_0, _6589};
  wire [2:0] _12646 = {_0, _12644} + {_0, _12645};
  wire [1:0] _12647 = {_0, _9054} + {_0, _11581};
  wire [3:0] _12648 = {_0, _12646} + {_0, _0, _12647};
  wire _12649 = _12301 < _12648;
  wire _12650 = r2009 ^ _12649;
  wire _12651 = _12298 ? coded_block[2009] : r2009;
  wire _12652 = _12296 ? _12650 : _12651;
  always @ (posedge reset or posedge clock) if (reset) r2009 <= 1'd0; else if (_12300) r2009 <= _12652;
  wire [1:0] _12653 = {_0, _1057} + {_0, _2336};
  wire [1:0] _12654 = {_0, _4319} + {_0, _7485};
  wire [2:0] _12655 = {_0, _12653} + {_0, _12654};
  wire [1:0] _12656 = {_0, _10204} + {_0, _11837};
  wire [3:0] _12657 = {_0, _12655} + {_0, _0, _12656};
  wire _12658 = _12301 < _12657;
  wire _12659 = r2008 ^ _12658;
  wire _12660 = _12298 ? coded_block[2008] : r2008;
  wire _12661 = _12296 ? _12659 : _12660;
  always @ (posedge reset or posedge clock) if (reset) r2008 <= 1'd0; else if (_12300) r2008 <= _12661;
  wire [1:0] _12662 = {_0, _97} + {_0, _3517};
  wire [1:0] _12663 = {_0, _5949} + {_0, _7132};
  wire [2:0] _12664 = {_0, _12662} + {_0, _12663};
  wire [1:0] _12665 = {_0, _8957} + {_0, _11581};
  wire [3:0] _12666 = {_0, _12664} + {_0, _0, _12665};
  wire _12667 = _12301 < _12666;
  wire _12668 = r2007 ^ _12667;
  wire _12669 = _12298 ? coded_block[2007] : r2007;
  wire _12670 = _12296 ? _12668 : _12669;
  always @ (posedge reset or posedge clock) if (reset) r2007 <= 1'd0; else if (_12300) r2007 <= _12670;
  wire [1:0] _12671 = {_0, _545} + {_0, _3870};
  wire [1:0] _12672 = {_0, _5246} + {_0, _6525};
  wire [2:0] _12673 = {_0, _12671} + {_0, _12672};
  wire [1:0] _12674 = {_0, _8543} + {_0, _11422};
  wire [3:0] _12675 = {_0, _12673} + {_0, _0, _12674};
  wire _12676 = _12301 < _12675;
  wire _12677 = r2006 ^ _12676;
  wire _12678 = _12298 ? coded_block[2006] : r2006;
  wire _12679 = _12296 ? _12677 : _12678;
  always @ (posedge reset or posedge clock) if (reset) r2006 <= 1'd0; else if (_12300) r2006 <= _12679;
  wire [1:0] _12680 = {_0, _1568} + {_0, _2813};
  wire [1:0] _12681 = {_0, _4350} + {_0, _7389};
  wire [2:0] _12682 = {_0, _12680} + {_0, _12681};
  wire [1:0] _12683 = {_0, _10204} + {_0, _11422};
  wire [3:0] _12684 = {_0, _12682} + {_0, _0, _12683};
  wire _12685 = _12301 < _12684;
  wire _12686 = r2005 ^ _12685;
  wire _12687 = _12298 ? coded_block[2005] : r2005;
  wire _12688 = _12296 ? _12686 : _12687;
  always @ (posedge reset or posedge clock) if (reset) r2005 <= 1'd0; else if (_12300) r2005 <= _12688;
  wire [1:0] _12689 = {_0, _1568} + {_0, _3294};
  wire [1:0] _12690 = {_0, _6108} + {_0, _7326};
  wire [2:0] _12691 = {_0, _12689} + {_0, _12690};
  wire [1:0] _12692 = {_0, _8894} + {_0, _11069};
  wire [3:0] _12693 = {_0, _12691} + {_0, _0, _12692};
  wire _12694 = _12301 < _12693;
  wire _12695 = r2004 ^ _12694;
  wire _12696 = _12298 ? coded_block[2004] : r2004;
  wire _12697 = _12296 ? _12695 : _12696;
  always @ (posedge reset or posedge clock) if (reset) r2004 <= 1'd0; else if (_12300) r2004 <= _12697;
  wire [1:0] _12698 = {_0, _97} + {_0, _2336};
  wire [1:0] _12699 = {_0, _4574} + {_0, _7262};
  wire [2:0] _12700 = {_0, _12698} + {_0, _12699};
  wire [1:0] _12701 = {_0, _9054} + {_0, _10303};
  wire [3:0] _12702 = {_0, _12700} + {_0, _0, _12701};
  wire _12703 = _12301 < _12702;
  wire _12704 = r2003 ^ _12703;
  wire _12705 = _12298 ? coded_block[2003] : r2003;
  wire _12706 = _12296 ? _12704 : _12705;
  always @ (posedge reset or posedge clock) if (reset) r2003 <= 1'd0; else if (_12300) r2003 <= _12706;
  wire [1:0] _12707 = {_0, _1184} + {_0, _3262};
  wire [1:0] _12708 = {_0, _6108} + {_0, _6845};
  wire [2:0] _12709 = {_0, _12707} + {_0, _12708};
  wire [1:0] _12710 = {_0, _8799} + {_0, _11358};
  wire [3:0] _12711 = {_0, _12709} + {_0, _0, _12710};
  wire _12712 = _12301 < _12711;
  wire _12713 = r2002 ^ _12712;
  wire _12714 = _12298 ? coded_block[2002] : r2002;
  wire _12715 = _12296 ? _12713 : _12714;
  always @ (posedge reset or posedge clock) if (reset) r2002 <= 1'd0; else if (_12300) r2002 <= _12715;
  wire [1:0] _12716 = {_0, _1533} + {_0, _2782};
  wire [1:0] _12717 = {_0, _4319} + {_0, _7357};
  wire [2:0] _12718 = {_0, _12716} + {_0, _12717};
  wire [1:0] _12719 = {_0, _10172} + {_0, _11389};
  wire [3:0] _12720 = {_0, _12718} + {_0, _0, _12719};
  wire _12721 = _12301 < _12720;
  wire _12722 = r2001 ^ _12721;
  wire _12723 = _12298 ? coded_block[2001] : r2001;
  wire _12724 = _12296 ? _12722 : _12723;
  always @ (posedge reset or posedge clock) if (reset) r2001 <= 1'd0; else if (_12300) r2001 <= _12724;
  wire [1:0] _12725 = {_0, _1662} + {_0, _2813};
  wire [1:0] _12726 = {_0, _5407} + {_0, _6525};
  wire [2:0] _12727 = {_0, _12725} + {_0, _12726};
  wire [1:0] _12728 = {_0, _8894} + {_0, _11389};
  wire [3:0] _12729 = {_0, _12727} + {_0, _0, _12728};
  wire _12730 = _12301 < _12729;
  wire _12731 = r2000 ^ _12730;
  wire _12732 = _12298 ? coded_block[2000] : r2000;
  wire _12733 = _12296 ? _12731 : _12732;
  always @ (posedge reset or posedge clock) if (reset) r2000 <= 1'd0; else if (_12300) r2000 <= _12733;
  wire [1:0] _12734 = {_0, _1057} + {_0, _2941};
  wire [1:0] _12735 = {_0, _4958} + {_0, _7837};
  wire [2:0] _12736 = {_0, _12734} + {_0, _12735};
  wire [1:0] _12737 = {_0, _10172} + {_0, _11613};
  wire [3:0] _12738 = {_0, _12736} + {_0, _0, _12737};
  wire _12739 = _12301 < _12738;
  wire _12740 = r1999 ^ _12739;
  wire _12741 = _12298 ? coded_block[1999] : r1999;
  wire _12742 = _12296 ? _12740 : _12741;
  always @ (posedge reset or posedge clock) if (reset) r1999 <= 1'd0; else if (_12300) r1999 <= _12742;
  wire [1:0] _12743 = {_0, _1662} + {_0, _3742};
  wire [1:0] _12744 = {_0, _4574} + {_0, _7326};
  wire [2:0] _12745 = {_0, _12743} + {_0, _12744};
  wire [1:0] _12746 = {_0, _9279} + {_0, _11837};
  wire [3:0] _12747 = {_0, _12745} + {_0, _0, _12746};
  wire _12748 = _12301 < _12747;
  wire _12749 = r1998 ^ _12748;
  wire _12750 = _12298 ? coded_block[1998] : r1998;
  wire _12751 = _12296 ? _12749 : _12750;
  always @ (posedge reset or posedge clock) if (reset) r1998 <= 1'd0; else if (_12300) r1998 <= _12751;
  wire [1:0] _12752 = {_0, _289} + {_0, _3262};
  wire [1:0] _12753 = {_0, _4703} + {_0, _6589};
  wire [2:0] _12754 = {_0, _12752} + {_0, _12753};
  wire [1:0] _12755 = {_0, _8225} + {_0, _10717};
  wire [3:0] _12756 = {_0, _12754} + {_0, _0, _12755};
  wire _12757 = _12301 < _12756;
  wire _12758 = r1997 ^ _12757;
  wire _12759 = _12298 ? coded_block[1997] : r1997;
  wire _12760 = _12296 ? _12758 : _12759;
  always @ (posedge reset or posedge clock) if (reset) r1997 <= 1'd0; else if (_12300) r1997 <= _12760;
  wire [1:0] _12761 = {_0, _65} + {_0, _2782};
  wire [1:0] _12762 = {_0, _5407} + {_0, _7389};
  wire [2:0] _12763 = {_0, _12761} + {_0, _12762};
  wire [1:0] _12764 = {_0, _8543} + {_0, _11259};
  wire [3:0] _12765 = {_0, _12763} + {_0, _0, _12764};
  wire _12766 = _12301 < _12765;
  wire _12767 = r1996 ^ _12766;
  wire _12768 = _12298 ? coded_block[1996] : r1996;
  wire _12769 = _12296 ? _12767 : _12768;
  always @ (posedge reset or posedge clock) if (reset) r1996 <= 1'd0; else if (_12300) r1996 <= _12769;
  wire [1:0] _12770 = {_0, _1184} + {_0, _2144};
  wire [1:0] _12771 = {_0, _5597} + {_0, _7485};
  wire [2:0] _12772 = {_0, _12770} + {_0, _12771};
  wire [1:0] _12773 = {_0, _8225} + {_0, _11613};
  wire [3:0] _12774 = {_0, _12772} + {_0, _0, _12773};
  wire _12775 = _12301 < _12774;
  wire _12776 = r1995 ^ _12775;
  wire _12777 = _12298 ? coded_block[1995] : r1995;
  wire _12778 = _12296 ? _12776 : _12777;
  always @ (posedge reset or posedge clock) if (reset) r1995 <= 1'd0; else if (_12300) r1995 <= _12778;
  wire [1:0] _12779 = {_0, _65} + {_0, _2081};
  wire [1:0] _12780 = {_0, _4350} + {_0, _6589};
  wire [2:0] _12781 = {_0, _12779} + {_0, _12780};
  wire [1:0] _12782 = {_0, _9279} + {_0, _11069};
  wire [3:0] _12783 = {_0, _12781} + {_0, _0, _12782};
  wire _12784 = _12301 < _12783;
  wire _12785 = r1994 ^ _12784;
  wire _12786 = _12298 ? coded_block[1994] : r1994;
  wire _12787 = _12296 ? _12785 : _12786;
  always @ (posedge reset or posedge clock) if (reset) r1994 <= 1'd0; else if (_12300) r1994 <= _12787;
  wire [1:0] _12788 = {_0, _352} + {_0, _2782};
  wire [1:0] _12789 = {_0, _5470} + {_0, _7262};
  wire [2:0] _12790 = {_0, _12788} + {_0, _12789};
  wire [1:0] _12791 = {_0, _8511} + {_0, _10621};
  wire [3:0] _12792 = {_0, _12790} + {_0, _0, _12791};
  wire _12793 = _12301 < _12792;
  wire _12794 = r1993 ^ _12793;
  wire _12795 = _12298 ? coded_block[1993] : r1993;
  wire _12796 = _12296 ? _12794 : _12795;
  always @ (posedge reset or posedge clock) if (reset) r1993 <= 1'd0; else if (_12300) r1993 <= _12796;
  wire [1:0] _12797 = {_0, _1312} + {_0, _2081};
  wire [1:0] _12798 = {_0, _5597} + {_0, _7837};
  wire [2:0] _12799 = {_0, _12797} + {_0, _12798};
  wire [1:0] _12800 = {_0, _8511} + {_0, _10303};
  wire [3:0] _12801 = {_0, _12799} + {_0, _0, _12800};
  wire _12802 = _12301 < _12801;
  wire _12803 = r1992 ^ _12802;
  wire _12804 = _12298 ? coded_block[1992] : r1992;
  wire _12805 = _12296 ? _12803 : _12804;
  always @ (posedge reset or posedge clock) if (reset) r1992 <= 1'd0; else if (_12300) r1992 <= _12805;
  wire [1:0] _12806 = {_0, _1312} + {_0, _3933};
  wire [1:0] _12807 = {_0, _4703} + {_0, _7357};
  wire [2:0] _12808 = {_0, _12806} + {_0, _12807};
  wire [1:0] _12809 = {_0, _8957} + {_0, _10621};
  wire [3:0] _12810 = {_0, _12808} + {_0, _0, _12809};
  wire _12811 = _12301 < _12810;
  wire _12812 = r1991 ^ _12811;
  wire _12813 = _12298 ? coded_block[1991] : r1991;
  wire _12814 = _12296 ? _12812 : _12813;
  always @ (posedge reset or posedge clock) if (reset) r1991 <= 1'd0; else if (_12300) r1991 <= _12814;
  wire [1:0] _12815 = {_0, _958} + {_0, _3933};
  wire [1:0] _12816 = {_0, _5373} + {_0, _7262};
  wire [2:0] _12817 = {_0, _12815} + {_0, _12816};
  wire [1:0] _12818 = {_0, _8225} + {_0, _11389};
  wire [3:0] _12819 = {_0, _12817} + {_0, _0, _12818};
  wire _12820 = _12301 < _12819;
  wire _12821 = r1990 ^ _12820;
  wire _12822 = _12298 ? coded_block[1990] : r1990;
  wire _12823 = _12296 ? _12821 : _12822;
  always @ (posedge reset or posedge clock) if (reset) r1990 <= 1'd0; else if (_12300) r1990 <= _12823;
  wire [1:0] _12824 = {_0, _639} + {_0, _3294};
  wire [1:0] _12825 = {_0, _4574} + {_0, _6589};
  wire [2:0] _12826 = {_0, _12824} + {_0, _12825};
  wire [1:0] _12827 = {_0, _9469} + {_0, _11806};
  wire [3:0] _12828 = {_0, _12826} + {_0, _0, _12827};
  wire _12829 = _12301 < _12828;
  wire _12830 = r1989 ^ _12829;
  wire _12831 = _12298 ? coded_block[1989] : r1989;
  wire _12832 = _12296 ? _12830 : _12831;
  always @ (posedge reset or posedge clock) if (reset) r1989 <= 1'd0; else if (_12300) r1989 <= _12832;
  wire [1:0] _12833 = {_0, _958} + {_0, _3964};
  wire [1:0] _12834 = {_0, _5597} + {_0, _7357};
  wire [2:0] _12835 = {_0, _12833} + {_0, _12834};
  wire [1:0] _12836 = {_0, _8352} + {_0, _11900};
  wire [3:0] _12837 = {_0, _12835} + {_0, _0, _12836};
  wire _12838 = _12301 < _12837;
  wire _12839 = r1988 ^ _12838;
  wire _12840 = _12298 ? coded_block[1988] : r1988;
  wire _12841 = _12296 ? _12839 : _12840;
  always @ (posedge reset or posedge clock) if (reset) r1988 <= 1'd0; else if (_12300) r1988 <= _12841;
  wire [1:0] _12842 = {_0, _735} + {_0, _3964};
  wire [1:0] _12843 = {_0, _5116} + {_0, _7837};
  wire [2:0] _12844 = {_0, _12842} + {_0, _12843};
  wire [1:0] _12845 = {_0, _9469} + {_0, _11228};
  wire [3:0] _12846 = {_0, _12844} + {_0, _0, _12845};
  wire _12847 = _12301 < _12846;
  wire _12848 = r1987 ^ _12847;
  wire _12849 = _12298 ? coded_block[1987] : r1987;
  wire _12850 = _12296 ? _12848 : _12849;
  always @ (posedge reset or posedge clock) if (reset) r1987 <= 1'd0; else if (_12300) r1987 <= _12850;
  wire [1:0] _12851 = {_0, _639} + {_0, _2336};
  wire [1:0] _12852 = {_0, _5470} + {_0, _7837};
  wire [2:0] _12853 = {_0, _12851} + {_0, _12852};
  wire [1:0] _12854 = {_0, _8319} + {_0, _11740};
  wire [3:0] _12855 = {_0, _12853} + {_0, _0, _12854};
  wire _12856 = _12301 < _12855;
  wire _12857 = r1986 ^ _12856;
  wire _12858 = _12298 ? coded_block[1986] : r1986;
  wire _12859 = _12296 ? _12857 : _12858;
  always @ (posedge reset or posedge clock) if (reset) r1986 <= 1'd0; else if (_12300) r1986 <= _12859;
  wire [1:0] _12860 = {_0, _958} + {_0, _3805};
  wire [1:0] _12861 = {_0, _5116} + {_0, _6207};
  wire [2:0] _12862 = {_0, _12860} + {_0, _12861};
  wire [1:0] _12863 = {_0, _8799} + {_0, _11933};
  wire [3:0] _12864 = {_0, _12862} + {_0, _0, _12863};
  wire _12865 = _12301 < _12864;
  wire _12866 = r1985 ^ _12865;
  wire _12867 = _12298 ? coded_block[1985] : r1985;
  wire _12868 = _12296 ? _12866 : _12867;
  always @ (posedge reset or posedge clock) if (reset) r1985 <= 1'd0; else if (_12300) r1985 <= _12868;
  wire [1:0] _12869 = {_0, _1312} + {_0, _3805};
  wire [1:0] _12870 = {_0, _5022} + {_0, _6589};
  wire [2:0] _12871 = {_0, _12869} + {_0, _12870};
  wire [1:0] _12872 = {_0, _8767} + {_0, _12155};
  wire [3:0] _12873 = {_0, _12871} + {_0, _0, _12872};
  wire _12874 = _12301 < _12873;
  wire _12875 = r1984 ^ _12874;
  wire _12876 = _12298 ? coded_block[1984] : r1984;
  wire _12877 = _12296 ? _12875 : _12876;
  always @ (posedge reset or posedge clock) if (reset) r1984 <= 1'd0; else if (_12300) r1984 <= _12877;
  wire [1:0] _12878 = {_0, _1917} + {_0, _2782};
  wire [1:0] _12879 = {_0, _5534} + {_0, _7485};
  wire [2:0] _12880 = {_0, _12878} + {_0, _12879};
  wire [1:0] _12881 = {_0, _10045} + {_0, _10941};
  wire [3:0] _12882 = {_0, _12880} + {_0, _0, _12881};
  wire _12883 = _12301 < _12882;
  wire _12884 = r1983 ^ _12883;
  wire _12885 = _12298 ? coded_block[1983] : r1983;
  wire _12886 = _12296 ? _12884 : _12885;
  always @ (posedge reset or posedge clock) if (reset) r1983 <= 1'd0; else if (_12300) r1983 <= _12886;
  wire [1:0] _12887 = {_0, _352} + {_0, _2239};
  wire [1:0] _12888 = {_0, _4256} + {_0, _7132};
  wire [2:0] _12889 = {_0, _12887} + {_0, _12888};
  wire [1:0] _12890 = {_0, _9469} + {_0, _10910};
  wire [3:0] _12891 = {_0, _12889} + {_0, _0, _12890};
  wire _12892 = _12301 < _12891;
  wire _12893 = r1982 ^ _12892;
  wire _12894 = _12298 ? coded_block[1982] : r1982;
  wire _12895 = _12296 ? _12893 : _12894;
  always @ (posedge reset or posedge clock) if (reset) r1982 <= 1'd0; else if (_12300) r1982 <= _12895;
  wire [1:0] _12896 = {_0, _352} + {_0, _3453};
  wire [1:0] _12897 = {_0, _5949} + {_0, _7357};
  wire [2:0] _12898 = {_0, _12896} + {_0, _12897};
  wire [1:0] _12899 = {_0, _8319} + {_0, _10462};
  wire [3:0] _12900 = {_0, _12898} + {_0, _0, _12899};
  wire _12901 = _12301 < _12900;
  wire _12902 = r1981 ^ _12901;
  wire _12903 = _12298 ? coded_block[1981] : r1981;
  wire _12904 = _12296 ? _12902 : _12903;
  always @ (posedge reset or posedge clock) if (reset) r1981 <= 1'd0; else if (_12300) r1981 <= _12904;
  wire [1:0] _12905 = {_0, _958} + {_0, _2112};
  wire [1:0] _12906 = {_0, _4703} + {_0, _7837};
  wire [2:0] _12907 = {_0, _12905} + {_0, _12906};
  wire [1:0] _12908 = {_0, _10204} + {_0, _10685};
  wire [3:0] _12909 = {_0, _12907} + {_0, _0, _12908};
  wire _12910 = _12301 < _12909;
  wire _12911 = r1980 ^ _12910;
  wire _12912 = _12298 ? coded_block[1980] : r1980;
  wire _12913 = _12296 ? _12911 : _12912;
  always @ (posedge reset or posedge clock) if (reset) r1980 <= 1'd0; else if (_12300) r1980 <= _12913;
  wire [1:0] _12914 = {_0, _1568} + {_0, _2941};
  wire [1:0] _12915 = {_0, _5246} + {_0, _8186};
  wire [2:0] _12916 = {_0, _12914} + {_0, _12915};
  wire [1:0] _12917 = {_0, _9886} + {_0, _12155};
  wire [3:0] _12918 = {_0, _12916} + {_0, _0, _12917};
  wire _12919 = _12301 < _12918;
  wire _12920 = r1979 ^ _12919;
  wire _12921 = _12298 ? coded_block[1979] : r1979;
  wire _12922 = _12296 ? _12920 : _12921;
  always @ (posedge reset or posedge clock) if (reset) r1979 <= 1'd0; else if (_12300) r1979 <= _12922;
  wire [1:0] _12923 = {_0, _161} + {_0, _2112};
  wire [1:0] _12924 = {_0, _5726} + {_0, _7389};
  wire [2:0] _12925 = {_0, _12923} + {_0, _12924};
  wire [1:0] _12926 = {_0, _8446} + {_0, _10910};
  wire [3:0] _12927 = {_0, _12925} + {_0, _0, _12926};
  wire _12928 = _12301 < _12927;
  wire _12929 = r1978 ^ _12928;
  wire _12930 = _12298 ? coded_block[1978] : r1978;
  wire _12931 = _12296 ? _12929 : _12930;
  always @ (posedge reset or posedge clock) if (reset) r1978 <= 1'd0; else if (_12300) r1978 <= _12931;
  wire [1:0] _12932 = {_0, _161} + {_0, _3453};
  wire [1:0] _12933 = {_0, _5438} + {_0, _6589};
  wire [2:0] _12934 = {_0, _12932} + {_0, _12933};
  wire [1:0] _12935 = {_0, _9311} + {_0, _10941};
  wire [3:0] _12936 = {_0, _12934} + {_0, _0, _12935};
  wire _12937 = _12301 < _12936;
  wire _12938 = r1977 ^ _12937;
  wire _12939 = _12298 ? coded_block[1977] : r1977;
  wire _12940 = _12296 ? _12938 : _12939;
  always @ (posedge reset or posedge clock) if (reset) r1977 <= 1'd0; else if (_12300) r1977 <= _12940;
  wire [1:0] _12941 = {_0, _1184} + {_0, _3997};
  wire [1:0] _12942 = {_0, _5246} + {_0, _7357};
  wire [2:0] _12943 = {_0, _12941} + {_0, _12942};
  wire [1:0] _12944 = {_0, _10204} + {_0, _10941};
  wire [3:0] _12945 = {_0, _12943} + {_0, _0, _12944};
  wire _12946 = _12301 < _12945;
  wire _12947 = r1976 ^ _12946;
  wire _12948 = _12298 ? coded_block[1976] : r1976;
  wire _12949 = _12296 ? _12947 : _12948;
  always @ (posedge reset or posedge clock) if (reset) r1976 <= 1'd0; else if (_12300) r1976 <= _12949;
  wire [1:0] _12950 = {_0, _2044} + {_0, _3836};
  wire [1:0] _12951 = {_0, _5022} + {_0, _6845};
  wire [2:0] _12952 = {_0, _12950} + {_0, _12951};
  wire [1:0] _12953 = {_0, _9469} + {_0, _11453};
  wire [3:0] _12954 = {_0, _12952} + {_0, _0, _12953};
  wire _12955 = _12301 < _12954;
  wire _12956 = r1975 ^ _12955;
  wire _12957 = _12298 ? coded_block[1975] : r1975;
  wire _12958 = _12296 ? _12956 : _12957;
  always @ (posedge reset or posedge clock) if (reset) r1975 <= 1'd0; else if (_12300) r1975 <= _12958;
  wire [1:0] _12959 = {_0, _1312} + {_0, _3773};
  wire [1:0] _12960 = {_0, _5116} + {_0, _6845};
  wire [2:0] _12961 = {_0, _12959} + {_0, _12960};
  wire [1:0] _12962 = {_0, _9054} + {_0, _10910};
  wire [3:0] _12963 = {_0, _12961} + {_0, _0, _12962};
  wire _12964 = _12301 < _12963;
  wire _12965 = r1974 ^ _12964;
  wire _12966 = _12298 ? coded_block[1974] : r1974;
  wire _12967 = _12296 ? _12965 : _12966;
  always @ (posedge reset or posedge clock) if (reset) r1974 <= 1'd0; else if (_12300) r1974 <= _12967;
  wire [1:0] _12968 = {_0, _1057} + {_0, _2623};
  wire [1:0] _12969 = {_0, _4574} + {_0, _7132};
  wire [2:0] _12970 = {_0, _12968} + {_0, _12969};
  wire [1:0] _12971 = {_0, _10045} + {_0, _11358};
  wire [3:0] _12972 = {_0, _12970} + {_0, _0, _12971};
  wire _12973 = _12301 < _12972;
  wire _12974 = r1973 ^ _12973;
  wire _12975 = _12298 ? coded_block[1973] : r1973;
  wire _12976 = _12296 ? _12974 : _12975;
  always @ (posedge reset or posedge clock) if (reset) r1973 <= 1'd0; else if (_12300) r1973 <= _12976;
  wire [1:0] _12977 = {_0, _1950} + {_0, _2878};
  wire [1:0] _12978 = {_0, _4703} + {_0, _7326};
  wire [2:0] _12979 = {_0, _12977} + {_0, _12978};
  wire [1:0] _12980 = {_0, _9311} + {_0, _10462};
  wire [3:0] _12981 = {_0, _12979} + {_0, _0, _12980};
  wire _12982 = _12301 < _12981;
  wire _12983 = r1972 ^ _12982;
  wire _12984 = _12298 ? coded_block[1972] : r1972;
  wire _12985 = _12296 ? _12983 : _12984;
  always @ (posedge reset or posedge clock) if (reset) r1972 <= 1'd0; else if (_12300) r1972 <= _12985;
  wire [1:0] _12986 = {_0, _352} + {_0, _2623};
  wire [1:0] _12987 = {_0, _5022} + {_0, _7804};
  wire [2:0] _12988 = {_0, _12986} + {_0, _12987};
  wire [1:0] _12989 = {_0, _8446} + {_0, _12061};
  wire [3:0] _12990 = {_0, _12988} + {_0, _0, _12989};
  wire _12991 = _12301 < _12990;
  wire _12992 = r1971 ^ _12991;
  wire _12993 = _12298 ? coded_block[1971] : r1971;
  wire _12994 = _12296 ? _12992 : _12993;
  always @ (posedge reset or posedge clock) if (reset) r1971 <= 1'd0; else if (_12300) r1971 <= _12994;
  wire [1:0] _12995 = {_0, _2044} + {_0, _3997};
  wire [1:0] _12996 = {_0, _5597} + {_0, _7262};
  wire [2:0] _12997 = {_0, _12995} + {_0, _12996};
  wire [1:0] _12998 = {_0, _8319} + {_0, _10783};
  wire [3:0] _12999 = {_0, _12997} + {_0, _0, _12998};
  wire _13000 = _12301 < _12999;
  wire _13001 = r1970 ^ _13000;
  wire _13002 = _12298 ? coded_block[1970] : r1970;
  wire _13003 = _12296 ? _13001 : _13002;
  always @ (posedge reset or posedge clock) if (reset) r1970 <= 1'd0; else if (_12300) r1970 <= _13003;
  wire [1:0] _13004 = {_0, _1184} + {_0, _3836};
  wire [1:0] _13005 = {_0, _5116} + {_0, _7132};
  wire [2:0] _13006 = {_0, _13004} + {_0, _13005};
  wire [1:0] _13007 = {_0, _10014} + {_0, _10335};
  wire [3:0] _13008 = {_0, _13006} + {_0, _0, _13007};
  wire _13009 = _12301 < _13008;
  wire _13010 = r1969 ^ _13009;
  wire _13011 = _12298 ? coded_block[1969] : r1969;
  wire _13012 = _12296 ? _13010 : _13011;
  always @ (posedge reset or posedge clock) if (reset) r1969 <= 1'd0; else if (_12300) r1969 <= _13012;
  wire [1:0] _13013 = {_0, _1533} + {_0, _3167};
  wire [1:0] _13014 = {_0, _6108} + {_0, _7804};
  wire [2:0] _13015 = {_0, _13013} + {_0, _13014};
  wire [1:0] _13016 = {_0, _10077} + {_0, _11996};
  wire [3:0] _13017 = {_0, _13015} + {_0, _0, _13016};
  wire _13018 = _12301 < _13017;
  wire _13019 = r1968 ^ _13018;
  wire _13020 = _12298 ? coded_block[1968] : r1968;
  wire _13021 = _12296 ? _13019 : _13020;
  always @ (posedge reset or posedge clock) if (reset) r1968 <= 1'd0; else if (_12300) r1968 <= _13021;
  wire [1:0] _13022 = {_0, _2044} + {_0, _2592};
  wire [1:0] _13023 = {_0, _5116} + {_0, _6589};
  wire [2:0] _13024 = {_0, _13022} + {_0, _13023};
  wire [1:0] _13025 = {_0, _9949} + {_0, _11677};
  wire [3:0] _13026 = {_0, _13024} + {_0, _0, _13025};
  wire _13027 = _12301 < _13026;
  wire _13028 = r1967 ^ _13027;
  wire _13029 = _12298 ? coded_block[1967] : r1967;
  wire _13030 = _12296 ? _13028 : _13029;
  always @ (posedge reset or posedge clock) if (reset) r1967 <= 1'd0; else if (_12300) r1967 <= _13030;
  wire [1:0] _13031 = {_0, _1950} + {_0, _3390};
  wire [1:0] _13032 = {_0, _5597} + {_0, _7454};
  wire [2:0] _13033 = {_0, _13031} + {_0, _13032};
  wire [1:0] _13034 = {_0, _9886} + {_0, _11069};
  wire [3:0] _13035 = {_0, _13033} + {_0, _0, _13034};
  wire _13036 = _12301 < _13035;
  wire _13037 = r1966 ^ _13036;
  wire _13038 = _12298 ? coded_block[1966] : r1966;
  wire _13039 = _12296 ? _13037 : _13038;
  always @ (posedge reset or posedge clock) if (reset) r1966 <= 1'd0; else if (_12300) r1966 <= _13039;
  wire [1:0] _13040 = {_0, _289} + {_0, _3773};
  wire [1:0] _13041 = {_0, _4319} + {_0, _7230};
  wire [2:0] _13042 = {_0, _13040} + {_0, _13041};
  wire [1:0] _13043 = {_0, _8543} + {_0, _11644};
  wire [3:0] _13044 = {_0, _13042} + {_0, _0, _13043};
  wire _13045 = _12301 < _13044;
  wire _13046 = r1965 ^ _13045;
  wire _13047 = _12298 ? coded_block[1965] : r1965;
  wire _13048 = _12296 ? _13046 : _13047;
  always @ (posedge reset or posedge clock) if (reset) r1965 <= 1'd0; else if (_12300) r1965 <= _13048;
  wire [1:0] _13049 = {_0, _639} + {_0, _4028};
  wire [1:0] _13050 = {_0, _4319} + {_0, _7262};
  wire [2:0] _13051 = {_0, _13049} + {_0, _13050};
  wire [1:0] _13052 = {_0, _8957} + {_0, _11228};
  wire [3:0] _13053 = {_0, _13051} + {_0, _0, _13052};
  wire _13054 = _12301 < _13053;
  wire _13055 = r1964 ^ _13054;
  wire _13056 = _12298 ? coded_block[1964] : r1964;
  wire _13057 = _12296 ? _13055 : _13056;
  always @ (posedge reset or posedge clock) if (reset) r1964 <= 1'd0; else if (_12300) r1964 <= _13057;
  wire [1:0] _13058 = {_0, _2044} + {_0, _3422};
  wire [1:0] _13059 = {_0, _5726} + {_0, _6652};
  wire [2:0] _13060 = {_0, _13058} + {_0, _13059};
  wire [1:0] _13061 = {_0, _8352} + {_0, _10621};
  wire [3:0] _13062 = {_0, _13060} + {_0, _0, _13061};
  wire _13063 = _12301 < _13062;
  wire _13064 = r1963 ^ _13063;
  wire _13065 = _12298 ? coded_block[1963] : r1963;
  wire _13066 = _12296 ? _13064 : _13065;
  always @ (posedge reset or posedge clock) if (reset) r1963 <= 1'd0; else if (_12300) r1963 <= _13066;
  wire [1:0] _13067 = {_0, _1021} + {_0, _3997};
  wire [1:0] _13068 = {_0, _5438} + {_0, _7326};
  wire [2:0] _13069 = {_0, _13067} + {_0, _13068};
  wire [1:0] _13070 = {_0, _8225} + {_0, _11453};
  wire [3:0] _13071 = {_0, _13069} + {_0, _0, _13070};
  wire _13072 = _12301 < _13071;
  wire _13073 = r1962 ^ _13072;
  wire _13074 = _12298 ? coded_block[1962] : r1962;
  wire _13075 = _12296 ? _13073 : _13074;
  always @ (posedge reset or posedge clock) if (reset) r1962 <= 1'd0; else if (_12300) r1962 <= _13075;
  wire [1:0] _13076 = {_0, _510} + {_0, _2592};
  wire [1:0] _13077 = {_0, _5438} + {_0, _8186};
  wire [2:0] _13078 = {_0, _13076} + {_0, _13077};
  wire [1:0] _13079 = {_0, _10141} + {_0, _10685};
  wire [3:0] _13080 = {_0, _13078} + {_0, _0, _13079};
  wire _13081 = _12301 < _13080;
  wire _13082 = r1961 ^ _13081;
  wire _13083 = _12298 ? coded_block[1961] : r1961;
  wire _13084 = _12296 ? _13082 : _13083;
  always @ (posedge reset or posedge clock) if (reset) r1961 <= 1'd0; else if (_12300) r1961 <= _13084;
  wire [1:0] _13085 = {_0, _958} + {_0, _2081};
  wire [1:0] _13086 = {_0, _5246} + {_0, _7485};
  wire [2:0] _13087 = {_0, _13085} + {_0, _13086};
  wire [1:0] _13088 = {_0, _10172} + {_0, _11964};
  wire [3:0] _13089 = {_0, _13087} + {_0, _0, _13088};
  wire _13090 = _12301 < _13089;
  wire _13091 = r1960 ^ _13090;
  wire _13092 = _12298 ? coded_block[1960] : r1960;
  wire _13093 = _12296 ? _13091 : _13092;
  always @ (posedge reset or posedge clock) if (reset) r1960 <= 1'd0; else if (_12300) r1960 <= _13093;
  wire [1:0] _13094 = {_0, _1057} + {_0, _4028};
  wire [1:0] _13095 = {_0, _5470} + {_0, _7357};
  wire [2:0] _13096 = {_0, _13094} + {_0, _13095};
  wire [1:0] _13097 = {_0, _8225} + {_0, _11485};
  wire [3:0] _13098 = {_0, _13096} + {_0, _0, _13097};
  wire _13099 = _12301 < _13098;
  wire _13100 = r1959 ^ _13099;
  wire _13101 = _12298 ? coded_block[1959] : r1959;
  wire _13102 = _12296 ? _13100 : _13101;
  always @ (posedge reset or posedge clock) if (reset) r1959 <= 1'd0; else if (_12300) r1959 <= _13102;
  wire [1:0] _13103 = {_0, _1057} + {_0, _3870};
  wire [1:0] _13104 = {_0, _5116} + {_0, _7230};
  wire [2:0] _13105 = {_0, _13103} + {_0, _13104};
  wire [1:0] _13106 = {_0, _10077} + {_0, _10814};
  wire [3:0] _13107 = {_0, _13105} + {_0, _0, _13106};
  wire _13108 = _12301 < _13107;
  wire _13109 = r1958 ^ _13108;
  wire _13110 = _12298 ? coded_block[1958] : r1958;
  wire _13111 = _12296 ? _13109 : _13110;
  always @ (posedge reset or posedge clock) if (reset) r1958 <= 1'd0; else if (_12300) r1958 <= _13111;
  wire [1:0] _13112 = {_0, _639} + {_0, _2623};
  wire [1:0] _13113 = {_0, _5534} + {_0, _6845};
  wire [2:0] _13114 = {_0, _13112} + {_0, _13113};
  wire [1:0] _13115 = {_0, _9949} + {_0, _10527};
  wire [3:0] _13116 = {_0, _13114} + {_0, _0, _13115};
  wire _13117 = _12301 < _13116;
  wire _13118 = r1957 ^ _13117;
  wire _13119 = _12298 ? coded_block[1957] : r1957;
  wire _13120 = _12296 ? _13118 : _13119;
  always @ (posedge reset or posedge clock) if (reset) r1957 <= 1'd0; else if (_12300) r1957 <= _13120;
  wire [1:0] _13121 = {_0, _1533} + {_0, _2623};
  wire [1:0] _13122 = {_0, _5116} + {_0, _6525};
  wire [2:0] _13123 = {_0, _13121} + {_0, _13122};
  wire [1:0] _13124 = {_0, _9503} + {_0, _11644};
  wire [3:0] _13125 = {_0, _13123} + {_0, _0, _13124};
  wire _13126 = _12301 < _13125;
  wire _13127 = r1956 ^ _13126;
  wire _13128 = _12298 ? coded_block[1956] : r1956;
  wire _13129 = _12296 ? _13127 : _13128;
  always @ (posedge reset or posedge clock) if (reset) r1956 <= 1'd0; else if (_12300) r1956 <= _13129;
  wire [1:0] _13130 = {_0, _958} + {_0, _3836};
  wire [1:0] _13131 = {_0, _4574} + {_0, _6525};
  wire [2:0] _13132 = {_0, _13130} + {_0, _13131};
  wire [1:0] _13133 = {_0, _9085} + {_0, _11996};
  wire [3:0] _13134 = {_0, _13132} + {_0, _0, _13133};
  wire _13135 = _12301 < _13134;
  wire _13136 = r1955 ^ _13135;
  wire _13137 = _12298 ? coded_block[1955] : r1955;
  wire _13138 = _12296 ? _13136 : _13137;
  always @ (posedge reset or posedge clock) if (reset) r1955 <= 1'd0; else if (_12300) r1955 <= _13138;
  wire [1:0] _13139 = {_0, _1568} + {_0, _2782};
  wire [1:0] _13140 = {_0, _5949} + {_0, _6652};
  wire [2:0] _13141 = {_0, _13139} + {_0, _13140};
  wire [1:0] _13142 = {_0, _8288} + {_0, _12061};
  wire [3:0] _13143 = {_0, _13141} + {_0, _0, _13142};
  wire _13144 = _12301 < _13143;
  wire _13145 = r1954 ^ _13144;
  wire _13146 = _12298 ? coded_block[1954] : r1954;
  wire _13147 = _12296 ? _13145 : _13146;
  always @ (posedge reset or posedge clock) if (reset) r1954 <= 1'd0; else if (_12300) r1954 <= _13147;
  wire [1:0] _13148 = {_0, _510} + {_0, _3422};
  wire [1:0] _13149 = {_0, _4384} + {_0, _6525};
  wire [2:0] _13150 = {_0, _13148} + {_0, _13149};
  wire [1:0] _13151 = {_0, _10045} + {_0, _10335};
  wire [3:0] _13152 = {_0, _13150} + {_0, _0, _13151};
  wire _13153 = _12301 < _13152;
  wire _13154 = r1953 ^ _13153;
  wire _13155 = _12298 ? coded_block[1953] : r1953;
  wire _13156 = _12296 ? _13154 : _13155;
  always @ (posedge reset or posedge clock) if (reset) r1953 <= 1'd0; else if (_12300) r1953 <= _13156;
  wire [1:0] _13157 = {_0, _1021} + {_0, _2302};
  wire [1:0] _13158 = {_0, _4287} + {_0, _7454};
  wire [2:0] _13159 = {_0, _13157} + {_0, _13158};
  wire [1:0] _13160 = {_0, _10172} + {_0, _11806};
  wire [3:0] _13161 = {_0, _13159} + {_0, _0, _13160};
  wire _13162 = _12301 < _13161;
  wire _13163 = r1952 ^ _13162;
  wire _13164 = _12298 ? coded_block[1952] : r1952;
  wire _13165 = _12296 ? _13163 : _13164;
  always @ (posedge reset or posedge clock) if (reset) r1952 <= 1'd0; else if (_12300) r1952 <= _13165;
  wire [1:0] _13166 = {_0, _383} + {_0, _2239};
  wire [1:0] _13167 = {_0, _5116} + {_0, _7454};
  wire [2:0] _13168 = {_0, _13166} + {_0, _13167};
  wire [1:0] _13169 = {_0, _8894} + {_0, _10783};
  wire [3:0] _13170 = {_0, _13168} + {_0, _0, _13169};
  wire _13171 = _12301 < _13170;
  wire _13172 = r1951 ^ _13171;
  wire _13173 = _12298 ? coded_block[1951] : r1951;
  wire _13174 = _12296 ? _13172 : _13173;
  always @ (posedge reset or posedge clock) if (reset) r1951 <= 1'd0; else if (_12300) r1951 <= _13174;
  wire [1:0] _13175 = {_0, _1184} + {_0, _2557};
  wire [1:0] _13176 = {_0, _4861} + {_0, _7804};
  wire [2:0] _13177 = {_0, _13175} + {_0, _13176};
  wire [1:0] _13178 = {_0, _9503} + {_0, _11771};
  wire [3:0] _13179 = {_0, _13177} + {_0, _0, _13178};
  wire _13180 = _12301 < _13179;
  wire _13181 = r1950 ^ _13180;
  wire _13182 = _12298 ? coded_block[1950] : r1950;
  wire _13183 = _12296 ? _13181 : _13182;
  always @ (posedge reset or posedge clock) if (reset) r1950 <= 1'd0; else if (_12300) r1950 <= _13183;
  wire [1:0] _13184 = {_0, _2044} + {_0, _2623};
  wire [1:0] _13185 = {_0, _4384} + {_0, _7389};
  wire [2:0] _13186 = {_0, _13184} + {_0, _13185};
  wire [1:0] _13187 = {_0, _8926} + {_0, _11964};
  wire [3:0] _13188 = {_0, _13186} + {_0, _0, _13187};
  wire _13189 = _12301 < _13188;
  wire _13190 = r1949 ^ _13189;
  wire _13191 = _12298 ? coded_block[1949] : r1949;
  wire _13192 = _12296 ? _13190 : _13191;
  always @ (posedge reset or posedge clock) if (reset) r1949 <= 1'd0; else if (_12300) r1949 <= _13192;
  wire [1:0] _13193 = {_0, _97} + {_0, _2239};
  wire [1:0] _13194 = {_0, _4703} + {_0, _7230};
  wire [2:0] _13195 = {_0, _13193} + {_0, _13194};
  wire [1:0] _13196 = {_0, _8701} + {_0, _12061};
  wire [3:0] _13197 = {_0, _13195} + {_0, _0, _13196};
  wire _13198 = _12301 < _13197;
  wire _13199 = r1948 ^ _13198;
  wire _13200 = _12298 ? coded_block[1948] : r1948;
  wire _13201 = _12296 ? _13199 : _13200;
  always @ (posedge reset or posedge clock) if (reset) r1948 <= 1'd0; else if (_12300) r1948 <= _13201;
  wire [1:0] _13202 = {_0, _1184} + {_0, _3742};
  wire [1:0] _13203 = {_0, _4256} + {_0, _7741};
  wire [2:0] _13204 = {_0, _13202} + {_0, _13203};
  wire [1:0] _13205 = {_0, _9085} + {_0, _10814};
  wire [3:0] _13206 = {_0, _13204} + {_0, _0, _13205};
  wire _13207 = _12301 < _13206;
  wire _13208 = r1947 ^ _13207;
  wire _13209 = _12298 ? coded_block[1947] : r1947;
  wire _13210 = _12296 ? _13208 : _13209;
  always @ (posedge reset or posedge clock) if (reset) r1947 <= 1'd0; else if (_12300) r1947 <= _13210;
  wire [1:0] _13211 = {_0, _383} + {_0, _2782};
  wire [1:0] _13212 = {_0, _4703} + {_0, _7100};
  wire [2:0] _13213 = {_0, _13211} + {_0, _13212};
  wire [1:0] _13214 = {_0, _9886} + {_0, _10527};
  wire [3:0] _13215 = {_0, _13213} + {_0, _0, _13214};
  wire _13216 = _12301 < _13215;
  wire _13217 = r1946 ^ _13216;
  wire _13218 = _12298 ? coded_block[1946] : r1946;
  wire _13219 = _12296 ? _13217 : _13218;
  always @ (posedge reset or posedge clock) if (reset) r1946 <= 1'd0; else if (_12300) r1946 <= _13219;
  wire [1:0] _13220 = {_0, _1695} + {_0, _3836};
  wire [1:0] _13221 = {_0, _4287} + {_0, _6814};
  wire [2:0] _13222 = {_0, _13220} + {_0, _13221};
  wire [1:0] _13223 = {_0, _8288} + {_0, _11644};
  wire [3:0] _13224 = {_0, _13222} + {_0, _0, _13223};
  wire _13225 = _12301 < _13224;
  wire _13226 = r1945 ^ _13225;
  wire _13227 = _12298 ? coded_block[1945] : r1945;
  wire _13228 = _12296 ? _13226 : _13227;
  always @ (posedge reset or posedge clock) if (reset) r1945 <= 1'd0; else if (_12300) r1945 <= _13228;
  wire [1:0] _13229 = {_0, _161} + {_0, _2782};
  wire [1:0] _13230 = {_0, _5565} + {_0, _6207};
  wire [2:0] _13231 = {_0, _13229} + {_0, _13230};
  wire [1:0] _13232 = {_0, _9822} + {_0, _11485};
  wire [3:0] _13233 = {_0, _13231} + {_0, _0, _13232};
  wire _13234 = _12301 < _13233;
  wire _13235 = r1944 ^ _13234;
  wire _13236 = _12298 ? coded_block[1944] : r1944;
  wire _13237 = _12296 ? _13235 : _13236;
  always @ (posedge reset or posedge clock) if (reset) r1944 <= 1'd0; else if (_12300) r1944 <= _13237;
  wire [1:0] _13238 = {_0, _1057} + {_0, _3037};
  wire [1:0] _13239 = {_0, _5949} + {_0, _7262};
  wire [2:0] _13240 = {_0, _13238} + {_0, _13239};
  wire [1:0] _13241 = {_0, _8352} + {_0, _10941};
  wire [3:0] _13242 = {_0, _13240} + {_0, _0, _13241};
  wire _13243 = _12301 < _13242;
  wire _13244 = r1943 ^ _13243;
  wire _13245 = _12298 ? coded_block[1943] : r1943;
  wire _13246 = _12296 ? _13244 : _13245;
  always @ (posedge reset or posedge clock) if (reset) r1943 <= 1'd0; else if (_12300) r1943 <= _13246;
  wire [1:0] _13247 = {_0, _128} + {_0, _3836};
  wire [1:0] _13248 = {_0, _4958} + {_0, _7326};
  wire [2:0] _13249 = {_0, _13247} + {_0, _13248};
  wire [1:0] _13250 = {_0, _9822} + {_0, _11228};
  wire [3:0] _13251 = {_0, _13249} + {_0, _0, _13250};
  wire _13252 = _12301 < _13251;
  wire _13253 = r1942 ^ _13252;
  wire _13254 = _12298 ? coded_block[1942] : r1942;
  wire _13255 = _12296 ? _13253 : _13254;
  always @ (posedge reset or posedge clock) if (reset) r1942 <= 1'd0; else if (_12300) r1942 <= _13255;
  wire [1:0] _13256 = {_0, _735} + {_0, _3836};
  wire [1:0] _13257 = {_0, _4319} + {_0, _7741};
  wire [2:0] _13258 = {_0, _13256} + {_0, _13257};
  wire [1:0] _13259 = {_0, _8701} + {_0, _10846};
  wire [3:0] _13260 = {_0, _13258} + {_0, _0, _13259};
  wire _13261 = _12301 < _13260;
  wire _13262 = r1941 ^ _13261;
  wire _13263 = _12298 ? coded_block[1941] : r1941;
  wire _13264 = _12296 ? _13262 : _13263;
  always @ (posedge reset or posedge clock) if (reset) r1941 <= 1'd0; else if (_12300) r1941 <= _13264;
  wire [1:0] _13265 = {_0, _128} + {_0, _2144};
  wire [1:0] _13266 = {_0, _4256} + {_0, _7100};
  wire [2:0] _13267 = {_0, _13265} + {_0, _13266};
  wire [1:0] _13268 = {_0, _9853} + {_0, _11806};
  wire [3:0] _13269 = {_0, _13267} + {_0, _0, _13268};
  wire _13270 = _12301 < _13269;
  wire _13271 = r1940 ^ _13270;
  wire _13272 = _12298 ? coded_block[1940] : r1940;
  wire _13273 = _12296 ? _13271 : _13272;
  always @ (posedge reset or posedge clock) if (reset) r1940 <= 1'd0; else if (_12300) r1940 <= _13273;
  wire [1:0] _13274 = {_0, _1662} + {_0, _3517};
  wire [1:0] _13275 = {_0, _4384} + {_0, _6718};
  wire [2:0] _13276 = {_0, _13274} + {_0, _13275};
  wire [1:0] _13277 = {_0, _10172} + {_0, _12061};
  wire [3:0] _13278 = {_0, _13276} + {_0, _0, _13277};
  wire _13279 = _12301 < _13278;
  wire _13280 = r1939 ^ _13279;
  wire _13281 = _12298 ? coded_block[1939] : r1939;
  wire _13282 = _12296 ? _13280 : _13281;
  always @ (posedge reset or posedge clock) if (reset) r1939 <= 1'd0; else if (_12300) r1939 <= _13282;
  wire [1:0] _13283 = {_0, _1568} + {_0, _3422};
  wire [1:0] _13284 = {_0, _4287} + {_0, _6621};
  wire [2:0] _13285 = {_0, _13283} + {_0, _13284};
  wire [1:0] _13286 = {_0, _10077} + {_0, _11964};
  wire [3:0] _13287 = {_0, _13285} + {_0, _0, _13286};
  wire _13288 = _12301 < _13287;
  wire _13289 = r1938 ^ _13288;
  wire _13290 = _12298 ? coded_block[1938] : r1938;
  wire _13291 = _12296 ? _13289 : _13290;
  always @ (posedge reset or posedge clock) if (reset) r1938 <= 1'd0; else if (_12300) r1938 <= _13291;
  wire [1:0] _13292 = {_0, _510} + {_0, _2302};
  wire [1:0] _13293 = {_0, _5501} + {_0, _7326};
  wire [2:0] _13294 = {_0, _13292} + {_0, _13293};
  wire [1:0] _13295 = {_0, _9949} + {_0, _11933};
  wire [3:0] _13296 = {_0, _13294} + {_0, _0, _13295};
  wire _13297 = _12301 < _13296;
  wire _13298 = r1937 ^ _13297;
  wire _13299 = _12298 ? coded_block[1937] : r1937;
  wire _13300 = _12296 ? _13298 : _13299;
  always @ (posedge reset or posedge clock) if (reset) r1937 <= 1'd0; else if (_12300) r1937 <= _13300;
  wire [1:0] _13301 = {_0, _1758} + {_0, _3037};
  wire [1:0] _13302 = {_0, _5022} + {_0, _8186};
  wire [2:0] _13303 = {_0, _13301} + {_0, _13302};
  wire [1:0] _13304 = {_0, _8894} + {_0, _10527};
  wire [3:0] _13305 = {_0, _13303} + {_0, _0, _13304};
  wire _13306 = _12301 < _13305;
  wire _13307 = r1936 ^ _13306;
  wire _13308 = _12298 ? coded_block[1936] : r1936;
  wire _13309 = _12296 ? _13307 : _13308;
  always @ (posedge reset or posedge clock) if (reset) r1936 <= 1'd0; else if (_12300) r1936 <= _13309;
  wire [1:0] _13310 = {_0, _894} + {_0, _2878};
  wire [1:0] _13311 = {_0, _5790} + {_0, _7100};
  wire [2:0] _13312 = {_0, _13310} + {_0, _13311};
  wire [1:0] _13313 = {_0, _10204} + {_0, _10783};
  wire [3:0] _13314 = {_0, _13312} + {_0, _0, _13313};
  wire _13315 = _12301 < _13314;
  wire _13316 = r1935 ^ _13315;
  wire _13317 = _12298 ? coded_block[1935] : r1935;
  wire _13318 = _12296 ? _13316 : _13317;
  always @ (posedge reset or posedge clock) if (reset) r1935 <= 1'd0; else if (_12300) r1935 <= _13318;
  wire [1:0] _13319 = {_0, _703} + {_0, _3773};
  wire [1:0] _13320 = {_0, _5565} + {_0, _6814};
  wire [2:0] _13321 = {_0, _13319} + {_0, _13320};
  wire [1:0] _13322 = {_0, _8926} + {_0, _11771};
  wire [3:0] _13323 = {_0, _13321} + {_0, _0, _13322};
  wire _13324 = _12301 < _13323;
  wire _13325 = r1934 ^ _13324;
  wire _13326 = _12298 ? coded_block[1934] : r1934;
  wire _13327 = _12296 ? _13325 : _13326;
  always @ (posedge reset or posedge clock) if (reset) r1934 <= 1'd0; else if (_12300) r1934 <= _13327;
  wire [1:0] _13328 = {_0, _894} + {_0, _3037};
  wire [1:0] _13329 = {_0, _5501} + {_0, _8028};
  wire [2:0] _13330 = {_0, _13328} + {_0, _13329};
  wire [1:0] _13331 = {_0, _9503} + {_0, _10846};
  wire [3:0] _13332 = {_0, _13330} + {_0, _0, _13331};
  wire _13333 = _12301 < _13332;
  wire _13334 = r1933 ^ _13333;
  wire _13335 = _12298 ? coded_block[1933] : r1933;
  wire _13336 = _12296 ? _13334 : _13335;
  always @ (posedge reset or posedge clock) if (reset) r1933 <= 1'd0; else if (_12300) r1933 <= _13336;
  wire [1:0] _13337 = {_0, _703} + {_0, _3997};
  wire [1:0] _13338 = {_0, _5981} + {_0, _7132};
  wire [2:0] _13339 = {_0, _13337} + {_0, _13338};
  wire [1:0] _13340 = {_0, _9853} + {_0, _11485};
  wire [3:0] _13341 = {_0, _13339} + {_0, _0, _13340};
  wire _13342 = _12301 < _13341;
  wire _13343 = r1932 ^ _13342;
  wire _13344 = _12298 ? coded_block[1932] : r1932;
  wire _13345 = _12296 ? _13343 : _13344;
  always @ (posedge reset or posedge clock) if (reset) r1932 <= 1'd0; else if (_12300) r1932 <= _13345;
  wire [1:0] _13346 = {_0, _1758} + {_0, _3773};
  wire [1:0] _13347 = {_0, _5884} + {_0, _6718};
  wire [2:0] _13348 = {_0, _13346} + {_0, _13347};
  wire [1:0] _13349 = {_0, _9469} + {_0, _11422};
  wire [3:0] _13350 = {_0, _13348} + {_0, _0, _13349};
  wire _13351 = _12301 < _13350;
  wire _13352 = r1931 ^ _13351;
  wire _13353 = _12298 ? coded_block[1931] : r1931;
  wire _13354 = _12296 ? _13352 : _13353;
  always @ (posedge reset or posedge clock) if (reset) r1931 <= 1'd0; else if (_12300) r1931 <= _13354;
  wire [1:0] _13355 = {_0, _1726} + {_0, _2144};
  wire [1:0] _13356 = {_0, _4830} + {_0, _6621};
  wire [2:0] _13357 = {_0, _13355} + {_0, _13356};
  wire [1:0] _13358 = {_0, _9886} + {_0, _11996};
  wire [3:0] _13359 = {_0, _13357} + {_0, _0, _13358};
  wire _13360 = _12301 < _13359;
  wire _13361 = r1930 ^ _13360;
  wire _13362 = _12298 ? coded_block[1930] : r1930;
  wire _13363 = _12296 ? _13361 : _13362;
  always @ (posedge reset or posedge clock) if (reset) r1930 <= 1'd0; else if (_12300) r1930 <= _13363;
  wire [1:0] _13364 = {_0, _1886} + {_0, _2847};
  wire [1:0] _13365 = {_0, _4287} + {_0, _8186};
  wire [2:0] _13366 = {_0, _13364} + {_0, _13365};
  wire [1:0] _13367 = {_0, _8225} + {_0, _10303};
  wire [3:0] _13368 = {_0, _13366} + {_0, _0, _13367};
  wire _13369 = _12301 < _13368;
  wire _13370 = r1929 ^ _13369;
  wire _13371 = _12298 ? coded_block[1929] : r1929;
  wire _13372 = _12296 ? _13370 : _13371;
  always @ (posedge reset or posedge clock) if (reset) r1929 <= 1'd0; else if (_12300) r1929 <= _13372;
  wire [1:0] _13373 = {_0, _1886} + {_0, _3933};
  wire [1:0] _13374 = {_0, _5981} + {_0, _8028};
  wire [2:0] _13375 = {_0, _13373} + {_0, _13374};
  wire [1:0] _13376 = {_0, _10077} + {_0, _12124};
  wire [3:0] _13377 = {_0, _13375} + {_0, _0, _13376};
  wire _13378 = _12301 < _13377;
  wire _13379 = r1928 ^ _13378;
  wire _13380 = _12298 ? coded_block[1928] : r1928;
  wire _13381 = _12296 ? _13379 : _13380;
  always @ (posedge reset or posedge clock) if (reset) r1928 <= 1'd0; else if (_12300) r1928 <= _13381;
  wire [1:0] _13382 = {_0, _1917} + {_0, _3517};
  wire [1:0] _13383 = {_0, _5373} + {_0, _7804};
  wire [2:0] _13384 = {_0, _13382} + {_0, _13383};
  wire [1:0] _13385 = {_0, _8991} + {_0, _10814};
  wire [3:0] _13386 = {_0, _13384} + {_0, _0, _13385};
  wire _13387 = _12301 < _13386;
  wire _13388 = r1927 ^ _13387;
  wire _13389 = _12298 ? coded_block[1927] : r1927;
  wire _13390 = _12296 ? _13388 : _13389;
  always @ (posedge reset or posedge clock) if (reset) r1927 <= 1'd0; else if (_12300) r1927 <= _13390;
  wire [1:0] _13391 = {_0, _1662} + {_0, _2175};
  wire [1:0] _13392 = {_0, _5884} + {_0, _8155};
  wire [2:0] _13393 = {_0, _13391} + {_0, _13392};
  wire [1:0] _13394 = {_0, _10077} + {_0, _10462};
  wire [3:0] _13395 = {_0, _13393} + {_0, _0, _13394};
  wire _13396 = _12301 < _13395;
  wire _13397 = r1926 ^ _13396;
  wire _13398 = _12298 ? coded_block[1926] : r1926;
  wire _13399 = _12296 ? _13397 : _13398;
  always @ (posedge reset or posedge clock) if (reset) r1926 <= 1'd0; else if (_12300) r1926 <= _13399;
  wire [1:0] _13400 = {_0, _510} + {_0, _2910};
  wire [1:0] _13401 = {_0, _4830} + {_0, _7230};
  wire [2:0] _13402 = {_0, _13400} + {_0, _13401};
  wire [1:0] _13403 = {_0, _10014} + {_0, _10654};
  wire [3:0] _13404 = {_0, _13402} + {_0, _0, _13403};
  wire _13405 = _12301 < _13404;
  wire _13406 = r1925 ^ _13405;
  wire _13407 = _12298 ? coded_block[1925] : r1925;
  wire _13408 = _12296 ? _13406 : _13407;
  always @ (posedge reset or posedge clock) if (reset) r1925 <= 1'd0; else if (_12300) r1925 <= _13408;
  wire [1:0] _13409 = {_0, _289} + {_0, _3805};
  wire [1:0] _13410 = {_0, _5470} + {_0, _6525};
  wire [2:0] _13411 = {_0, _13409} + {_0, _13410};
  wire [1:0] _13412 = {_0, _8991} + {_0, _11516};
  wire [3:0] _13413 = {_0, _13411} + {_0, _0, _13412};
  wire _13414 = _12301 < _13413;
  wire _13415 = r1924 ^ _13414;
  wire _13416 = _12298 ? coded_block[1924] : r1924;
  wire _13417 = _12296 ? _13415 : _13416;
  always @ (posedge reset or posedge clock) if (reset) r1924 <= 1'd0; else if (_12300) r1924 <= _13417;
  wire [1:0] _13418 = {_0, _1533} + {_0, _2910};
  wire [1:0] _13419 = {_0, _5215} + {_0, _8155};
  wire [2:0] _13420 = {_0, _13418} + {_0, _13419};
  wire [1:0] _13421 = {_0, _9853} + {_0, _12124};
  wire [3:0] _13422 = {_0, _13420} + {_0, _0, _13421};
  wire _13423 = _12301 < _13422;
  wire _13424 = r1923 ^ _13423;
  wire _13425 = _12298 ? coded_block[1923] : r1923;
  wire _13426 = _12296 ? _13424 : _13425;
  always @ (posedge reset or posedge clock) if (reset) r1923 <= 1'd0; else if (_12300) r1923 <= _13426;
  wire [1:0] _13427 = {_0, _958} + {_0, _2686};
  wire [1:0] _13428 = {_0, _5501} + {_0, _6718};
  wire [2:0] _13429 = {_0, _13427} + {_0, _13428};
  wire [1:0] _13430 = {_0, _8288} + {_0, _10462};
  wire [3:0] _13431 = {_0, _13429} + {_0, _0, _13430};
  wire _13432 = _12301 < _13431;
  wire _13433 = r1922 ^ _13432;
  wire _13434 = _12298 ? coded_block[1922] : r1922;
  wire _13435 = _12296 ? _13433 : _13434;
  always @ (posedge reset or posedge clock) if (reset) r1922 <= 1'd0; else if (_12300) r1922 <= _13435;
  wire [1:0] _13436 = {_0, _1021} + {_0, _2367};
  wire [1:0] _13437 = {_0, _5022} + {_0, _6621};
  wire [2:0] _13438 = {_0, _13436} + {_0, _13437};
  wire [1:0] _13439 = {_0, _8288} + {_0, _11358};
  wire [3:0] _13440 = {_0, _13438} + {_0, _0, _13439};
  wire _13441 = _12301 < _13440;
  wire _13442 = r1921 ^ _13441;
  wire _13443 = _12298 ? coded_block[1921] : r1921;
  wire _13444 = _12296 ? _13442 : _13443;
  always @ (posedge reset or posedge clock) if (reset) r1921 <= 1'd0; else if (_12300) r1921 <= _13444;
  wire [1:0] _13445 = {_0, _1917} + {_0, _2367};
  wire [1:0] _13446 = {_0, _5726} + {_0, _7454};
  wire [2:0] _13447 = {_0, _13445} + {_0, _13446};
  wire [1:0] _13448 = {_0, _9661} + {_0, _11516};
  wire [3:0] _13449 = {_0, _13447} + {_0, _0, _13448};
  wire _13450 = _12301 < _13449;
  wire _13451 = r1920 ^ _13450;
  wire _13452 = _12298 ? coded_block[1920] : r1920;
  wire _13453 = _12296 ? _13451 : _13452;
  always @ (posedge reset or posedge clock) if (reset) r1920 <= 1'd0; else if (_12300) r1920 <= _13453;
  wire [1:0] _13454 = {_0, _128} + {_0, _2686};
  wire [1:0] _13455 = {_0, _5215} + {_0, _6687};
  wire [2:0] _13456 = {_0, _13454} + {_0, _13455};
  wire [1:0] _13457 = {_0, _10045} + {_0, _11771};
  wire [3:0] _13458 = {_0, _13456} + {_0, _0, _13457};
  wire _13459 = _12301 < _13458;
  wire _13460 = r1919 ^ _13459;
  wire _13461 = _12298 ? coded_block[1919] : r1919;
  wire _13462 = _12296 ? _13460 : _13461;
  always @ (posedge reset or posedge clock) if (reset) r1919 <= 1'd0; else if (_12300) r1919 <= _13462;
  wire [1:0] _13463 = {_0, _352} + {_0, _2878};
  wire [1:0] _13464 = {_0, _4574} + {_0, _6845};
  wire [2:0] _13465 = {_0, _13463} + {_0, _13464};
  wire [1:0] _13466 = {_0, _8767} + {_0, _11165};
  wire [3:0] _13467 = {_0, _13465} + {_0, _0, _13466};
  wire _13468 = _12301 < _13467;
  wire _13469 = r1918 ^ _13468;
  wire _13470 = _12298 ? coded_block[1918] : r1918;
  wire _13471 = _12296 ? _13469 : _13470;
  always @ (posedge reset or posedge clock) if (reset) r1918 <= 1'd0; else if (_12300) r1918 <= _13471;
  wire [1:0] _13472 = {_0, _1726} + {_0, _2813};
  wire [1:0] _13473 = {_0, _5310} + {_0, _6718};
  wire [2:0] _13474 = {_0, _13472} + {_0, _13473};
  wire [1:0] _13475 = {_0, _9693} + {_0, _11837};
  wire [3:0] _13476 = {_0, _13474} + {_0, _0, _13475};
  wire _13477 = _12301 < _13476;
  wire _13478 = r1917 ^ _13477;
  wire _13479 = _12298 ? coded_block[1917] : r1917;
  wire _13480 = _12296 ? _13478 : _13479;
  always @ (posedge reset or posedge clock) if (reset) r1917 <= 1'd0; else if (_12300) r1917 <= _13480;
  wire [1:0] _13481 = {_0, _1695} + {_0, _2782};
  wire [1:0] _13482 = {_0, _5279} + {_0, _6687};
  wire [2:0] _13483 = {_0, _13481} + {_0, _13482};
  wire [1:0] _13484 = {_0, _9661} + {_0, _11806};
  wire [3:0] _13485 = {_0, _13483} + {_0, _0, _13484};
  wire _13486 = _12301 < _13485;
  wire _13487 = r1916 ^ _13486;
  wire _13488 = _12298 ? coded_block[1916] : r1916;
  wire _13489 = _12296 ? _13487 : _13488;
  always @ (posedge reset or posedge clock) if (reset) r1916 <= 1'd0; else if (_12300) r1916 <= _13489;
  wire [1:0] _13490 = {_0, _1247} + {_0, _2592};
  wire [1:0] _13491 = {_0, _5246} + {_0, _6845};
  wire [2:0] _13492 = {_0, _13490} + {_0, _13491};
  wire [1:0] _13493 = {_0, _8511} + {_0, _11581};
  wire [3:0] _13494 = {_0, _13492} + {_0, _0, _13493};
  wire _13495 = _12301 < _13494;
  wire _13496 = r1915 ^ _13495;
  wire _13497 = _12298 ? coded_block[1915] : r1915;
  wire _13498 = _12296 ? _13496 : _13497;
  always @ (posedge reset or posedge clock) if (reset) r1915 <= 1'd0; else if (_12300) r1915 <= _13498;
  wire [1:0] _13499 = {_0, _383} + {_0, _2367};
  wire [1:0] _13500 = {_0, _5279} + {_0, _6589};
  wire [2:0] _13501 = {_0, _13499} + {_0, _13500};
  wire [1:0] _13502 = {_0, _9693} + {_0, _12282};
  wire [3:0] _13503 = {_0, _13501} + {_0, _0, _13502};
  wire _13504 = _12301 < _13503;
  wire _13505 = r1914 ^ _13504;
  wire _13506 = _12298 ? coded_block[1914] : r1914;
  wire _13507 = _12296 ? _13505 : _13506;
  always @ (posedge reset or posedge clock) if (reset) r1914 <= 1'd0; else if (_12300) r1914 <= _13507;
  wire [1:0] _13508 = {_0, _958} + {_0, _3773};
  wire [1:0] _13509 = {_0, _5022} + {_0, _7132};
  wire [2:0] _13510 = {_0, _13508} + {_0, _13509};
  wire [1:0] _13511 = {_0, _9980} + {_0, _10717};
  wire [3:0] _13512 = {_0, _13510} + {_0, _0, _13511};
  wire _13513 = _12301 < _13512;
  wire _13514 = r1913 ^ _13513;
  wire _13515 = _12298 ? coded_block[1913] : r1913;
  wire _13516 = _12296 ? _13514 : _13515;
  always @ (posedge reset or posedge clock) if (reset) r1913 <= 1'd0; else if (_12300) r1913 <= _13516;
  wire [1:0] _13517 = {_0, _1312} + {_0, _3262};
  wire [1:0] _13518 = {_0, _4861} + {_0, _6525};
  wire [2:0] _13519 = {_0, _13517} + {_0, _13518};
  wire [1:0] _13520 = {_0, _9597} + {_0, _12061};
  wire [3:0] _13521 = {_0, _13519} + {_0, _0, _13520};
  wire _13522 = _12301 < _13521;
  wire _13523 = r1912 ^ _13522;
  wire _13524 = _12298 ? coded_block[1912] : r1912;
  wire _13525 = _12296 ? _13523 : _13524;
  always @ (posedge reset or posedge clock) if (reset) r1912 <= 1'd0; else if (_12300) r1912 <= _13525;
  wire [1:0] _13526 = {_0, _1568} + {_0, _2847};
  wire [1:0] _13527 = {_0, _4830} + {_0, _7996};
  wire [2:0] _13528 = {_0, _13526} + {_0, _13527};
  wire [1:0] _13529 = {_0, _8701} + {_0, _10335};
  wire [3:0] _13530 = {_0, _13528} + {_0, _0, _13529};
  wire _13531 = _12301 < _13530;
  wire _13532 = r1911 ^ _13531;
  wire _13533 = _12298 ? coded_block[1911] : r1911;
  wire _13534 = _12296 ? _13532 : _13533;
  always @ (posedge reset or posedge clock) if (reset) r1911 <= 1'd0; else if (_12300) r1911 <= _13534;
  wire [1:0] _13535 = {_0, _510} + {_0, _3997};
  wire [1:0] _13536 = {_0, _4542} + {_0, _7454};
  wire [2:0] _13537 = {_0, _13535} + {_0, _13536};
  wire [1:0] _13538 = {_0, _8767} + {_0, _11869};
  wire [3:0] _13539 = {_0, _13537} + {_0, _0, _13538};
  wire _13540 = _12301 < _13539;
  wire _13541 = r1910 ^ _13540;
  wire _13542 = _12298 ? coded_block[1910] : r1910;
  wire _13543 = _12296 ? _13541 : _13542;
  always @ (posedge reset or posedge clock) if (reset) r1910 <= 1'd0; else if (_12300) r1910 <= _13543;
  wire [1:0] _13544 = {_0, _1247} + {_0, _2750};
  wire [1:0] _13545 = {_0, _4415} + {_0, _7485};
  wire [2:0] _13546 = {_0, _13544} + {_0, _13545};
  wire [1:0] _13547 = {_0, _9949} + {_0, _10462};
  wire [3:0] _13548 = {_0, _13546} + {_0, _0, _13547};
  wire _13549 = _12301 < _13548;
  wire _13550 = r1909 ^ _13549;
  wire _13551 = _12298 ? coded_block[1909] : r1909;
  wire _13552 = _12296 ? _13550 : _13551;
  always @ (posedge reset or posedge clock) if (reset) r1909 <= 1'd0; else if (_12300) r1909 <= _13552;
  wire [1:0] _13553 = {_0, _1695} + {_0, _3104};
  wire [1:0] _13554 = {_0, _5534} + {_0, _6718};
  wire [2:0] _13555 = {_0, _13553} + {_0, _13554};
  wire [1:0] _13556 = {_0, _8543} + {_0, _11165};
  wire [3:0] _13557 = {_0, _13555} + {_0, _0, _13556};
  wire _13558 = _12301 < _13557;
  wire _13559 = r1908 ^ _13558;
  wire _13560 = _12298 ? coded_block[1908] : r1908;
  wire _13561 = _12296 ? _13559 : _13560;
  always @ (posedge reset or posedge clock) if (reset) r1908 <= 1'd0; else if (_12300) r1908 <= _13561;
  wire [1:0] _13562 = {_0, _161} + {_0, _2719};
  wire [1:0] _13563 = {_0, _5246} + {_0, _6718};
  wire [2:0] _13564 = {_0, _13562} + {_0, _13563};
  wire [1:0] _13565 = {_0, _10077} + {_0, _11806};
  wire [3:0] _13566 = {_0, _13564} + {_0, _0, _13565};
  wire _13567 = _12301 < _13566;
  wire _13568 = r1907 ^ _13567;
  wire _13569 = _12298 ? coded_block[1907] : r1907;
  wire _13570 = _12296 ? _13568 : _13569;
  always @ (posedge reset or posedge clock) if (reset) r1907 <= 1'd0; else if (_12300) r1907 <= _13570;
  wire [1:0] _13571 = {_0, _1406} + {_0, _3294};
  wire [1:0] _13572 = {_0, _5310} + {_0, _8186};
  wire [2:0] _13573 = {_0, _13571} + {_0, _13572};
  wire [1:0] _13574 = {_0, _8511} + {_0, _11964};
  wire [3:0] _13575 = {_0, _13573} + {_0, _0, _13574};
  wire _13576 = _12301 < _13575;
  wire _13577 = r1906 ^ _13576;
  wire _13578 = _12298 ? coded_block[1906] : r1906;
  wire _13579 = _12296 ? _13577 : _13578;
  always @ (posedge reset or posedge clock) if (reset) r1906 <= 1'd0; else if (_12300) r1906 <= _13579;
  wire [1:0] _13580 = {_0, _1726} + {_0, _2941};
  wire [1:0] _13581 = {_0, _6108} + {_0, _6814};
  wire [2:0] _13582 = {_0, _13580} + {_0, _13581};
  wire [1:0] _13583 = {_0, _8446} + {_0, _12219};
  wire [3:0] _13584 = {_0, _13582} + {_0, _0, _13583};
  wire _13585 = _12301 < _13584;
  wire _13586 = r1905 ^ _13585;
  wire _13587 = _12298 ? coded_block[1905] : r1905;
  wire _13588 = _12296 ? _13586 : _13587;
  always @ (posedge reset or posedge clock) if (reset) r1905 <= 1'd0; else if (_12300) r1905 <= _13588;
  wire [1:0] _13589 = {_0, _97} + {_0, _3870};
  wire [1:0] _13590 = {_0, _5597} + {_0, _7804};
  wire [2:0] _13591 = {_0, _13589} + {_0, _13590};
  wire [1:0] _13592 = {_0, _9661} + {_0, _12092};
  wire [3:0] _13593 = {_0, _13591} + {_0, _0, _13592};
  wire _13594 = _12301 < _13593;
  wire _13595 = r1904 ^ _13594;
  wire _13596 = _12298 ? coded_block[1904] : r1904;
  wire _13597 = _12296 ? _13595 : _13596;
  always @ (posedge reset or posedge clock) if (reset) r1904 <= 1'd0; else if (_12300) r1904 <= _13597;
  wire [1:0] _13598 = {_0, _735} + {_0, _2847};
  wire [1:0] _13599 = {_0, _5949} + {_0, _6525};
  wire [2:0] _13600 = {_0, _13598} + {_0, _13599};
  wire [1:0] _13601 = {_0, _9661} + {_0, _12027};
  wire [3:0] _13602 = {_0, _13600} + {_0, _0, _13601};
  wire _13603 = _12301 < _13602;
  wire _13604 = r1903 ^ _13603;
  wire _13605 = _12298 ? coded_block[1903] : r1903;
  wire _13606 = _12296 ? _13604 : _13605;
  always @ (posedge reset or posedge clock) if (reset) r1903 <= 1'd0; else if (_12300) r1903 <= _13606;
  wire [1:0] _13607 = {_0, _289} + {_0, _2081};
  wire [1:0] _13608 = {_0, _4574} + {_0, _6814};
  wire [2:0] _13609 = {_0, _13607} + {_0, _13608};
  wire [1:0] _13610 = {_0, _9503} + {_0, _11295};
  wire [3:0] _13611 = {_0, _13609} + {_0, _0, _13610};
  wire _13612 = _12301 < _13611;
  wire _13613 = r1902 ^ _13612;
  wire _13614 = _12298 ? coded_block[1902] : r1902;
  wire _13615 = _12296 ? _13613 : _13614;
  always @ (posedge reset or posedge clock) if (reset) r1902 <= 1'd0; else if (_12300) r1902 <= _13615;
  wire [1:0] _13616 = {_0, _161} + {_0, _3037};
  wire [1:0] _13617 = {_0, _5790} + {_0, _7741};
  wire [2:0] _13618 = {_0, _13616} + {_0, _13617};
  wire [1:0] _13619 = {_0, _8288} + {_0, _11196};
  wire [3:0] _13620 = {_0, _13618} + {_0, _0, _13619};
  wire _13621 = _12301 < _13620;
  wire _13622 = r1901 ^ _13621;
  wire _13623 = _12298 ? coded_block[1901] : r1901;
  wire _13624 = _12296 ? _13622 : _13623;
  always @ (posedge reset or posedge clock) if (reset) r1901 <= 1'd0; else if (_12300) r1901 <= _13624;
  wire [1:0] _13625 = {_0, _545} + {_0, _2175};
  wire [1:0] _13626 = {_0, _5116} + {_0, _6814};
  wire [2:0] _13627 = {_0, _13625} + {_0, _13626};
  wire [1:0] _13628 = {_0, _9085} + {_0, _11004};
  wire [3:0] _13629 = {_0, _13627} + {_0, _0, _13628};
  wire _13630 = _12301 < _13629;
  wire _13631 = r1900 ^ _13630;
  wire _13632 = _12298 ? coded_block[1900] : r1900;
  wire _13633 = _12296 ? _13631 : _13632;
  always @ (posedge reset or posedge clock) if (reset) r1900 <= 1'd0; else if (_12300) r1900 <= _13633;
  wire [1:0] _13634 = {_0, _1533} + {_0, _3870};
  wire [1:0] _13635 = {_0, _4574} + {_0, _6207};
  wire [2:0] _13636 = {_0, _13634} + {_0, _13635};
  wire [1:0] _13637 = {_0, _9980} + {_0, _10973};
  wire [3:0] _13638 = {_0, _13636} + {_0, _0, _13637};
  wire _13639 = _12301 < _13638;
  wire _13640 = r1899 ^ _13639;
  wire _13641 = _12298 ? coded_block[1899] : r1899;
  wire _13642 = _12296 ? _13640 : _13641;
  always @ (posedge reset or posedge clock) if (reset) r1899 <= 1'd0; else if (_12300) r1899 <= _13642;
  wire [1:0] _13643 = {_0, _958} + {_0, _3997};
  wire [1:0] _13644 = {_0, _5470} + {_0, _6814};
  wire [2:0] _13645 = {_0, _13643} + {_0, _13644};
  wire [1:0] _13646 = {_0, _8543} + {_0, _10748};
  wire [3:0] _13647 = {_0, _13645} + {_0, _0, _13646};
  wire _13648 = _12301 < _13647;
  wire _13649 = r1898 ^ _13648;
  wire _13650 = _12298 ? coded_block[1898] : r1898;
  wire _13651 = _12296 ? _13649 : _13650;
  always @ (posedge reset or posedge clock) if (reset) r1898 <= 1'd0; else if (_12300) r1898 <= _13651;
  wire [1:0] _13652 = {_0, _1247} + {_0, _2719};
  wire [1:0] _13653 = {_0, _5279} + {_0, _8186};
  wire [2:0] _13654 = {_0, _13652} + {_0, _13653};
  wire [1:0] _13655 = {_0, _9503} + {_0, _10590};
  wire [3:0] _13656 = {_0, _13654} + {_0, _0, _13655};
  wire _13657 = _12301 < _13656;
  wire _13658 = r1897 ^ _13657;
  wire _13659 = _12298 ? coded_block[1897] : r1897;
  wire _13660 = _12296 ? _13658 : _13659;
  always @ (posedge reset or posedge clock) if (reset) r1897 <= 1'd0; else if (_12300) r1897 <= _13660;
  wire [1:0] _13661 = {_0, _1533} + {_0, _4028};
  wire [1:0] _13662 = {_0, _5246} + {_0, _6814};
  wire [2:0] _13663 = {_0, _13661} + {_0, _13662};
  wire [1:0] _13664 = {_0, _8991} + {_0, _10366};
  wire [3:0] _13665 = {_0, _13663} + {_0, _0, _13664};
  wire _13666 = _12301 < _13665;
  wire _13667 = r1896 ^ _13666;
  wire _13668 = _12298 ? coded_block[1896] : r1896;
  wire _13669 = _12296 ? _13667 : _13668;
  always @ (posedge reset or posedge clock) if (reset) r1896 <= 1'd0; else if (_12300) r1896 <= _13669;
  wire [1:0] _13670 = {_0, _352} + {_0, _3037};
  wire [1:0] _13671 = {_0, _5373} + {_0, _6814};
  wire [2:0] _13672 = {_0, _13670} + {_0, _13671};
  wire [1:0] _13673 = {_0, _8701} + {_0, _10272};
  wire [3:0] _13674 = {_0, _13672} + {_0, _0, _13673};
  wire _13675 = _12301 < _13674;
  wire _13676 = r1895 ^ _13675;
  wire _13677 = _12298 ? coded_block[1895] : r1895;
  wire _13678 = _12296 ? _13676 : _13677;
  always @ (posedge reset or posedge clock) if (reset) r1895 <= 1'd0; else if (_12300) r1895 <= _13678;
  wire [1:0] _13679 = {_0, _958} + {_0, _2878};
  wire [1:0] _13680 = {_0, _4384} + {_0, _6687};
  wire [2:0] _13681 = {_0, _13679} + {_0, _13680};
  wire [1:0] _13682 = {_0, _9630} + {_0, _11326};
  wire [3:0] _13683 = {_0, _13681} + {_0, _0, _13682};
  wire _13684 = _12301 < _13683;
  wire _13685 = r1894 ^ _13684;
  wire _13686 = _12298 ? coded_block[1894] : r1894;
  wire _13687 = _12296 ? _13685 : _13686;
  always @ (posedge reset or posedge clock) if (reset) r1894 <= 1'd0; else if (_12300) r1894 <= _13687;
  wire [1:0] _13688 = {_0, _1533} + {_0, _3517};
  wire [1:0] _13689 = {_0, _4415} + {_0, _7741};
  wire [2:0] _13690 = {_0, _13688} + {_0, _13689};
  wire [1:0] _13691 = {_0, _8830} + {_0, _11422};
  wire [3:0] _13692 = {_0, _13690} + {_0, _0, _13691};
  wire _13693 = _12301 < _13692;
  wire _13694 = r1893 ^ _13693;
  wire _13695 = _12298 ? coded_block[1893] : r1893;
  wire _13696 = _12296 ? _13694 : _13695;
  always @ (posedge reset or posedge clock) if (reset) r1893 <= 1'd0; else if (_12300) r1893 <= _13696;
  wire [1:0] _13697 = {_0, _161} + {_0, _2878};
  wire [1:0] _13698 = {_0, _5501} + {_0, _7485};
  wire [2:0] _13699 = {_0, _13697} + {_0, _13698};
  wire [1:0] _13700 = {_0, _8638} + {_0, _11358};
  wire [3:0] _13701 = {_0, _13699} + {_0, _0, _13700};
  wire _13702 = _12301 < _13701;
  wire _13703 = r1892 ^ _13702;
  wire _13704 = _12298 ? coded_block[1892] : r1892;
  wire _13705 = _12296 ? _13703 : _13704;
  always @ (posedge reset or posedge clock) if (reset) r1892 <= 1'd0; else if (_12300) r1892 <= _13705;
  wire [1:0] _13706 = {_0, _289} + {_0, _2557};
  wire [1:0] _13707 = {_0, _4958} + {_0, _7741};
  wire [2:0] _13708 = {_0, _13706} + {_0, _13707};
  wire [1:0] _13709 = {_0, _8383} + {_0, _11996};
  wire [3:0] _13710 = {_0, _13708} + {_0, _0, _13709};
  wire _13711 = _12301 < _13710;
  wire _13712 = r1891 ^ _13711;
  wire _13713 = _12298 ? coded_block[1891] : r1891;
  wire _13714 = _12296 ? _13712 : _13713;
  always @ (posedge reset or posedge clock) if (reset) r1891 <= 1'd0; else if (_12300) r1891 <= _13714;
  wire [1:0] _13715 = {_0, _1758} + {_0, _3294};
  wire [1:0] _13716 = {_0, _4703} + {_0, _7675};
  wire [2:0] _13717 = {_0, _13715} + {_0, _13716};
  wire [1:0] _13718 = {_0, _9822} + {_0, _11326};
  wire [3:0] _13719 = {_0, _13717} + {_0, _0, _13718};
  wire _13720 = _12301 < _13719;
  wire _13721 = r1890 ^ _13720;
  wire _13722 = _12298 ? coded_block[1890] : r1890;
  wire _13723 = _12296 ? _13721 : _13722;
  always @ (posedge reset or posedge clock) if (reset) r1890 <= 1'd0; else if (_12300) r1890 <= _13723;
  wire [1:0] _13724 = {_0, _1406} + {_0, _3453};
  wire [1:0] _13725 = {_0, _5501} + {_0, _7548};
  wire [2:0] _13726 = {_0, _13724} + {_0, _13725};
  wire [1:0] _13727 = {_0, _9597} + {_0, _11644};
  wire [3:0] _13728 = {_0, _13726} + {_0, _0, _13727};
  wire _13729 = _12301 < _13728;
  wire _13730 = r1889 ^ _13729;
  wire _13731 = _12298 ? coded_block[1889] : r1889;
  wire _13732 = _12296 ? _13730 : _13731;
  always @ (posedge reset or posedge clock) if (reset) r1889 <= 1'd0; else if (_12300) r1889 <= _13732;
  wire [1:0] _13733 = {_0, _1184} + {_0, _2910};
  wire [1:0] _13734 = {_0, _5726} + {_0, _6942};
  wire [2:0] _13735 = {_0, _13733} + {_0, _13734};
  wire [1:0] _13736 = {_0, _8511} + {_0, _10685};
  wire [3:0] _13737 = {_0, _13735} + {_0, _0, _13736};
  wire _13738 = _12301 < _13737;
  wire _13739 = r1888 ^ _13738;
  wire _13740 = _12298 ? coded_block[1888] : r1888;
  wire _13741 = _12296 ? _13739 : _13740;
  always @ (posedge reset or posedge clock) if (reset) r1888 <= 1'd0; else if (_12300) r1888 <= _13741;
  wire [1:0] _13742 = {_0, _1568} + {_0, _3037};
  wire [1:0] _13743 = {_0, _5597} + {_0, _6494};
  wire [2:0] _13744 = {_0, _13742} + {_0, _13743};
  wire [1:0] _13745 = {_0, _9822} + {_0, _10910};
  wire [3:0] _13746 = {_0, _13744} + {_0, _0, _13745};
  wire _13747 = _12301 < _13746;
  wire _13748 = r1887 ^ _13747;
  wire _13749 = _12298 ? coded_block[1887] : r1887;
  wire _13750 = _12296 ? _13748 : _13749;
  always @ (posedge reset or posedge clock) if (reset) r1887 <= 1'd0; else if (_12300) r1887 <= _13750;
  wire [1:0] _13751 = {_0, _289} + {_0, _3104};
  wire [1:0] _13752 = {_0, _4350} + {_0, _6462};
  wire [2:0] _13753 = {_0, _13751} + {_0, _13752};
  wire [1:0] _13754 = {_0, _9311} + {_0, _12061};
  wire [3:0] _13755 = {_0, _13753} + {_0, _0, _13754};
  wire _13756 = _12301 < _13755;
  wire _13757 = r1886 ^ _13756;
  wire _13758 = _12298 ? coded_block[1886] : r1886;
  wire _13759 = _12296 ? _13757 : _13758;
  always @ (posedge reset or posedge clock) if (reset) r1886 <= 1'd0; else if (_12300) r1886 <= _13759;
  wire [1:0] _13760 = {_0, _639} + {_0, _3422};
  wire [1:0] _13761 = {_0, _5790} + {_0, _6270};
  wire [2:0] _13762 = {_0, _13760} + {_0, _13761};
  wire [1:0] _13763 = {_0, _9693} + {_0, _10654};
  wire [3:0] _13764 = {_0, _13762} + {_0, _0, _13763};
  wire _13765 = _12301 < _13764;
  wire _13766 = r1885 ^ _13765;
  wire _13767 = _12298 ? coded_block[1885] : r1885;
  wire _13768 = _12296 ? _13766 : _13767;
  always @ (posedge reset or posedge clock) if (reset) r1885 <= 1'd0; else if (_12300) r1885 <= _13768;
  wire [1:0] _13769 = {_0, _639} + {_0, _3262};
  wire [1:0] _13770 = {_0, _6045} + {_0, _6687};
  wire [2:0] _13771 = {_0, _13769} + {_0, _13770};
  wire [1:0] _13772 = {_0, _8288} + {_0, _11964};
  wire [3:0] _13773 = {_0, _13771} + {_0, _0, _13772};
  wire _13774 = _12301 < _13773;
  wire _13775 = r1884 ^ _13774;
  wire _13776 = _12298 ? coded_block[1884] : r1884;
  wire _13777 = _12296 ? _13775 : _13776;
  always @ (posedge reset or posedge clock) if (reset) r1884 <= 1'd0; else if (_12300) r1884 <= _13777;
  wire [1:0] _13778 = {_0, _1950} + {_0, _2557};
  wire [1:0] _13779 = {_0, _5342} + {_0, _7996};
  wire [2:0] _13780 = {_0, _13778} + {_0, _13779};
  wire [1:0] _13781 = {_0, _9597} + {_0, _11259};
  wire [3:0] _13782 = {_0, _13780} + {_0, _0, _13781};
  wire _13783 = _12301 < _13782;
  wire _13784 = r1883 ^ _13783;
  wire _13785 = _12298 ? coded_block[1883] : r1883;
  wire _13786 = _12296 ? _13784 : _13785;
  always @ (posedge reset or posedge clock) if (reset) r1883 <= 1'd0; else if (_12300) r1883 <= _13786;
  wire [1:0] _13787 = {_0, _735} + {_0, _2910};
  wire [1:0] _13788 = {_0, _5183} + {_0, _7100};
  wire [2:0] _13789 = {_0, _13787} + {_0, _13788};
  wire [1:0] _13790 = {_0, _9503} + {_0, _12282};
  wire [3:0] _13791 = {_0, _13789} + {_0, _0, _13790};
  wire _13792 = _12301 < _13791;
  wire _13793 = r1882 ^ _13792;
  wire _13794 = _12298 ? coded_block[1882] : r1882;
  wire _13795 = _12296 ? _13793 : _13794;
  always @ (posedge reset or posedge clock) if (reset) r1882 <= 1'd0; else if (_12300) r1882 <= _13795;
  wire [1:0] _13796 = {_0, _1247} + {_0, _2910};
  wire [1:0] _13797 = {_0, _4478} + {_0, _6652};
  wire [2:0] _13798 = {_0, _13796} + {_0, _13797};
  wire [1:0] _13799 = {_0, _10045} + {_0, _11326};
  wire [3:0] _13800 = {_0, _13798} + {_0, _0, _13799};
  wire _13801 = _12301 < _13800;
  wire _13802 = r1881 ^ _13801;
  wire _13803 = _12298 ? coded_block[1881] : r1881;
  wire _13804 = _12296 ? _13802 : _13803;
  always @ (posedge reset or posedge clock) if (reset) r1881 <= 1'd0; else if (_12300) r1881 <= _13804;
  wire [1:0] _13805 = {_0, _2013} + {_0, _2399};
  wire [1:0] _13806 = {_0, _4319} + {_0, _6718};
  wire [2:0] _13807 = {_0, _13805} + {_0, _13806};
  wire [1:0] _13808 = {_0, _9503} + {_0, _12155};
  wire [3:0] _13809 = {_0, _13807} + {_0, _0, _13808};
  wire _13810 = _12301 < _13809;
  wire _13811 = r1880 ^ _13810;
  wire _13812 = _12298 ? coded_block[1880] : r1880;
  wire _13813 = _12296 ? _13811 : _13812;
  always @ (posedge reset or posedge clock) if (reset) r1880 <= 1'd0; else if (_12300) r1880 <= _13813;
  wire [1:0] _13814 = {_0, _1502} + {_0, _3836};
  wire [1:0] _13815 = {_0, _4542} + {_0, _8186};
  wire [2:0] _13816 = {_0, _13814} + {_0, _13815};
  wire [1:0] _13817 = {_0, _9949} + {_0, _10941};
  wire [3:0] _13818 = {_0, _13816} + {_0, _0, _13817};
  wire _13819 = _12301 < _13818;
  wire _13820 = r1879 ^ _13819;
  wire _13821 = _12298 ? coded_block[1879] : r1879;
  wire _13822 = _12296 ? _13820 : _13821;
  always @ (posedge reset or posedge clock) if (reset) r1879 <= 1'd0; else if (_12300) r1879 <= _13822;
  wire [1:0] _13823 = {_0, _1120} + {_0, _2623};
  wire [1:0] _13824 = {_0, _4287} + {_0, _7357};
  wire [2:0] _13825 = {_0, _13823} + {_0, _13824};
  wire [1:0] _13826 = {_0, _9822} + {_0, _10335};
  wire [3:0] _13827 = {_0, _13825} + {_0, _0, _13826};
  wire _13828 = _12301 < _13827;
  wire _13829 = r1878 ^ _13828;
  wire _13830 = _12298 ? coded_block[1878] : r1878;
  wire _13831 = _12296 ? _13829 : _13830;
  always @ (posedge reset or posedge clock) if (reset) r1878 <= 1'd0; else if (_12300) r1878 <= _13831;
  wire [1:0] _13832 = {_0, _831} + {_0, _3773};
  wire [1:0] _13833 = {_0, _5597} + {_0, _6207};
  wire [2:0] _13834 = {_0, _13832} + {_0, _13833};
  wire [1:0] _13835 = {_0, _10204} + {_0, _11358};
  wire [3:0] _13836 = {_0, _13834} + {_0, _0, _13835};
  wire _13837 = _12301 < _13836;
  wire _13838 = r1877 ^ _13837;
  wire _13839 = _12298 ? coded_block[1877] : r1877;
  wire _13840 = _12296 ? _13838 : _13839;
  always @ (posedge reset or posedge clock) if (reset) r1877 <= 1'd0; else if (_12300) r1877 <= _13840;
  wire [1:0] _13841 = {_0, _672} + {_0, _3964};
  wire [1:0] _13842 = {_0, _5949} + {_0, _7100};
  wire [2:0] _13843 = {_0, _13841} + {_0, _13842};
  wire [1:0] _13844 = {_0, _9822} + {_0, _11453};
  wire [3:0] _13845 = {_0, _13843} + {_0, _0, _13844};
  wire _13846 = _12301 < _13845;
  wire _13847 = r1876 ^ _13846;
  wire _13848 = _12298 ? coded_block[1876] : r1876;
  wire _13849 = _12296 ? _13847 : _13848;
  always @ (posedge reset or posedge clock) if (reset) r1876 <= 1'd0; else if (_12300) r1876 <= _13849;
  wire [1:0] _13850 = {_0, _831} + {_0, _2144};
  wire [1:0] _13851 = {_0, _5534} + {_0, _6814};
  wire [2:0] _13852 = {_0, _13850} + {_0, _13851};
  wire [1:0] _13853 = {_0, _8830} + {_0, _11708};
  wire [3:0] _13854 = {_0, _13852} + {_0, _0, _13853};
  wire _13855 = _12301 < _13854;
  wire _13856 = r1875 ^ _13855;
  wire _13857 = _12298 ? coded_block[1875] : r1875;
  wire _13858 = _12296 ? _13856 : _13857;
  always @ (posedge reset or posedge clock) if (reset) r1875 <= 1'd0; else if (_12300) r1875 <= _13858;
  wire [1:0] _13859 = {_0, _1917} + {_0, _2623};
  wire [1:0] _13860 = {_0, _5246} + {_0, _7230};
  wire [2:0] _13861 = {_0, _13859} + {_0, _13860};
  wire [1:0] _13862 = {_0, _8383} + {_0, _11101};
  wire [3:0] _13863 = {_0, _13861} + {_0, _0, _13862};
  wire _13864 = _12301 < _13863;
  wire _13865 = r1874 ^ _13864;
  wire _13866 = _12298 ? coded_block[1874] : r1874;
  wire _13867 = _12296 ? _13865 : _13866;
  always @ (posedge reset or posedge clock) if (reset) r1874 <= 1'd0; else if (_12300) r1874 <= _13867;
  wire [1:0] _13868 = {_0, _1184} + {_0, _3805};
  wire [1:0] _13869 = {_0, _4574} + {_0, _7230};
  wire [2:0] _13870 = {_0, _13868} + {_0, _13869};
  wire [1:0] _13871 = {_0, _8830} + {_0, _10493};
  wire [3:0] _13872 = {_0, _13870} + {_0, _0, _13871};
  wire _13873 = _12301 < _13872;
  wire _13874 = r1873 ^ _13873;
  wire _13875 = _12298 ? coded_block[1873] : r1873;
  wire _13876 = _12296 ? _13874 : _13875;
  always @ (posedge reset or posedge clock) if (reset) r1873 <= 1'd0; else if (_12300) r1873 <= _13876;
  wire [1:0] _13877 = {_0, _1695} + {_0, _2750};
  wire [1:0] _13878 = {_0, _4542} + {_0, _7804};
  wire [2:0] _13879 = {_0, _13877} + {_0, _13878};
  wire [1:0] _13880 = {_0, _9917} + {_0, _10748};
  wire [3:0] _13881 = {_0, _13879} + {_0, _0, _13880};
  wire _13882 = _12301 < _13881;
  wire _13883 = r1872 ^ _13882;
  wire _13884 = _12298 ? coded_block[1872] : r1872;
  wire _13885 = _12296 ? _13883 : _13884;
  always @ (posedge reset or posedge clock) if (reset) r1872 <= 1'd0; else if (_12300) r1872 <= _13885;
  wire [1:0] _13886 = {_0, _1950} + {_0, _2686};
  wire [1:0] _13887 = {_0, _5726} + {_0, _6525};
  wire [2:0] _13888 = {_0, _13886} + {_0, _13887};
  wire [1:0] _13889 = {_0, _9759} + {_0, _11326};
  wire [3:0] _13890 = {_0, _13888} + {_0, _0, _13889};
  wire _13891 = _12301 < _13890;
  wire _13892 = r1871 ^ _13891;
  wire _13893 = _12298 ? coded_block[1871] : r1871;
  wire _13894 = _12296 ? _13892 : _13893;
  always @ (posedge reset or posedge clock) if (reset) r1871 <= 1'd0; else if (_12300) r1871 <= _13894;
  wire [1:0] _13895 = {_0, _1886} + {_0, _2719};
  wire [1:0] _13896 = {_0, _6045} + {_0, _7132};
  wire [2:0] _13897 = {_0, _13895} + {_0, _13896};
  wire [1:0] _13898 = {_0, _9724} + {_0, _10846};
  wire [3:0] _13899 = {_0, _13897} + {_0, _0, _13898};
  wire _13900 = _12301 < _13899;
  wire _13901 = r1870 ^ _13900;
  wire _13902 = _12298 ? coded_block[1870] : r1870;
  wire _13903 = _12296 ? _13901 : _13902;
  always @ (posedge reset or posedge clock) if (reset) r1870 <= 1'd0; else if (_12300) r1870 <= _13903;
  wire [1:0] _13904 = {_0, _894} + {_0, _2813};
  wire [1:0] _13905 = {_0, _4319} + {_0, _6621};
  wire [2:0] _13906 = {_0, _13904} + {_0, _13905};
  wire [1:0] _13907 = {_0, _9566} + {_0, _11259};
  wire [3:0] _13908 = {_0, _13906} + {_0, _0, _13907};
  wire _13909 = _12301 < _13908;
  wire _13910 = r1869 ^ _13909;
  wire _13911 = _12298 ? coded_block[1869] : r1869;
  wire _13912 = _12296 ? _13910 : _13911;
  always @ (posedge reset or posedge clock) if (reset) r1869 <= 1'd0; else if (_12300) r1869 <= _13912;
  wire [1:0] _13913 = {_0, _1662} + {_0, _3964};
  wire [1:0] _13914 = {_0, _4958} + {_0, _6494};
  wire [2:0] _13915 = {_0, _13913} + {_0, _13914};
  wire [1:0] _13916 = {_0, _9534} + {_0, _10335};
  wire [3:0] _13917 = {_0, _13915} + {_0, _0, _13916};
  wire _13918 = _12301 < _13917;
  wire _13919 = r1868 ^ _13918;
  wire _13920 = _12298 ? coded_block[1868] : r1868;
  wire _13921 = _12296 ? _13919 : _13920;
  always @ (posedge reset or posedge clock) if (reset) r1868 <= 1'd0; else if (_12300) r1868 <= _13921;
  wire [1:0] _13922 = {_0, _383} + {_0, _2623};
  wire [1:0] _13923 = {_0, _4861} + {_0, _7548};
  wire [2:0] _13924 = {_0, _13922} + {_0, _13923};
  wire [1:0] _13925 = {_0, _9342} + {_0, _10590};
  wire [3:0] _13926 = {_0, _13924} + {_0, _0, _13925};
  wire _13927 = _12301 < _13926;
  wire _13928 = r1867 ^ _13927;
  wire _13929 = _12298 ? coded_block[1867] : r1867;
  wire _13930 = _12296 ? _13928 : _13929;
  always @ (posedge reset or posedge clock) if (reset) r1867 <= 1'd0; else if (_12300) r1867 <= _13930;
  wire [1:0] _13931 = {_0, _1662} + {_0, _2557};
  wire [1:0] _13932 = {_0, _5534} + {_0, _7675};
  wire [2:0] _13933 = {_0, _13931} + {_0, _13932};
  wire [1:0] _13934 = {_0, _9181} + {_0, _11485};
  wire [3:0] _13935 = {_0, _13933} + {_0, _0, _13934};
  wire _13936 = _12301 < _13935;
  wire _13937 = r1866 ^ _13936;
  wire _13938 = _12298 ? coded_block[1866] : r1866;
  wire _13939 = _12296 ? _13937 : _13938;
  always @ (posedge reset or posedge clock) if (reset) r1866 <= 1'd0; else if (_12300) r1866 <= _13939;
  wire [1:0] _13940 = {_0, _2044} + {_0, _3933};
  wire [1:0] _13941 = {_0, _5949} + {_0, _6814};
  wire [2:0] _13942 = {_0, _13940} + {_0, _13941};
  wire [1:0] _13943 = {_0, _9149} + {_0, _10590};
  wire [3:0] _13944 = {_0, _13942} + {_0, _0, _13943};
  wire _13945 = _12301 < _13944;
  wire _13946 = r1865 ^ _13945;
  wire _13947 = _12298 ? coded_block[1865] : r1865;
  wire _13948 = _12296 ? _13946 : _13947;
  always @ (posedge reset or posedge clock) if (reset) r1865 <= 1'd0; else if (_12300) r1865 <= _13948;
  wire [1:0] _13949 = {_0, _1662} + {_0, _3773};
  wire [1:0] _13950 = {_0, _4861} + {_0, _7454};
  wire [2:0] _13951 = {_0, _13949} + {_0, _13950};
  wire [1:0] _13952 = {_0, _8574} + {_0, _10941};
  wire [3:0] _13953 = {_0, _13951} + {_0, _0, _13952};
  wire _13954 = _12301 < _13953;
  wire _13955 = r1864 ^ _13954;
  wire _13956 = _12298 ? coded_block[1864] : r1864;
  wire _13957 = _12296 ? _13955 : _13956;
  always @ (posedge reset or posedge clock) if (reset) r1864 <= 1'd0; else if (_12300) r1864 <= _13957;
  wire [1:0] _13958 = {_0, _2013} + {_0, _2719};
  wire [1:0] _13959 = {_0, _5342} + {_0, _7326};
  wire [2:0] _13960 = {_0, _13958} + {_0, _13959};
  wire [1:0] _13961 = {_0, _8480} + {_0, _11196};
  wire [3:0] _13962 = {_0, _13960} + {_0, _0, _13961};
  wire _13963 = _12301 < _13962;
  wire _13964 = r1863 ^ _13963;
  wire _13965 = _12298 ? coded_block[1863] : r1863;
  wire _13966 = _12296 ? _13964 : _13965;
  always @ (posedge reset or posedge clock) if (reset) r1863 <= 1'd0; else if (_12300) r1863 <= _13966;
  wire [1:0] _13967 = {_0, _831} + {_0, _3870};
  wire [1:0] _13968 = {_0, _5342} + {_0, _6687};
  wire [2:0] _13969 = {_0, _13967} + {_0, _13968};
  wire [1:0] _13970 = {_0, _8415} + {_0, _10621};
  wire [3:0] _13971 = {_0, _13969} + {_0, _0, _13970};
  wire _13972 = _12301 < _13971;
  wire _13973 = r1862 ^ _13972;
  wire _13974 = _12298 ? coded_block[1862] : r1862;
  wire _13975 = _12296 ? _13973 : _13974;
  always @ (posedge reset or posedge clock) if (reset) r1862 <= 1'd0; else if (_12300) r1862 <= _13975;
  wire [1:0] _13976 = {_0, _1502} + {_0, _2878};
  wire [1:0] _13977 = {_0, _5183} + {_0, _8123};
  wire [2:0] _13978 = {_0, _13976} + {_0, _13977};
  wire [1:0] _13979 = {_0, _9822} + {_0, _12092};
  wire [3:0] _13980 = {_0, _13978} + {_0, _0, _13979};
  wire _13981 = _12301 < _13980;
  wire _13982 = r1861 ^ _13981;
  wire _13983 = _12298 ? coded_block[1861] : r1861;
  wire _13984 = _12296 ? _13982 : _13983;
  always @ (posedge reset or posedge clock) if (reset) r1861 <= 1'd0; else if (_12300) r1861 <= _13984;
  wire [1:0] _13985 = {_0, _383} + {_0, _2144};
  wire [1:0] _13986 = {_0, _5884} + {_0, _8092};
  wire [2:0] _13987 = {_0, _13985} + {_0, _13986};
  wire [1:0] _13988 = {_0, _9949} + {_0, _10366};
  wire [3:0] _13989 = {_0, _13987} + {_0, _0, _13988};
  wire _13990 = _12301 < _13989;
  wire _13991 = r1860 ^ _13990;
  wire _13992 = _12298 ? coded_block[1860] : r1860;
  wire _13993 = _12296 ? _13991 : _13992;
  always @ (posedge reset or posedge clock) if (reset) r1860 <= 1'd0; else if (_12300) r1860 <= _13993;
  wire [1:0] _13994 = {_0, _289} + {_0, _4028};
  wire [1:0] _13995 = {_0, _4830} + {_0, _8059};
  wire [2:0] _13996 = {_0, _13994} + {_0, _13995};
  wire [1:0] _13997 = {_0, _9630} + {_0, _11806};
  wire [3:0] _13998 = {_0, _13996} + {_0, _0, _13997};
  wire _13999 = _12301 < _13998;
  wire _14000 = r1859 ^ _13999;
  wire _14001 = _12298 ? coded_block[1859] : r1859;
  wire _14002 = _12296 ? _14000 : _14001;
  always @ (posedge reset or posedge clock) if (reset) r1859 <= 1'd0; else if (_12300) r1859 <= _14002;
  wire [1:0] _14003 = {_0, _672} + {_0, _3517};
  wire [1:0] _14004 = {_0, _4830} + {_0, _7931};
  wire [2:0] _14005 = {_0, _14003} + {_0, _14004};
  wire [1:0] _14006 = {_0, _8511} + {_0, _11644};
  wire [3:0] _14007 = {_0, _14005} + {_0, _0, _14006};
  wire _14008 = _12301 < _14007;
  wire _14009 = r1858 ^ _14008;
  wire _14010 = _12298 ? coded_block[1858] : r1858;
  wire _14011 = _12296 ? _14009 : _14010;
  always @ (posedge reset or posedge clock) if (reset) r1858 <= 1'd0; else if (_12300) r1858 <= _14011;
  wire [1:0] _14012 = {_0, _672} + {_0, _2367};
  wire [1:0] _14013 = {_0, _5501} + {_0, _7868};
  wire [2:0] _14014 = {_0, _14012} + {_0, _14013};
  wire [1:0] _14015 = {_0, _8352} + {_0, _11771};
  wire [3:0] _14016 = {_0, _14014} + {_0, _0, _14015};
  wire _14017 = _12301 < _14016;
  wire _14018 = r1857 ^ _14017;
  wire _14019 = _12298 ? coded_block[1857] : r1857;
  wire _14020 = _12296 ? _14018 : _14019;
  always @ (posedge reset or posedge clock) if (reset) r1857 <= 1'd0; else if (_12300) r1857 <= _14020;
  wire [1:0] _14021 = {_0, _1312} + {_0, _3997};
  wire [1:0] _14022 = {_0, _4319} + {_0, _7773};
  wire [2:0] _14023 = {_0, _14021} + {_0, _14022};
  wire [1:0] _14024 = {_0, _9661} + {_0, _10272};
  wire [3:0] _14025 = {_0, _14023} + {_0, _0, _14024};
  wire _14026 = _12301 < _14025;
  wire _14027 = r1856 ^ _14026;
  wire _14028 = _12298 ? coded_block[1856] : r1856;
  wire _14029 = _12296 ? _14027 : _14028;
  always @ (posedge reset or posedge clock) if (reset) r1856 <= 1'd0; else if (_12300) r1856 <= _14029;
  wire [1:0] _14030 = {_0, _2044} + {_0, _2112};
  wire [1:0] _14031 = {_0, _4958} + {_0, _7710};
  wire [2:0] _14032 = {_0, _14030} + {_0, _14031};
  wire [1:0] _14033 = {_0, _9661} + {_0, _12219};
  wire [3:0] _14034 = {_0, _14032} + {_0, _0, _14033};
  wire _14035 = _12301 < _14034;
  wire _14036 = r1855 ^ _14035;
  wire _14037 = _12298 ? coded_block[1855] : r1855;
  wire _14038 = _12296 ? _14036 : _14037;
  always @ (posedge reset or posedge clock) if (reset) r1855 <= 1'd0; else if (_12300) r1855 <= _14038;
  wire [1:0] _14039 = {_0, _672} + {_0, _2144};
  wire [1:0] _14040 = {_0, _4703} + {_0, _7612};
  wire [2:0] _14041 = {_0, _14039} + {_0, _14040};
  wire [1:0] _14042 = {_0, _8926} + {_0, _12027};
  wire [3:0] _14043 = {_0, _14041} + {_0, _0, _14042};
  wire _14044 = _12301 < _14043;
  wire _14045 = r1854 ^ _14044;
  wire _14046 = _12298 ? coded_block[1854] : r1854;
  wire _14047 = _12296 ? _14045 : _14046;
  always @ (posedge reset or posedge clock) if (reset) r1854 <= 1'd0; else if (_12300) r1854 <= _14047;
  wire [1:0] _14048 = {_0, _1950} + {_0, _2813};
  wire [1:0] _14049 = {_0, _5565} + {_0, _7517};
  wire [2:0] _14050 = {_0, _14048} + {_0, _14049};
  wire [1:0] _14051 = {_0, _10077} + {_0, _10973};
  wire [3:0] _14052 = {_0, _14050} + {_0, _0, _14051};
  wire _14053 = _12301 < _14052;
  wire _14054 = r1853 ^ _14053;
  wire _14055 = _12298 ? coded_block[1853] : r1853;
  wire _14056 = _12296 ? _14054 : _14055;
  always @ (posedge reset or posedge clock) if (reset) r1853 <= 1'd0; else if (_12300) r1853 <= _14056;
  wire [1:0] _14057 = {_0, _672} + {_0, _3870};
  wire [1:0] _14058 = {_0, _6045} + {_0, _7420};
  wire [2:0] _14059 = {_0, _14057} + {_0, _14058};
  wire [1:0] _14060 = {_0, _8701} + {_0, _10717};
  wire [3:0] _14061 = {_0, _14059} + {_0, _0, _14060};
  wire _14062 = _12301 < _14061;
  wire _14063 = r1852 ^ _14062;
  wire _14064 = _12298 ? coded_block[1852] : r1852;
  wire _14065 = _12296 ? _14063 : _14064;
  always @ (posedge reset or posedge clock) if (reset) r1852 <= 1'd0; else if (_12300) r1852 <= _14065;
  wire [1:0] _14066 = {_0, _1886} + {_0, _2112};
  wire [1:0] _14067 = {_0, _4350} + {_0, _7036};
  wire [2:0] _14068 = {_0, _14066} + {_0, _14067};
  wire [1:0] _14069 = {_0, _8830} + {_0, _12092};
  wire [3:0] _14070 = {_0, _14068} + {_0, _0, _14069};
  wire _14071 = _12301 < _14070;
  wire _14072 = r1851 ^ _14071;
  wire _14073 = _12298 ? coded_block[1851] : r1851;
  wire _14074 = _12296 ? _14072 : _14073;
  always @ (posedge reset or posedge clock) if (reset) r1851 <= 1'd0; else if (_12300) r1851 <= _14074;
  wire [1:0] _14075 = {_0, _128} + {_0, _3262};
  wire [1:0] _14076 = {_0, _4319} + {_0, _6781};
  wire [2:0] _14077 = {_0, _14075} + {_0, _14076};
  wire [1:0] _14078 = {_0, _9311} + {_0, _10783};
  wire [3:0] _14079 = {_0, _14077} + {_0, _0, _14078};
  wire _14080 = _12301 < _14079;
  wire _14081 = r1850 ^ _14080;
  wire _14082 = _12298 ? coded_block[1850] : r1850;
  wire _14083 = _12296 ? _14081 : _14082;
  always @ (posedge reset or posedge clock) if (reset) r1850 <= 1'd0; else if (_12300) r1850 <= _14083;
  wire [1:0] _14084 = {_0, _639} + {_0, _2175};
  wire [1:0] _14085 = {_0, _5597} + {_0, _6558};
  wire [2:0] _14086 = {_0, _14084} + {_0, _14085};
  wire [1:0] _14087 = {_0, _8701} + {_0, _12219};
  wire [3:0] _14088 = {_0, _14086} + {_0, _0, _14087};
  wire _14089 = _12301 < _14088;
  wire _14090 = r1849 ^ _14089;
  wire _14091 = _12298 ? coded_block[1849] : r1849;
  wire _14092 = _12296 ? _14090 : _14091;
  always @ (posedge reset or posedge clock) if (reset) r1849 <= 1'd0; else if (_12300) r1849 <= _14092;
  wire [1:0] _14093 = {_0, _894} + {_0, _2336};
  wire [1:0] _14094 = {_0, _4542} + {_0, _6397};
  wire [2:0] _14095 = {_0, _14093} + {_0, _14094};
  wire [1:0] _14096 = {_0, _8830} + {_0, _12027};
  wire [3:0] _14097 = {_0, _14095} + {_0, _0, _14096};
  wire _14098 = _12301 < _14097;
  wire _14099 = r1848 ^ _14098;
  wire _14100 = _12298 ? coded_block[1848] : r1848;
  wire _14101 = _12296 ? _14099 : _14100;
  always @ (posedge reset or posedge clock) if (reset) r1848 <= 1'd0; else if (_12300) r1848 <= _14101;
  wire [1:0] _14102 = {_0, _1758} + {_0, _2302};
  wire [1:0] _14103 = {_0, _4830} + {_0, _6303};
  wire [2:0] _14104 = {_0, _14102} + {_0, _14103};
  wire [1:0] _14105 = {_0, _9661} + {_0, _11389};
  wire [3:0] _14106 = {_0, _14104} + {_0, _0, _14105};
  wire _14107 = _12301 < _14106;
  wire _14108 = r1847 ^ _14107;
  wire _14109 = _12298 ? coded_block[1847] : r1847;
  wire _14110 = _12296 ? _14108 : _14109;
  always @ (posedge reset or posedge clock) if (reset) r1847 <= 1'd0; else if (_12300) r1847 <= _14110;
  wire [1:0] _14111 = {_0, _1950} + {_0, _2910};
  wire [1:0] _14112 = {_0, _4350} + {_0, _6239};
  wire [2:0] _14113 = {_0, _14111} + {_0, _14112};
  wire [1:0] _14114 = {_0, _8225} + {_0, _10366};
  wire [3:0] _14115 = {_0, _14113} + {_0, _0, _14114};
  wire _14116 = _12301 < _14115;
  wire _14117 = r1846 ^ _14116;
  wire _14118 = _12298 ? coded_block[1846] : r1846;
  wire _14119 = _12296 ? _14117 : _14118;
  always @ (posedge reset or posedge clock) if (reset) r1846 <= 1'd0; else if (_12300) r1846 <= _14119;
  wire [1:0] _14120 = {_0, _128} + {_0, _2494};
  wire [1:0] _14121 = {_0, _4384} + {_0, _6176};
  wire [2:0] _14122 = {_0, _14120} + {_0, _14121};
  wire [1:0] _14123 = {_0, _8511} + {_0, _10748};
  wire [3:0] _14124 = {_0, _14122} + {_0, _0, _14123};
  wire _14125 = _12301 < _14124;
  wire _14126 = r1845 ^ _14125;
  wire _14127 = _12298 ? coded_block[1845] : r1845;
  wire _14128 = _12296 ? _14126 : _14127;
  always @ (posedge reset or posedge clock) if (reset) r1845 <= 1'd0; else if (_12300) r1845 <= _14128;
  wire [1:0] _14129 = {_0, _672} + {_0, _3294};
  wire [1:0] _14130 = {_0, _6076} + {_0, _6718};
  wire [2:0] _14131 = {_0, _14129} + {_0, _14130};
  wire [1:0] _14132 = {_0, _8319} + {_0, _11996};
  wire [3:0] _14133 = {_0, _14131} + {_0, _0, _14132};
  wire _14134 = _12301 < _14133;
  wire _14135 = r1844 ^ _14134;
  wire _14136 = _12298 ? coded_block[1844] : r1844;
  wire _14137 = _12296 ? _14135 : _14136;
  always @ (posedge reset or posedge clock) if (reset) r1844 <= 1'd0; else if (_12300) r1844 <= _14137;
  wire [1:0] _14138 = {_0, _383} + {_0, _3997};
  wire [1:0] _14139 = {_0, _5853} + {_0, _6270};
  wire [2:0] _14140 = {_0, _14138} + {_0, _14139};
  wire [1:0] _14141 = {_0, _9469} + {_0, _11295};
  wire [3:0] _14142 = {_0, _14140} + {_0, _0, _14141};
  wire _14143 = _12301 < _14142;
  wire _14144 = r1843 ^ _14143;
  wire _14145 = _12298 ? coded_block[1843] : r1843;
  wire _14146 = _12296 ? _14144 : _14145;
  always @ (posedge reset or posedge clock) if (reset) r1843 <= 1'd0; else if (_12300) r1843 <= _14146;
  wire [1:0] _14147 = {_0, _510} + {_0, _2813};
  wire [1:0] _14148 = {_0, _5821} + {_0, _7357};
  wire [2:0] _14149 = {_0, _14147} + {_0, _14148};
  wire [1:0] _14150 = {_0, _8383} + {_0, _11196};
  wire [3:0] _14151 = {_0, _14149} + {_0, _0, _14150};
  wire _14152 = _12301 < _14151;
  wire _14153 = r1842 ^ _14152;
  wire _14154 = _12298 ? coded_block[1842] : r1842;
  wire _14155 = _12296 ? _14153 : _14154;
  always @ (posedge reset or posedge clock) if (reset) r1842 <= 1'd0; else if (_12300) r1842 <= _14155;
  wire [1:0] _14156 = {_0, _831} + {_0, _2910};
  wire [1:0] _14157 = {_0, _5757} + {_0, _6494};
  wire [2:0] _14158 = {_0, _14156} + {_0, _14157};
  wire [1:0] _14159 = {_0, _8446} + {_0, _11004};
  wire [3:0] _14160 = {_0, _14158} + {_0, _0, _14159};
  wire _14161 = _12301 < _14160;
  wire _14162 = r1841 ^ _14161;
  wire _14163 = _12298 ? coded_block[1841] : r1841;
  wire _14164 = _12296 ? _14162 : _14163;
  always @ (posedge reset or posedge clock) if (reset) r1841 <= 1'd0; else if (_12300) r1841 <= _14164;
  wire [1:0] _14165 = {_0, _1758} + {_0, _3262};
  wire [1:0] _14166 = {_0, _4926} + {_0, _7996};
  wire [2:0] _14167 = {_0, _14165} + {_0, _14166};
  wire [1:0] _14168 = {_0, _8446} + {_0, _10973};
  wire [3:0] _14169 = {_0, _14167} + {_0, _0, _14168};
  wire _14170 = _12301 < _14169;
  wire _14171 = r1840 ^ _14170;
  wire _14172 = _12298 ? coded_block[1840] : r1840;
  wire _14173 = _12296 ? _14171 : _14172;
  always @ (posedge reset or posedge clock) if (reset) r1840 <= 1'd0; else if (_12300) r1840 <= _14173;
  wire [1:0] _14174 = {_0, _894} + {_0, _2239};
  wire [1:0] _14175 = {_0, _4895} + {_0, _6494};
  wire [2:0] _14176 = {_0, _14174} + {_0, _14175};
  wire [1:0] _14177 = {_0, _10172} + {_0, _11228};
  wire [3:0] _14178 = {_0, _14176} + {_0, _0, _14177};
  wire _14179 = _12301 < _14178;
  wire _14180 = r1839 ^ _14179;
  wire _14181 = _12298 ? coded_block[1839] : r1839;
  wire _14182 = _12296 ? _14180 : _14181;
  always @ (posedge reset or posedge clock) if (reset) r1839 <= 1'd0; else if (_12300) r1839 <= _14182;
  wire [1:0] _14183 = {_0, _1886} + {_0, _3964};
  wire [1:0] _14184 = {_0, _4798} + {_0, _7548};
  wire [2:0] _14185 = {_0, _14183} + {_0, _14184};
  wire [1:0] _14186 = {_0, _9503} + {_0, _12061};
  wire [3:0] _14187 = {_0, _14185} + {_0, _0, _14186};
  wire _14188 = _12301 < _14187;
  wire _14189 = r1838 ^ _14188;
  wire _14190 = _12298 ? coded_block[1838] : r1838;
  wire _14191 = _12296 ? _14189 : _14190;
  always @ (posedge reset or posedge clock) if (reset) r1838 <= 1'd0; else if (_12300) r1838 <= _14191;
  wire [1:0] _14192 = {_0, _97} + {_0, _2367};
  wire [1:0] _14193 = {_0, _4767} + {_0, _7548};
  wire [2:0] _14194 = {_0, _14192} + {_0, _14193};
  wire [1:0] _14195 = {_0, _10204} + {_0, _11806};
  wire [3:0] _14196 = {_0, _14194} + {_0, _0, _14195};
  wire _14197 = _12301 < _14196;
  wire _14198 = r1837 ^ _14197;
  wire _14199 = _12298 ? coded_block[1837] : r1837;
  wire _14200 = _12296 ? _14198 : _14199;
  always @ (posedge reset or posedge clock) if (reset) r1837 <= 1'd0; else if (_12300) r1837 <= _14200;
  wire [1:0] _14201 = {_0, _1726} + {_0, _2399};
  wire [1:0] _14202 = {_0, _4734} + {_0, _8186};
  wire [2:0] _14203 = {_0, _14201} + {_0, _14202};
  wire [1:0] _14204 = {_0, _10077} + {_0, _10272};
  wire [3:0] _14205 = {_0, _14203} + {_0, _0, _14204};
  wire _14206 = _12301 < _14205;
  wire _14207 = r1836 ^ _14206;
  wire _14208 = _12298 ? coded_block[1836] : r1836;
  wire _14209 = _12296 ? _14207 : _14208;
  always @ (posedge reset or posedge clock) if (reset) r1836 <= 1'd0; else if (_12300) r1836 <= _14209;
  wire [1:0] _14210 = {_0, _1662} + {_0, _3453};
  wire [1:0] _14211 = {_0, _4640} + {_0, _6462};
  wire [2:0] _14212 = {_0, _14210} + {_0, _14211};
  wire [1:0] _14213 = {_0, _9085} + {_0, _11069};
  wire [3:0] _14214 = {_0, _14212} + {_0, _0, _14213};
  wire _14215 = _12301 < _14214;
  wire _14216 = r1835 ^ _14215;
  wire _14217 = _12298 ? coded_block[1835] : r1835;
  wire _14218 = _12296 ? _14216 : _14217;
  always @ (posedge reset or posedge clock) if (reset) r1835 <= 1'd0; else if (_12300) r1835 <= _14218;
  wire [1:0] _14219 = {_0, _1662} + {_0, _2910};
  wire [1:0] _14220 = {_0, _4447} + {_0, _7485};
  wire [2:0] _14221 = {_0, _14219} + {_0, _14220};
  wire [1:0] _14222 = {_0, _8288} + {_0, _11516};
  wire [3:0] _14223 = {_0, _14221} + {_0, _0, _14222};
  wire _14224 = _12301 < _14223;
  wire _14225 = r1834 ^ _14224;
  wire _14226 = _12298 ? coded_block[1834] : r1834;
  wire _14227 = _12296 ? _14225 : _14226;
  always @ (posedge reset or posedge clock) if (reset) r1834 <= 1'd0; else if (_12300) r1834 <= _14227;
  wire [1:0] _14228 = {_0, _128} + {_0, _2175};
  wire [1:0] _14229 = {_0, _4223} + {_0, _6270};
  wire [2:0] _14230 = {_0, _14228} + {_0, _14229};
  wire [1:0] _14231 = {_0, _8319} + {_0, _10366};
  wire [3:0] _14232 = {_0, _14230} + {_0, _0, _14231};
  wire _14233 = _12301 < _14232;
  wire _14234 = r1833 ^ _14233;
  wire _14235 = _12298 ? coded_block[1833] : r1833;
  wire _14236 = _12296 ? _14234 : _14235;
  always @ (posedge reset or posedge clock) if (reset) r1833 <= 1'd0; else if (_12300) r1833 <= _14236;
  wire [1:0] _14237 = {_0, _1502} + {_0, _2813};
  wire [1:0] _14238 = {_0, _4192} + {_0, _7485};
  wire [2:0] _14239 = {_0, _14237} + {_0, _14238};
  wire [1:0] _14240 = {_0, _9503} + {_0, _10366};
  wire [3:0] _14241 = {_0, _14239} + {_0, _0, _14240};
  wire _14242 = _12301 < _14241;
  wire _14243 = r1832 ^ _14242;
  wire _14244 = _12298 ? coded_block[1832] : r1832;
  wire _14245 = _12296 ? _14243 : _14244;
  always @ (posedge reset or posedge clock) if (reset) r1832 <= 1'd0; else if (_12300) r1832 <= _14245;
  wire [1:0] _14246 = {_0, _1057} + {_0, _3262};
  wire [1:0] _14247 = {_0, _4129} + {_0, _7389};
  wire [2:0] _14248 = {_0, _14246} + {_0, _14247};
  wire [1:0] _14249 = {_0, _9630} + {_0, _10303};
  wire [3:0] _14250 = {_0, _14248} + {_0, _0, _14249};
  wire _14251 = _12301 < _14250;
  wire _14252 = r1831 ^ _14251;
  wire _14253 = _12298 ? coded_block[1831] : r1831;
  wire _14254 = _12296 ? _14252 : _14253;
  always @ (posedge reset or posedge clock) if (reset) r1831 <= 1'd0; else if (_12300) r1831 <= _14254;
  wire [1:0] _14255 = {_0, _352} + {_0, _4060};
  wire [1:0] _14256 = {_0, _5183} + {_0, _7548};
  wire [2:0] _14257 = {_0, _14255} + {_0, _14256};
  wire [1:0] _14258 = {_0, _10045} + {_0, _11453};
  wire [3:0] _14259 = {_0, _14257} + {_0, _0, _14258};
  wire _14260 = _12301 < _14259;
  wire _14261 = r1830 ^ _14260;
  wire _14262 = _12298 ? coded_block[1830] : r1830;
  wire _14263 = _12296 ? _14261 : _14262;
  always @ (posedge reset or posedge clock) if (reset) r1830 <= 1'd0; else if (_12300) r1830 <= _14263;
  wire [1:0] _14264 = {_0, _383} + {_0, _3901};
  wire [1:0] _14265 = {_0, _5565} + {_0, _6621};
  wire [2:0] _14266 = {_0, _14264} + {_0, _14265};
  wire [1:0] _14267 = {_0, _9085} + {_0, _11613};
  wire [3:0] _14268 = {_0, _14266} + {_0, _0, _14267};
  wire _14269 = _12301 < _14268;
  wire _14270 = r1829 ^ _14269;
  wire _14271 = _12298 ? coded_block[1829] : r1829;
  wire _14272 = _12296 ? _14270 : _14271;
  always @ (posedge reset or posedge clock) if (reset) r1829 <= 1'd0; else if (_12300) r1829 <= _14272;
  wire [1:0] _14273 = {_0, _894} + {_0, _3678};
  wire [1:0] _14274 = {_0, _6045} + {_0, _6525};
  wire [2:0] _14275 = {_0, _14273} + {_0, _14274};
  wire [1:0] _14276 = {_0, _9949} + {_0, _10910};
  wire [3:0] _14277 = {_0, _14275} + {_0, _0, _14276};
  wire _14278 = _12301 < _14277;
  wire _14279 = r1828 ^ _14278;
  wire _14280 = _12298 ? coded_block[1828] : r1828;
  wire _14281 = _12296 ? _14279 : _14280;
  always @ (posedge reset or posedge clock) if (reset) r1828 <= 1'd0; else if (_12300) r1828 <= _14281;
  wire [1:0] _14282 = {_0, _2013} + {_0, _3646};
  wire [1:0] _14283 = {_0, _4574} + {_0, _6270};
  wire [2:0] _14284 = {_0, _14282} + {_0, _14283};
  wire [1:0] _14285 = {_0, _8543} + {_0, _10462};
  wire [3:0] _14286 = {_0, _14284} + {_0, _0, _14285};
  wire _14287 = _12301 < _14286;
  wire _14288 = r1827 ^ _14287;
  wire _14289 = _12298 ? coded_block[1827] : r1827;
  wire _14290 = _12296 ? _14288 : _14289;
  always @ (posedge reset or posedge clock) if (reset) r1827 <= 1'd0; else if (_12300) r1827 <= _14290;
  wire [1:0] _14291 = {_0, _1057} + {_0, _3580};
  wire [1:0] _14292 = {_0, _5279} + {_0, _7548};
  wire [2:0] _14293 = {_0, _14291} + {_0, _14292};
  wire [1:0] _14294 = {_0, _9469} + {_0, _11869};
  wire [3:0] _14295 = {_0, _14293} + {_0, _0, _14294};
  wire _14296 = _12301 < _14295;
  wire _14297 = r1826 ^ _14296;
  wire _14298 = _12298 ? coded_block[1826] : r1826;
  wire _14299 = _12296 ? _14297 : _14298;
  always @ (posedge reset or posedge clock) if (reset) r1826 <= 1'd0; else if (_12300) r1826 <= _14299;
  wire [1:0] _14300 = {_0, _1502} + {_0, _3231};
  wire [1:0] _14301 = {_0, _6045} + {_0, _7262};
  wire [2:0] _14302 = {_0, _14300} + {_0, _14301};
  wire [1:0] _14303 = {_0, _8830} + {_0, _11004};
  wire [3:0] _14304 = {_0, _14302} + {_0, _0, _14303};
  wire _14305 = _12301 < _14304;
  wire _14306 = r1825 ^ _14305;
  wire _14307 = _12298 ? coded_block[1825] : r1825;
  wire _14308 = _12296 ? _14306 : _14307;
  always @ (posedge reset or posedge clock) if (reset) r1825 <= 1'd0; else if (_12300) r1825 <= _14308;
  wire [1:0] _14309 = {_0, _128} + {_0, _2655};
  wire [1:0] _14310 = {_0, _4350} + {_0, _6621};
  wire [2:0] _14311 = {_0, _14309} + {_0, _14310};
  wire [1:0] _14312 = {_0, _8543} + {_0, _10941};
  wire [3:0] _14313 = {_0, _14311} + {_0, _0, _14312};
  wire _14314 = _12301 < _14313;
  wire _14315 = r1824 ^ _14314;
  wire _14316 = _12298 ? coded_block[1824] : r1824;
  wire _14317 = _12296 ? _14315 : _14316;
  always @ (posedge reset or posedge clock) if (reset) r1824 <= 1'd0; else if (_12300) r1824 <= _14317;
  wire [1:0] _14318 = {_0, _1568} + {_0, _2430};
  wire [1:0] _14319 = {_0, _5183} + {_0, _7132};
  wire [2:0] _14320 = {_0, _14318} + {_0, _14319};
  wire [1:0] _14321 = {_0, _9693} + {_0, _10590};
  wire [3:0] _14322 = {_0, _14320} + {_0, _0, _14321};
  wire _14323 = _12301 < _14322;
  wire _14324 = r1823 ^ _14323;
  wire _14325 = _12298 ? coded_block[1823] : r1823;
  wire _14326 = _12296 ? _14324 : _14325;
  always @ (posedge reset or posedge clock) if (reset) r1823 <= 1'd0; else if (_12300) r1823 <= _14326;
  wire [1:0] _14327 = {_0, _1120} + {_0, _2271};
  wire [1:0] _14328 = {_0, _4861} + {_0, _7996};
  wire [2:0] _14329 = {_0, _14327} + {_0, _14328};
  wire [1:0] _14330 = {_0, _8352} + {_0, _10846};
  wire [3:0] _14331 = {_0, _14329} + {_0, _0, _14330};
  wire _14332 = _12301 < _14331;
  wire _14333 = r1822 ^ _14332;
  wire _14334 = _12298 ? coded_block[1822] : r1822;
  wire _14335 = _12296 ? _14333 : _14334;
  always @ (posedge reset or posedge clock) if (reset) r1822 <= 1'd0; else if (_12300) r1822 <= _14335;
  wire [1:0] _14336 = {_0, _1981} + {_0, _3997};
  wire [1:0] _14337 = {_0, _6108} + {_0, _6942};
  wire [2:0] _14338 = {_0, _14336} + {_0, _14337};
  wire [1:0] _14339 = {_0, _9693} + {_0, _11644};
  wire [3:0] _14340 = {_0, _14338} + {_0, _0, _14339};
  wire _14341 = _12301 < _14340;
  wire _14342 = r1821 ^ _14341;
  wire _14343 = _12298 ? coded_block[1821] : r1821;
  wire _14344 = _12296 ? _14342 : _14343;
  always @ (posedge reset or posedge clock) if (reset) r1821 <= 1'd0; else if (_12300) r1821 <= _14344;
  wire [1:0] _14345 = {_0, _1854} + {_0, _2336};
  wire [1:0] _14346 = {_0, _5565} + {_0, _7132};
  wire [2:0] _14347 = {_0, _14345} + {_0, _14346};
  wire [1:0] _14348 = {_0, _9311} + {_0, _10685};
  wire [3:0] _14349 = {_0, _14347} + {_0, _0, _14348};
  wire _14350 = _12301 < _14349;
  wire _14351 = r1820 ^ _14350;
  wire _14352 = _12298 ? coded_block[1820] : r1820;
  wire _14353 = _12296 ? _14351 : _14352;
  always @ (posedge reset or posedge clock) if (reset) r1820 <= 1'd0; else if (_12300) r1820 <= _14353;
  wire [1:0] _14354 = {_0, _1823} + {_0, _2686};
  wire [1:0] _14355 = {_0, _5438} + {_0, _7389};
  wire [2:0] _14356 = {_0, _14354} + {_0, _14355};
  wire [1:0] _14357 = {_0, _9949} + {_0, _10846};
  wire [3:0] _14358 = {_0, _14356} + {_0, _0, _14357};
  wire _14359 = _12301 < _14358;
  wire _14360 = r1819 ^ _14359;
  wire _14361 = _12298 ? coded_block[1819] : r1819;
  wire _14362 = _12296 ? _14360 : _14361;
  always @ (posedge reset or posedge clock) if (reset) r1819 <= 1'd0; else if (_12300) r1819 <= _14362;
  wire [1:0] _14363 = {_0, _1631} + {_0, _3167};
  wire [1:0] _14364 = {_0, _4574} + {_0, _7548};
  wire [2:0] _14365 = {_0, _14363} + {_0, _14364};
  wire [1:0] _14366 = {_0, _9693} + {_0, _11196};
  wire [3:0] _14367 = {_0, _14365} + {_0, _0, _14366};
  wire _14368 = _12301 < _14367;
  wire _14369 = r1818 ^ _14368;
  wire _14370 = _12298 ? coded_block[1818] : r1818;
  wire _14371 = _12296 ? _14369 : _14370;
  always @ (posedge reset or posedge clock) if (reset) r1818 <= 1'd0; else if (_12300) r1818 <= _14371;
  wire [1:0] _14372 = {_0, _1470} + {_0, _3453};
  wire [1:0] _14373 = {_0, _4350} + {_0, _7675};
  wire [2:0] _14374 = {_0, _14372} + {_0, _14373};
  wire [1:0] _14375 = {_0, _8767} + {_0, _11358};
  wire [3:0] _14376 = {_0, _14374} + {_0, _0, _14375};
  wire _14377 = _12301 < _14376;
  wire _14378 = r1817 ^ _14377;
  wire _14379 = _12298 ? coded_block[1817] : r1817;
  wire _14380 = _12296 ? _14378 : _14379;
  always @ (posedge reset or posedge clock) if (reset) r1817 <= 1'd0; else if (_12300) r1817 <= _14380;
  wire [1:0] _14381 = {_0, _1343} + {_0, _4028};
  wire [1:0] _14382 = {_0, _4350} + {_0, _7804};
  wire [2:0] _14383 = {_0, _14381} + {_0, _14382};
  wire [1:0] _14384 = {_0, _9693} + {_0, _10272};
  wire [3:0] _14385 = {_0, _14383} + {_0, _0, _14384};
  wire _14386 = _12301 < _14385;
  wire _14387 = r1816 ^ _14386;
  wire _14388 = _12298 ? coded_block[1816] : r1816;
  wire _14389 = _12296 ? _14387 : _14388;
  always @ (posedge reset or posedge clock) if (reset) r1816 <= 1'd0; else if (_12300) r1816 <= _14389;
  wire [1:0] _14390 = {_0, _990} + {_0, _2750};
  wire [1:0] _14391 = {_0, _4478} + {_0, _6687};
  wire [2:0] _14392 = {_0, _14390} + {_0, _14391};
  wire [1:0] _14393 = {_0, _8543} + {_0, _10973};
  wire [3:0] _14394 = {_0, _14392} + {_0, _0, _14393};
  wire _14395 = _12301 < _14394;
  wire _14396 = r1815 ^ _14395;
  wire _14397 = _12298 ? coded_block[1815] : r1815;
  wire _14398 = _12296 ? _14396 : _14397;
  always @ (posedge reset or posedge clock) if (reset) r1815 <= 1'd0; else if (_12300) r1815 <= _14398;
  wire [1:0] _14399 = {_0, _800} + {_0, _3964};
  wire [1:0] _14400 = {_0, _4542} + {_0, _7675};
  wire [2:0] _14401 = {_0, _14399} + {_0, _14400};
  wire [1:0] _14402 = {_0, _10045} + {_0, _10527};
  wire [3:0] _14403 = {_0, _14401} + {_0, _0, _14402};
  wire _14404 = _12301 < _14403;
  wire _14405 = r1814 ^ _14404;
  wire _14406 = _12298 ? coded_block[1814] : r1814;
  wire _14407 = _12296 ? _14405 : _14406;
  always @ (posedge reset or posedge clock) if (reset) r1814 <= 1'd0; else if (_12300) r1814 <= _14407;
  wire [1:0] _14408 = {_0, _766} + {_0, _2302};
  wire [1:0] _14409 = {_0, _5726} + {_0, _6687};
  wire [2:0] _14410 = {_0, _14408} + {_0, _14409};
  wire [1:0] _14411 = {_0, _8830} + {_0, _10335};
  wire [3:0] _14412 = {_0, _14410} + {_0, _0, _14411};
  wire _14413 = _12301 < _14412;
  wire _14414 = r1813 ^ _14413;
  wire _14415 = _12298 ? coded_block[1813] : r1813;
  wire _14416 = _12296 ? _14414 : _14415;
  always @ (posedge reset or posedge clock) if (reset) r1813 <= 1'd0; else if (_12300) r1813 <= _14416;
  wire [1:0] _14417 = {_0, _576} + {_0, _2175};
  wire [1:0] _14418 = {_0, _6045} + {_0, _6462};
  wire [2:0] _14419 = {_0, _14417} + {_0, _14418};
  wire [1:0] _14420 = {_0, _9661} + {_0, _11485};
  wire [3:0] _14421 = {_0, _14419} + {_0, _0, _14420};
  wire _14422 = _12301 < _14421;
  wire _14423 = r1812 ^ _14422;
  wire _14424 = _12298 ? coded_block[1812] : r1812;
  wire _14425 = _12296 ? _14423 : _14424;
  always @ (posedge reset or posedge clock) if (reset) r1812 <= 1'd0; else if (_12300) r1812 <= _14425;
  wire [1:0] _14426 = {_0, _479} + {_0, _2175};
  wire [1:0] _14427 = {_0, _5310} + {_0, _7675};
  wire [2:0] _14428 = {_0, _14426} + {_0, _14427};
  wire [1:0] _14429 = {_0, _10172} + {_0, _11581};
  wire [3:0] _14430 = {_0, _14428} + {_0, _0, _14429};
  wire _14431 = _12301 < _14430;
  wire _14432 = r1811 ^ _14431;
  wire _14433 = _12298 ? coded_block[1811] : r1811;
  wire _14434 = _12296 ? _14432 : _14433;
  always @ (posedge reset or posedge clock) if (reset) r1811 <= 1'd0; else if (_12300) r1811 <= _14434;
  wire [1:0] _14435 = {_0, _447} + {_0, _2494};
  wire [1:0] _14436 = {_0, _4542} + {_0, _6589};
  wire [2:0] _14437 = {_0, _14435} + {_0, _14436};
  wire [1:0] _14438 = {_0, _8638} + {_0, _10685};
  wire [3:0] _14439 = {_0, _14437} + {_0, _0, _14438};
  wire _14440 = _12301 < _14439;
  wire _14441 = r1810 ^ _14440;
  wire _14442 = _12298 ? coded_block[1810] : r1810;
  wire _14443 = _12296 ? _14441 : _14442;
  always @ (posedge reset or posedge clock) if (reset) r1810 <= 1'd0; else if (_12300) r1810 <= _14443;
  wire [1:0] _14444 = {_0, _510} + {_0, _3678};
  wire [1:0] _14445 = {_0, _4256} + {_0, _7389};
  wire [2:0] _14446 = {_0, _14444} + {_0, _14445};
  wire [1:0] _14447 = {_0, _9759} + {_0, _12251};
  wire [3:0] _14448 = {_0, _14446} + {_0, _0, _14447};
  wire _14449 = _12301 < _14448;
  wire _14450 = r1809 ^ _14449;
  wire _14451 = _12298 ? coded_block[1809] : r1809;
  wire _14452 = _12296 ? _14450 : _14451;
  always @ (posedge reset or posedge clock) if (reset) r1809 <= 1'd0; else if (_12300) r1809 <= _14452;
  wire [1:0] _14453 = {_0, _97} + {_0, _3773};
  wire [1:0] _14454 = {_0, _5342} + {_0, _7517};
  wire [2:0] _14455 = {_0, _14453} + {_0, _14454};
  wire [1:0] _14456 = {_0, _8894} + {_0, _12188};
  wire [3:0] _14457 = {_0, _14455} + {_0, _0, _14456};
  wire _14458 = _12301 < _14457;
  wire _14459 = r1808 ^ _14458;
  wire _14460 = _12298 ? coded_block[1808] : r1808;
  wire _14461 = _12296 ? _14459 : _14460;
  always @ (posedge reset or posedge clock) if (reset) r1808 <= 1'd0; else if (_12300) r1808 <= _14461;
  wire [1:0] _14462 = {_0, _576} + {_0, _3422};
  wire [1:0] _14463 = {_0, _4734} + {_0, _7837};
  wire [2:0] _14464 = {_0, _14462} + {_0, _14463};
  wire [1:0] _14465 = {_0, _8415} + {_0, _11550};
  wire [3:0] _14466 = {_0, _14464} + {_0, _0, _14465};
  wire _14467 = _12301 < _14466;
  wire _14468 = r1807 ^ _14467;
  wire _14469 = _12298 ? coded_block[1807] : r1807;
  wire _14470 = _12296 ? _14468 : _14469;
  always @ (posedge reset or posedge clock) if (reset) r1807 <= 1'd0; else if (_12300) r1807 <= _14470;
  wire [1:0] _14471 = {_0, _990} + {_0, _3390};
  wire [1:0] _14472 = {_0, _5310} + {_0, _7710};
  wire [2:0] _14473 = {_0, _14471} + {_0, _14472};
  wire [1:0] _14474 = {_0, _8480} + {_0, _11132};
  wire [3:0] _14475 = {_0, _14473} + {_0, _0, _14474};
  wire _14476 = _12301 < _14475;
  wire _14477 = r1806 ^ _14476;
  wire _14478 = _12298 ? coded_block[1806] : r1806;
  wire _14479 = _12296 ? _14477 : _14478;
  always @ (posedge reset or posedge clock) if (reset) r1806 <= 1'd0; else if (_12300) r1806 <= _14479;
  wire [1:0] _14480 = {_0, _1981} + {_0, _3037};
  wire [1:0] _14481 = {_0, _4830} + {_0, _8092};
  wire [2:0] _14482 = {_0, _14480} + {_0, _14481};
  wire [1:0] _14483 = {_0, _10204} + {_0, _11038};
  wire [3:0] _14484 = {_0, _14482} + {_0, _0, _14483};
  wire _14485 = _12301 < _14484;
  wire _14486 = r1805 ^ _14485;
  wire _14487 = _12298 ? coded_block[1805] : r1805;
  wire _14488 = _12296 ? _14486 : _14487;
  always @ (posedge reset or posedge clock) if (reset) r1805 <= 1'd0; else if (_12300) r1805 <= _14488;
  wire [1:0] _14489 = {_0, _1854} + {_0, _2719};
  wire [1:0] _14490 = {_0, _5470} + {_0, _7420};
  wire [2:0] _14491 = {_0, _14489} + {_0, _14490};
  wire [1:0] _14492 = {_0, _9980} + {_0, _10877};
  wire [3:0] _14493 = {_0, _14491} + {_0, _0, _14492};
  wire _14494 = _12301 < _14493;
  wire _14495 = r1804 ^ _14494;
  wire _14496 = _12298 ? coded_block[1804] : r1804;
  wire _14497 = _12296 ? _14495 : _14496;
  always @ (posedge reset or posedge clock) if (reset) r1804 <= 1'd0; else if (_12300) r1804 <= _14497;
  wire [1:0] _14498 = {_0, _958} + {_0, _3422};
  wire [1:0] _14499 = {_0, _4767} + {_0, _6494};
  wire [2:0] _14500 = {_0, _14498} + {_0, _14499};
  wire [1:0] _14501 = {_0, _8701} + {_0, _10558};
  wire [3:0] _14502 = {_0, _14500} + {_0, _0, _14501};
  wire _14503 = _12301 < _14502;
  wire _14504 = r1803 ^ _14503;
  wire _14505 = _12298 ? coded_block[1803] : r1803;
  wire _14506 = _12296 ? _14504 : _14505;
  always @ (posedge reset or posedge clock) if (reset) r1803 <= 1'd0; else if (_12300) r1803 <= _14506;
  wire [1:0] _14507 = {_0, _766} + {_0, _2782};
  wire [1:0] _14508 = {_0, _4895} + {_0, _7741};
  wire [2:0] _14509 = {_0, _14507} + {_0, _14508};
  wire [1:0] _14510 = {_0, _8480} + {_0, _10430};
  wire [3:0] _14511 = {_0, _14509} + {_0, _0, _14510};
  wire _14512 = _12301 < _14511;
  wire _14513 = r1802 ^ _14512;
  wire _14514 = _12298 ? coded_block[1802] : r1802;
  wire _14515 = _12296 ? _14513 : _14514;
  always @ (posedge reset or posedge clock) if (reset) r1802 <= 1'd0; else if (_12300) r1802 <= _14515;
  wire [1:0] _14516 = {_0, _128} + {_0, _2557};
  wire [1:0] _14517 = {_0, _5246} + {_0, _7036};
  wire [2:0] _14518 = {_0, _14516} + {_0, _14517};
  wire [1:0] _14519 = {_0, _8288} + {_0, _10399};
  wire [3:0] _14520 = {_0, _14518} + {_0, _0, _14519};
  wire _14521 = _12301 < _14520;
  wire _14522 = r1801 ^ _14521;
  wire _14523 = _12298 ? coded_block[1801] : r1801;
  wire _14524 = _12296 ? _14522 : _14523;
  always @ (posedge reset or posedge clock) if (reset) r1801 <= 1'd0; else if (_12300) r1801 <= _14524;
  wire [1:0] _14525 = {_0, _831} + {_0, _3836};
  wire [1:0] _14526 = {_0, _5470} + {_0, _7230};
  wire [2:0] _14527 = {_0, _14525} + {_0, _14526};
  wire [1:0] _14528 = {_0, _10235} + {_0, _11771};
  wire [3:0] _14529 = {_0, _14527} + {_0, _0, _14528};
  wire _14530 = _12301 < _14529;
  wire _14531 = r1800 ^ _14530;
  wire _14532 = _12298 ? coded_block[1800] : r1800;
  wire _14533 = _12296 ? _14531 : _14532;
  always @ (posedge reset or posedge clock) if (reset) r1800 <= 1'd0; else if (_12300) r1800 <= _14533;
  wire [1:0] _14534 = {_0, _1981} + {_0, _2847};
  wire [1:0] _14535 = {_0, _5597} + {_0, _7548};
  wire [2:0] _14536 = {_0, _14534} + {_0, _14535};
  wire [1:0] _14537 = {_0, _10108} + {_0, _11004};
  wire [3:0] _14538 = {_0, _14536} + {_0, _0, _14537};
  wire _14539 = _12301 < _14538;
  wire _14540 = r1799 ^ _14539;
  wire _14541 = _12298 ? coded_block[1799] : r1799;
  wire _14542 = _12296 ? _14540 : _14541;
  always @ (posedge reset or posedge clock) if (reset) r1799 <= 1'd0; else if (_12300) r1799 <= _14542;
  wire [1:0] _14543 = {_0, _1854} + {_0, _3294};
  wire [1:0] _14544 = {_0, _5501} + {_0, _7357};
  wire [2:0] _14545 = {_0, _14543} + {_0, _14544};
  wire [1:0] _14546 = {_0, _9790} + {_0, _10973};
  wire [3:0] _14547 = {_0, _14545} + {_0, _0, _14546};
  wire _14548 = _12301 < _14547;
  wire _14549 = r1798 ^ _14548;
  wire _14550 = _12298 ? coded_block[1798] : r1798;
  wire _14551 = _12296 ? _14549 : _14550;
  always @ (posedge reset or posedge clock) if (reset) r1798 <= 1'd0; else if (_12300) r1798 <= _14551;
  wire [1:0] _14552 = {_0, _1758} + {_0, _3453};
  wire [1:0] _14553 = {_0, _4574} + {_0, _6942};
  wire [2:0] _14554 = {_0, _14552} + {_0, _14553};
  wire [1:0] _14555 = {_0, _9438} + {_0, _10846};
  wire [3:0] _14556 = {_0, _14554} + {_0, _0, _14555};
  wire _14557 = _12301 < _14556;
  wire _14558 = r1797 ^ _14557;
  wire _14559 = _12298 ? coded_block[1797] : r1797;
  wire _14560 = _12296 ? _14558 : _14559;
  always @ (posedge reset or posedge clock) if (reset) r1797 <= 1'd0; else if (_12300) r1797 <= _14560;
  wire [1:0] _14561 = {_0, _1568} + {_0, _2399};
  wire [1:0] _14562 = {_0, _5726} + {_0, _6814};
  wire [2:0] _14563 = {_0, _14561} + {_0, _14562};
  wire [1:0] _14564 = {_0, _9406} + {_0, _10527};
  wire [3:0] _14565 = {_0, _14563} + {_0, _0, _14564};
  wire _14566 = _12301 < _14565;
  wire _14567 = r1796 ^ _14566;
  wire _14568 = _12298 ? coded_block[1796] : r1796;
  wire _14569 = _12296 ? _14567 : _14568;
  always @ (posedge reset or posedge clock) if (reset) r1796 <= 1'd0; else if (_12300) r1796 <= _14569;
  wire [1:0] _14570 = {_0, _735} + {_0, _3997};
  wire [1:0] _14571 = {_0, _5534} + {_0, _6558};
  wire [2:0] _14572 = {_0, _14570} + {_0, _14571};
  wire [1:0] _14573 = {_0, _9375} + {_0, _10590};
  wire [3:0] _14574 = {_0, _14572} + {_0, _0, _14573};
  wire _14575 = _12301 < _14574;
  wire _14576 = r1795 ^ _14575;
  wire _14577 = _12298 ? coded_block[1795] : r1795;
  wire _14578 = _12296 ? _14576 : _14577;
  always @ (posedge reset or posedge clock) if (reset) r1795 <= 1'd0; else if (_12300) r1795 <= _14578;
  wire [1:0] _14579 = {_0, _1917} + {_0, _3646};
  wire [1:0] _14580 = {_0, _4447} + {_0, _7675};
  wire [2:0] _14581 = {_0, _14579} + {_0, _14580};
  wire [1:0] _14582 = {_0, _9248} + {_0, _11422};
  wire [3:0] _14583 = {_0, _14581} + {_0, _0, _14582};
  wire _14584 = _12301 < _14583;
  wire _14585 = r1794 ^ _14584;
  wire _14586 = _12298 ? coded_block[1794] : r1794;
  wire _14587 = _12296 ? _14585 : _14586;
  always @ (posedge reset or posedge clock) if (reset) r1794 <= 1'd0; else if (_12300) r1794 <= _14587;
  wire [1:0] _14588 = {_0, _735} + {_0, _3453};
  wire [1:0] _14589 = {_0, _6076} + {_0, _8059};
  wire [2:0] _14590 = {_0, _14588} + {_0, _14589};
  wire [1:0] _14591 = {_0, _9212} + {_0, _11933};
  wire [3:0] _14592 = {_0, _14590} + {_0, _0, _14591};
  wire _14593 = _12301 < _14592;
  wire _14594 = r1793 ^ _14593;
  wire _14595 = _12298 ? coded_block[1793] : r1793;
  wire _14596 = _12296 ? _14594 : _14595;
  always @ (posedge reset or posedge clock) if (reset) r1793 <= 1'd0; else if (_12300) r1793 <= _14596;
  wire [1:0] _14597 = {_0, _289} + {_0, _2941};
  wire [1:0] _14598 = {_0, _4223} + {_0, _6239};
  wire [2:0] _14599 = {_0, _14597} + {_0, _14598};
  wire [1:0] _14600 = {_0, _9118} + {_0, _11453};
  wire [3:0] _14601 = {_0, _14599} + {_0, _0, _14600};
  wire _14602 = _12301 < _14601;
  wire _14603 = r1792 ^ _14602;
  wire _14604 = _12298 ? coded_block[1792] : r1792;
  wire _14605 = _12296 ? _14603 : _14604;
  always @ (posedge reset or posedge clock) if (reset) r1792 <= 1'd0; else if (_12300) r1792 <= _14605;
  wire [1:0] _14606 = {_0, _1502} + {_0, _2399};
  wire [1:0] _14607 = {_0, _5373} + {_0, _7517};
  wire [2:0] _14608 = {_0, _14606} + {_0, _14607};
  wire [1:0] _14609 = {_0, _9022} + {_0, _11326};
  wire [3:0] _14610 = {_0, _14608} + {_0, _0, _14609};
  wire _14611 = _12301 < _14610;
  wire _14612 = r1791 ^ _14611;
  wire _14613 = _12298 ? coded_block[1791] : r1791;
  wire _14614 = _12296 ? _14612 : _14613;
  always @ (posedge reset or posedge clock) if (reset) r1791 <= 1'd0; else if (_12300) r1791 <= _14614;
  wire [1:0] _14615 = {_0, _1021} + {_0, _3870};
  wire [1:0] _14616 = {_0, _5183} + {_0, _6270};
  wire [2:0] _14617 = {_0, _14615} + {_0, _14616};
  wire [1:0] _14618 = {_0, _8863} + {_0, _11996};
  wire [3:0] _14619 = {_0, _14617} + {_0, _0, _14618};
  wire _14620 = _12301 < _14619;
  wire _14621 = r1790 ^ _14620;
  wire _14622 = _12298 ? coded_block[1790] : r1790;
  wire _14623 = _12296 ? _14621 : _14622;
  always @ (posedge reset or posedge clock) if (reset) r1790 <= 1'd0; else if (_12300) r1790 <= _14623;
  wire [1:0] _14624 = {_0, _1823} + {_0, _3933};
  wire [1:0] _14625 = {_0, _5022} + {_0, _7612};
  wire [2:0] _14626 = {_0, _14624} + {_0, _14625};
  wire [1:0] _14627 = {_0, _8736} + {_0, _11101};
  wire [3:0] _14628 = {_0, _14626} + {_0, _0, _14627};
  wire _14629 = _12301 < _14628;
  wire _14630 = r1789 ^ _14629;
  wire _14631 = _12298 ? coded_block[1789] : r1789;
  wire _14632 = _12296 ? _14630 : _14631;
  always @ (posedge reset or posedge clock) if (reset) r1789 <= 1'd0; else if (_12300) r1789 <= _14632;
  wire [1:0] _14633 = {_0, _289} + {_0, _2655};
  wire [1:0] _14634 = {_0, _4542} + {_0, _6176};
  wire [2:0] _14635 = {_0, _14633} + {_0, _14634};
  wire [1:0] _14636 = {_0, _8670} + {_0, _10910};
  wire [3:0] _14637 = {_0, _14635} + {_0, _0, _14636};
  wire _14638 = _12301 < _14637;
  wire _14639 = r1788 ^ _14638;
  wire _14640 = _12298 ? coded_block[1788] : r1788;
  wire _14641 = _12296 ? _14639 : _14640;
  always @ (posedge reset or posedge clock) if (reset) r1788 <= 1'd0; else if (_12300) r1788 <= _14641;
  wire [1:0] _14642 = {_0, _672} + {_0, _2112};
  wire [1:0] _14643 = {_0, _4319} + {_0, _8186};
  wire [2:0] _14644 = {_0, _14642} + {_0, _14643};
  wire [1:0] _14645 = {_0, _8607} + {_0, _11806};
  wire [3:0] _14646 = {_0, _14644} + {_0, _0, _14645};
  wire _14647 = _12301 < _14646;
  wire _14648 = r1787 ^ _14647;
  wire _14649 = _12298 ? coded_block[1787] : r1787;
  wire _14650 = _12296 ? _14648 : _14649;
  always @ (posedge reset or posedge clock) if (reset) r1787 <= 1'd0; else if (_12300) r1787 <= _14650;
  wire [1:0] _14651 = {_0, _576} + {_0, _2271};
  wire [1:0] _14652 = {_0, _5407} + {_0, _7773};
  wire [2:0] _14653 = {_0, _14651} + {_0, _14652};
  wire [1:0] _14654 = {_0, _8256} + {_0, _11677};
  wire [3:0] _14655 = {_0, _14653} + {_0, _0, _14654};
  wire _14656 = _12301 < _14655;
  wire _14657 = r1786 ^ _14656;
  wire _14658 = _12298 ? coded_block[1786] : r1786;
  wire _14659 = _12296 ? _14657 : _14658;
  always @ (posedge reset or posedge clock) if (reset) r1786 <= 1'd0; else if (_12300) r1786 <= _14659;
  wire [1:0] _14660 = {_0, _1758} + {_0, _3742};
  wire [1:0] _14661 = {_0, _4640} + {_0, _7965};
  wire [2:0] _14662 = {_0, _14660} + {_0, _14661};
  wire [1:0] _14663 = {_0, _9054} + {_0, _11644};
  wire [3:0] _14664 = {_0, _14662} + {_0, _0, _14663};
  wire _14665 = _12301 < _14664;
  wire _14666 = r1785 ^ _14665;
  wire _14667 = _12298 ? coded_block[1785] : r1785;
  wire _14668 = _12296 ? _14666 : _14667;
  always @ (posedge reset or posedge clock) if (reset) r1785 <= 1'd0; else if (_12300) r1785 <= _14668;
  wire [1:0] _14669 = {_0, _800} + {_0, _4028};
  wire [1:0] _14670 = {_0, _5183} + {_0, _7900};
  wire [2:0] _14671 = {_0, _14669} + {_0, _14670};
  wire [1:0] _14672 = {_0, _9534} + {_0, _11295};
  wire [3:0] _14673 = {_0, _14671} + {_0, _0, _14672};
  wire _14674 = _12301 < _14673;
  wire _14675 = r1784 ^ _14674;
  wire _14676 = _12298 ? coded_block[1784] : r1784;
  wire _14677 = _12296 ? _14675 : _14676;
  always @ (posedge reset or posedge clock) if (reset) r1784 <= 1'd0; else if (_12300) r1784 <= _14677;
  wire [1:0] _14678 = {_0, _2044} + {_0, _3390};
  wire [1:0] _14679 = {_0, _6045} + {_0, _7644};
  wire [2:0] _14680 = {_0, _14678} + {_0, _14679};
  wire [1:0] _14681 = {_0, _9311} + {_0, _10366};
  wire [3:0] _14682 = {_0, _14680} + {_0, _0, _14681};
  wire _14683 = _12301 < _14682;
  wire _14684 = r1783 ^ _14683;
  wire _14685 = _12298 ? coded_block[1783] : r1783;
  wire _14686 = _12296 ? _14684 : _14685;
  always @ (posedge reset or posedge clock) if (reset) r1783 <= 1'd0; else if (_12300) r1783 <= _14686;
  wire [1:0] _14687 = {_0, _1021} + {_0, _3580};
  wire [1:0] _14688 = {_0, _6108} + {_0, _7581};
  wire [2:0] _14689 = {_0, _14687} + {_0, _14688};
  wire [1:0] _14690 = {_0, _8926} + {_0, _10654};
  wire [3:0] _14691 = {_0, _14689} + {_0, _0, _14690};
  wire _14692 = _12301 < _14691;
  wire _14693 = r1782 ^ _14692;
  wire _14694 = _12298 ? coded_block[1782] : r1782;
  wire _14695 = _12296 ? _14693 : _14694;
  always @ (posedge reset or posedge clock) if (reset) r1782 <= 1'd0; else if (_12300) r1782 <= _14695;
  wire [1:0] _14696 = {_0, _958} + {_0, _3167};
  wire [1:0] _14697 = {_0, _4129} + {_0, _7293};
  wire [2:0] _14698 = {_0, _14696} + {_0, _14697};
  wire [1:0] _14699 = {_0, _9534} + {_0, _12219};
  wire [3:0] _14700 = {_0, _14698} + {_0, _0, _14699};
  wire _14701 = _12301 < _14700;
  wire _14702 = r1781 ^ _14701;
  wire _14703 = _12298 ? coded_block[1781] : r1781;
  wire _14704 = _12296 ? _14702 : _14703;
  always @ (posedge reset or posedge clock) if (reset) r1781 <= 1'd0; else if (_12300) r1781 <= _14704;
  wire [1:0] _14705 = {_0, _894} + {_0, _3870};
  wire [1:0] _14706 = {_0, _5310} + {_0, _7199};
  wire [2:0] _14707 = {_0, _14705} + {_0, _14706};
  wire [1:0] _14708 = {_0, _8225} + {_0, _11326};
  wire [3:0] _14709 = {_0, _14707} + {_0, _0, _14708};
  wire _14710 = _12301 < _14709;
  wire _14711 = r1780 ^ _14710;
  wire _14712 = _12298 ? coded_block[1780] : r1780;
  wire _14713 = _12296 ? _14711 : _14712;
  always @ (posedge reset or posedge clock) if (reset) r1780 <= 1'd0; else if (_12300) r1780 <= _14713;
  wire [1:0] _14714 = {_0, _2013} + {_0, _2239};
  wire [1:0] _14715 = {_0, _4478} + {_0, _7163};
  wire [2:0] _14716 = {_0, _14714} + {_0, _14715};
  wire [1:0] _14717 = {_0, _8957} + {_0, _12219};
  wire [3:0] _14718 = {_0, _14716} + {_0, _0, _14717};
  wire _14719 = _12301 < _14718;
  wire _14720 = r1779 ^ _14719;
  wire _14721 = _12298 ? coded_block[1779] : r1779;
  wire _14722 = _12296 ? _14720 : _14721;
  always @ (posedge reset or posedge clock) if (reset) r1779 <= 1'd0; else if (_12300) r1779 <= _14722;
  wire [1:0] _14723 = {_0, _479} + {_0, _3231};
  wire [1:0] _14724 = {_0, _4256} + {_0, _7069};
  wire [2:0] _14725 = {_0, _14723} + {_0, _14724};
  wire [1:0] _14726 = {_0, _8288} + {_0, _11869};
  wire [3:0] _14727 = {_0, _14725} + {_0, _0, _14726};
  wire _14728 = _12301 < _14727;
  wire _14729 = r1778 ^ _14728;
  wire _14730 = _12298 ? coded_block[1778] : r1778;
  wire _14731 = _12296 ? _14729 : _14730;
  always @ (posedge reset or posedge clock) if (reset) r1778 <= 1'd0; else if (_12300) r1778 <= _14731;
  wire [1:0] _14732 = {_0, _1631} + {_0, _2557};
  wire [1:0] _14733 = {_0, _4384} + {_0, _7005};
  wire [2:0] _14734 = {_0, _14732} + {_0, _14733};
  wire [1:0] _14735 = {_0, _8991} + {_0, _12155};
  wire [3:0] _14736 = {_0, _14734} + {_0, _0, _14735};
  wire _14737 = _12301 < _14736;
  wire _14738 = r1777 ^ _14737;
  wire _14739 = _12298 ? coded_block[1777] : r1777;
  wire _14740 = _12296 ? _14738 : _14739;
  always @ (posedge reset or posedge clock) if (reset) r1777 <= 1'd0; else if (_12300) r1777 <= _14740;
  wire [1:0] _14741 = {_0, _1726} + {_0, _2557};
  wire [1:0] _14742 = {_0, _5884} + {_0, _6973};
  wire [2:0] _14743 = {_0, _14741} + {_0, _14742};
  wire [1:0] _14744 = {_0, _9566} + {_0, _10685};
  wire [3:0] _14745 = {_0, _14743} + {_0, _0, _14744};
  wire _14746 = _12301 < _14745;
  wire _14747 = r1776 ^ _14746;
  wire _14748 = _12298 ? coded_block[1776] : r1776;
  wire _14749 = _12296 ? _14747 : _14748;
  always @ (posedge reset or posedge clock) if (reset) r1776 <= 1'd0; else if (_12300) r1776 <= _14749;
  wire [1:0] _14750 = {_0, _2013} + {_0, _2430};
  wire [1:0] _14751 = {_0, _5116} + {_0, _6908};
  wire [2:0] _14752 = {_0, _14750} + {_0, _14751};
  wire [1:0] _14753 = {_0, _10172} + {_0, _12282};
  wire [3:0] _14754 = {_0, _14752} + {_0, _0, _14753};
  wire _14755 = _12301 < _14754;
  wire _14756 = r1775 ^ _14755;
  wire _14757 = _12298 ? coded_block[1775] : r1775;
  wire _14758 = _12296 ? _14756 : _14757;
  always @ (posedge reset or posedge clock) if (reset) r1775 <= 1'd0; else if (_12300) r1775 <= _14758;
  wire [1:0] _14759 = {_0, _1917} + {_0, _3933};
  wire [1:0] _14760 = {_0, _6045} + {_0, _6877};
  wire [2:0] _14761 = {_0, _14759} + {_0, _14760};
  wire [1:0] _14762 = {_0, _9630} + {_0, _11581};
  wire [3:0] _14763 = {_0, _14761} + {_0, _0, _14762};
  wire _14764 = _12301 < _14763;
  wire _14765 = r1774 ^ _14764;
  wire _14766 = _12298 ? coded_block[1774] : r1774;
  wire _14767 = _12296 ? _14765 : _14766;
  always @ (posedge reset or posedge clock) if (reset) r1774 <= 1'd0; else if (_12300) r1774 <= _14767;
  wire [1:0] _14768 = {_0, _672} + {_0, _2239};
  wire [1:0] _14769 = {_0, _4192} + {_0, _6750};
  wire [2:0] _14770 = {_0, _14768} + {_0, _14769};
  wire [1:0] _14771 = {_0, _9661} + {_0, _10973};
  wire [3:0] _14772 = {_0, _14770} + {_0, _0, _14771};
  wire _14773 = _12301 < _14772;
  wire _14774 = r1773 ^ _14773;
  wire _14775 = _12298 ? coded_block[1773] : r1773;
  wire _14776 = _12296 ? _14774 : _14775;
  always @ (posedge reset or posedge clock) if (reset) r1773 <= 1'd0; else if (_12300) r1773 <= _14776;
  wire [1:0] _14777 = {_0, _639} + {_0, _2750};
  wire [1:0] _14778 = {_0, _5853} + {_0, _6431};
  wire [2:0] _14779 = {_0, _14777} + {_0, _14778};
  wire [1:0] _14780 = {_0, _9566} + {_0, _11933};
  wire [3:0] _14781 = {_0, _14779} + {_0, _0, _14780};
  wire _14782 = _12301 < _14781;
  wire _14783 = r1772 ^ _14782;
  wire _14784 = _12298 ? coded_block[1772] : r1772;
  wire _14785 = _12296 ? _14783 : _14784;
  always @ (posedge reset or posedge clock) if (reset) r1772 <= 1'd0; else if (_12300) r1772 <= _14785;
  wire [1:0] _14786 = {_0, _990} + {_0, _3933};
  wire [1:0] _14787 = {_0, _5757} + {_0, _6366};
  wire [2:0] _14788 = {_0, _14786} + {_0, _14787};
  wire [1:0] _14789 = {_0, _8352} + {_0, _11516};
  wire [3:0] _14790 = {_0, _14788} + {_0, _0, _14789};
  wire _14791 = _12301 < _14790;
  wire _14792 = r1771 ^ _14791;
  wire _14793 = _12298 ? coded_block[1771] : r1771;
  wire _14794 = _12296 ? _14792 : _14793;
  always @ (posedge reset or posedge clock) if (reset) r1771 <= 1'd0; else if (_12300) r1771 <= _14794;
  wire [1:0] _14795 = {_0, _672} + {_0, _2750};
  wire [1:0] _14796 = {_0, _5597} + {_0, _6334};
  wire [2:0] _14797 = {_0, _14795} + {_0, _14796};
  wire [1:0] _14798 = {_0, _8288} + {_0, _10846};
  wire [3:0] _14799 = {_0, _14797} + {_0, _0, _14798};
  wire _14800 = _12301 < _14799;
  wire _14801 = r1770 ^ _14800;
  wire _14802 = _12298 ? coded_block[1770] : r1770;
  wire _14803 = _12296 ? _14801 : _14802;
  always @ (posedge reset or posedge clock) if (reset) r1770 <= 1'd0; else if (_12300) r1770 <= _14803;
  wire [1:0] _14804 = {_0, _894} + {_0, _2557};
  wire [1:0] _14805 = {_0, _6139} + {_0, _6303};
  wire [2:0] _14806 = {_0, _14804} + {_0, _14805};
  wire [1:0] _14807 = {_0, _9693} + {_0, _10973};
  wire [3:0] _14808 = {_0, _14806} + {_0, _0, _14807};
  wire _14809 = _12301 < _14808;
  wire _14810 = r1769 ^ _14809;
  wire _14811 = _12298 ? coded_block[1769] : r1769;
  wire _14812 = _12296 ? _14810 : _14811;
  always @ (posedge reset or posedge clock) if (reset) r1769 <= 1'd0; else if (_12300) r1769 <= _14812;
  wire [1:0] _14813 = {_0, _1950} + {_0, _2750};
  wire [1:0] _14814 = {_0, _6012} + {_0, _8123};
  wire [2:0] _14815 = {_0, _14813} + {_0, _14814};
  wire [1:0] _14816 = {_0, _8957} + {_0, _11708};
  wire [3:0] _14817 = {_0, _14815} + {_0, _0, _14816};
  wire _14818 = _12301 < _14817;
  wire _14819 = r1768 ^ _14818;
  wire _14820 = _12298 ? coded_block[1768] : r1768;
  wire _14821 = _12296 ? _14819 : _14820;
  always @ (posedge reset or posedge clock) if (reset) r1768 <= 1'd0; else if (_12300) r1768 <= _14821;
  wire [1:0] _14822 = {_0, _1247} + {_0, _3517};
  wire [1:0] _14823 = {_0, _5918} + {_0, _6687};
  wire [2:0] _14824 = {_0, _14822} + {_0, _14823};
  wire [1:0] _14825 = {_0, _9342} + {_0, _10941};
  wire [3:0] _14826 = {_0, _14824} + {_0, _0, _14825};
  wire _14827 = _12301 < _14826;
  wire _14828 = r1767 ^ _14827;
  wire _14829 = _12298 ? coded_block[1767] : r1767;
  wire _14830 = _12296 ? _14828 : _14829;
  always @ (posedge reset or posedge clock) if (reset) r1767 <= 1'd0; else if (_12300) r1767 <= _14830;
  wire [1:0] _14831 = {_0, _831} + {_0, _3901};
  wire [1:0] _14832 = {_0, _5694} + {_0, _6942};
  wire [2:0] _14833 = {_0, _14831} + {_0, _14832};
  wire [1:0] _14834 = {_0, _9054} + {_0, _11900};
  wire [3:0] _14835 = {_0, _14833} + {_0, _0, _14834};
  wire _14836 = _12301 < _14835;
  wire _14837 = r1766 ^ _14836;
  wire _14838 = _12298 ? coded_block[1766] : r1766;
  wire _14839 = _12296 ? _14837 : _14838;
  always @ (posedge reset or posedge clock) if (reset) r1766 <= 1'd0; else if (_12300) r1766 <= _14839;
  wire [1:0] _14840 = {_0, _735} + {_0, _2813};
  wire [1:0] _14841 = {_0, _5663} + {_0, _6397};
  wire [2:0] _14842 = {_0, _14840} + {_0, _14841};
  wire [1:0] _14843 = {_0, _8352} + {_0, _10910};
  wire [3:0] _14844 = {_0, _14842} + {_0, _0, _14843};
  wire _14845 = _12301 < _14844;
  wire _14846 = r1765 ^ _14845;
  wire _14847 = _12298 ? coded_block[1765] : r1765;
  wire _14848 = _12296 ? _14846 : _14847;
  always @ (posedge reset or posedge clock) if (reset) r1765 <= 1'd0; else if (_12300) r1765 <= _14848;
  wire [1:0] _14849 = {_0, _383} + {_0, _4060};
  wire [1:0] _14850 = {_0, _5628} + {_0, _7804};
  wire [2:0] _14851 = {_0, _14849} + {_0, _14850};
  wire [1:0] _14852 = {_0, _9181} + {_0, _10462};
  wire [3:0] _14853 = {_0, _14851} + {_0, _0, _14852};
  wire _14854 = _12301 < _14853;
  wire _14855 = r1764 ^ _14854;
  wire _14856 = _12298 ? coded_block[1764] : r1764;
  wire _14857 = _12296 ? _14855 : _14856;
  always @ (posedge reset or posedge clock) if (reset) r1764 <= 1'd0; else if (_12300) r1764 <= _14857;
  wire [1:0] _14858 = {_0, _1568} + {_0, _2655};
  wire [1:0] _14859 = {_0, _5152} + {_0, _6558};
  wire [2:0] _14860 = {_0, _14858} + {_0, _14859};
  wire [1:0] _14861 = {_0, _9534} + {_0, _11677};
  wire [3:0] _14862 = {_0, _14860} + {_0, _0, _14861};
  wire _14863 = _12301 < _14862;
  wire _14864 = r1763 ^ _14863;
  wire _14865 = _12298 ? coded_block[1763] : r1763;
  wire _14866 = _12296 ? _14864 : _14865;
  always @ (posedge reset or posedge clock) if (reset) r1763 <= 1'd0; else if (_12300) r1763 <= _14866;
  wire [1:0] _14867 = {_0, _1406} + {_0, _2782};
  wire [1:0] _14868 = {_0, _5085} + {_0, _8028};
  wire [2:0] _14869 = {_0, _14867} + {_0, _14868};
  wire [1:0] _14870 = {_0, _9724} + {_0, _11996};
  wire [3:0] _14871 = {_0, _14869} + {_0, _0, _14870};
  wire _14872 = _12301 < _14871;
  wire _14873 = r1762 ^ _14872;
  wire _14874 = _12298 ? coded_block[1762] : r1762;
  wire _14875 = _12296 ? _14873 : _14874;
  always @ (posedge reset or posedge clock) if (reset) r1762 <= 1'd0; else if (_12300) r1762 <= _14875;
  wire [1:0] _14876 = {_0, _2044} + {_0, _2719};
  wire [1:0] _14877 = {_0, _5053} + {_0, _6494};
  wire [2:0] _14878 = {_0, _14876} + {_0, _14877};
  wire [1:0] _14879 = {_0, _8383} + {_0, _10272};
  wire [3:0] _14880 = {_0, _14878} + {_0, _0, _14879};
  wire _14881 = _12301 < _14880;
  wire _14882 = r1761 ^ _14881;
  wire _14883 = _12298 ? coded_block[1761] : r1761;
  wire _14884 = _12296 ? _14882 : _14883;
  always @ (posedge reset or posedge clock) if (reset) r1761 <= 1'd0; else if (_12300) r1761 <= _14884;
  wire [1:0] _14885 = {_0, _800} + {_0, _3933};
  wire [1:0] _14886 = {_0, _4989} + {_0, _7454};
  wire [2:0] _14887 = {_0, _14885} + {_0, _14886};
  wire [1:0] _14888 = {_0, _9980} + {_0, _11453};
  wire [3:0] _14889 = {_0, _14887} + {_0, _0, _14888};
  wire _14890 = _12301 < _14889;
  wire _14891 = r1760 ^ _14890;
  wire _14892 = _12298 ? coded_block[1760] : r1760;
  wire _14893 = _12296 ? _14891 : _14892;
  always @ (posedge reset or posedge clock) if (reset) r1760 <= 1'd0; else if (_12300) r1760 <= _14893;
  wire [1:0] _14894 = {_0, _831} + {_0, _2239};
  wire [1:0] _14895 = {_0, _4671} + {_0, _7868};
  wire [2:0] _14896 = {_0, _14894} + {_0, _14895};
  wire [1:0] _14897 = {_0, _9693} + {_0, _10303};
  wire [3:0] _14898 = {_0, _14896} + {_0, _0, _14897};
  wire _14899 = _12301 < _14898;
  wire _14900 = r1759 ^ _14899;
  wire _14901 = _12298 ? coded_block[1759] : r1759;
  wire _14902 = _12296 ? _14900 : _14901;
  always @ (posedge reset or posedge clock) if (reset) r1759 <= 1'd0; else if (_12300) r1759 <= _14902;
  wire [1:0] _14903 = {_0, _958} + {_0, _2399};
  wire [1:0] _14904 = {_0, _4605} + {_0, _6462};
  wire [2:0] _14905 = {_0, _14903} + {_0, _14904};
  wire [1:0] _14906 = {_0, _8894} + {_0, _12092};
  wire [3:0] _14907 = {_0, _14905} + {_0, _0, _14906};
  wire _14908 = _12301 < _14907;
  wire _14909 = r1758 ^ _14908;
  wire _14910 = _12298 ? coded_block[1758] : r1758;
  wire _14911 = _12296 ? _14909 : _14910;
  always @ (posedge reset or posedge clock) if (reset) r1758 <= 1'd0; else if (_12300) r1758 <= _14911;
  wire [1:0] _14912 = {_0, _1917} + {_0, _4060};
  wire [1:0] _14913 = {_0, _4511} + {_0, _7036};
  wire [2:0] _14914 = {_0, _14912} + {_0, _14913};
  wire [1:0] _14915 = {_0, _8511} + {_0, _11869};
  wire [3:0] _14916 = {_0, _14914} + {_0, _0, _14915};
  wire _14917 = _12301 < _14916;
  wire _14918 = r1757 ^ _14917;
  wire _14919 = _12298 ? coded_block[1757] : r1757;
  wire _14920 = _12296 ? _14918 : _14919;
  always @ (posedge reset or posedge clock) if (reset) r1757 <= 1'd0; else if (_12300) r1757 <= _14920;
  wire [1:0] _14921 = {_0, _1470} + {_0, _2782};
  wire [1:0] _14922 = {_0, _4160} + {_0, _7454};
  wire [2:0] _14923 = {_0, _14921} + {_0, _14922};
  wire [1:0] _14924 = {_0, _9469} + {_0, _10335};
  wire [3:0] _14925 = {_0, _14923} + {_0, _0, _14924};
  wire _14926 = _12301 < _14925;
  wire _14927 = r1756 ^ _14926;
  wire _14928 = _12298 ? coded_block[1756] : r1756;
  wire _14929 = _12296 ? _14927 : _14928;
  always @ (posedge reset or posedge clock) if (reset) r1756 <= 1'd0; else if (_12300) r1756 <= _14929;
  wire [1:0] _14930 = {_0, _1343} + {_0, _4091};
  wire [1:0] _14931 = {_0, _5116} + {_0, _7931};
  wire [2:0] _14932 = {_0, _14930} + {_0, _14931};
  wire [1:0] _14933 = {_0, _9149} + {_0, _10717};
  wire [3:0] _14934 = {_0, _14932} + {_0, _0, _14933};
  wire _14935 = _12301 < _14934;
  wire _14936 = r1755 ^ _14935;
  wire _14937 = _12298 ? coded_block[1755] : r1755;
  wire _14938 = _12296 ? _14936 : _14937;
  always @ (posedge reset or posedge clock) if (reset) r1755 <= 1'd0; else if (_12300) r1755 <= _14938;
  wire [1:0] _14939 = {_0, _766} + {_0, _3709};
  wire [1:0] _14940 = {_0, _5534} + {_0, _8155};
  wire [2:0] _14941 = {_0, _14939} + {_0, _14940};
  wire [1:0] _14942 = {_0, _10141} + {_0, _11295};
  wire [3:0] _14943 = {_0, _14941} + {_0, _0, _14942};
  wire _14944 = _12301 < _14943;
  wire _14945 = r1754 ^ _14944;
  wire _14946 = _12298 ? coded_block[1754] : r1754;
  wire _14947 = _12296 ? _14945 : _14946;
  always @ (posedge reset or posedge clock) if (reset) r1754 <= 1'd0; else if (_12300) r1754 <= _14947;
  wire [1:0] _14948 = {_0, _510} + {_0, _3615};
  wire [1:0] _14949 = {_0, _6108} + {_0, _7517};
  wire [2:0] _14950 = {_0, _14948} + {_0, _14949};
  wire [1:0] _14951 = {_0, _8480} + {_0, _10621};
  wire [3:0] _14952 = {_0, _14950} + {_0, _0, _14951};
  wire _14953 = _12301 < _14952;
  wire _14954 = r1753 ^ _14953;
  wire _14955 = _12298 ? coded_block[1753] : r1753;
  wire _14956 = _12296 ? _14954 : _14955;
  always @ (posedge reset or posedge clock) if (reset) r1753 <= 1'd0; else if (_12300) r1753 <= _14956;
  wire [1:0] _14957 = {_0, _1758} + {_0, _3549};
  wire [1:0] _14958 = {_0, _4734} + {_0, _6558};
  wire [2:0] _14959 = {_0, _14957} + {_0, _14958};
  wire [1:0] _14960 = {_0, _9181} + {_0, _11165};
  wire [3:0] _14961 = {_0, _14959} + {_0, _0, _14960};
  wire _14962 = _12301 < _14961;
  wire _14963 = r1752 ^ _14962;
  wire _14964 = _12298 ? coded_block[1752] : r1752;
  wire _14965 = _12296 ? _14963 : _14964;
  always @ (posedge reset or posedge clock) if (reset) r1752 <= 1'd0; else if (_12300) r1752 <= _14965;
  wire [1:0] _14966 = {_0, _1917} + {_0, _3486};
  wire [1:0] _14967 = {_0, _5438} + {_0, _7996};
  wire [2:0] _14968 = {_0, _14966} + {_0, _14967};
  wire [1:0] _14969 = {_0, _8894} + {_0, _12219};
  wire [3:0] _14970 = {_0, _14968} + {_0, _0, _14969};
  wire _14971 = _12301 < _14970;
  wire _14972 = r1751 ^ _14971;
  wire _14973 = _12298 ? coded_block[1751] : r1751;
  wire _14974 = _12296 ? _14972 : _14973;
  always @ (posedge reset or posedge clock) if (reset) r1751 <= 1'd0; else if (_12300) r1751 <= _14974;
  wire [1:0] _14975 = {_0, _447} + {_0, _3359};
  wire [1:0] _14976 = {_0, _4319} + {_0, _6462};
  wire [2:0] _14977 = {_0, _14975} + {_0, _14976};
  wire [1:0] _14978 = {_0, _9980} + {_0, _12282};
  wire [3:0] _14979 = {_0, _14977} + {_0, _0, _14978};
  wire _14980 = _12301 < _14979;
  wire _14981 = r1750 ^ _14980;
  wire _14982 = _12298 ? coded_block[1750] : r1750;
  wire _14983 = _12296 ? _14981 : _14982;
  always @ (posedge reset or posedge clock) if (reset) r1750 <= 1'd0; else if (_12300) r1750 <= _14983;
  wire [1:0] _14984 = {_0, _1406} + {_0, _3325};
  wire [1:0] _14985 = {_0, _4830} + {_0, _7132};
  wire [2:0] _14986 = {_0, _14984} + {_0, _14985};
  wire [1:0] _14987 = {_0, _10077} + {_0, _11771};
  wire [3:0] _14988 = {_0, _14986} + {_0, _0, _14987};
  wire _14989 = _12301 < _14988;
  wire _14990 = r1749 ^ _14989;
  wire _14991 = _12298 ? coded_block[1749] : r1749;
  wire _14992 = _12296 ? _14990 : _14991;
  always @ (posedge reset or posedge clock) if (reset) r1749 <= 1'd0; else if (_12300) r1749 <= _14992;
  wire [1:0] _14993 = {_0, _1343} + {_0, _3198};
  wire [1:0] _14994 = {_0, _6076} + {_0, _6397};
  wire [2:0] _14995 = {_0, _14993} + {_0, _14994};
  wire [1:0] _14996 = {_0, _9853} + {_0, _11740};
  wire [3:0] _14997 = {_0, _14995} + {_0, _0, _14996};
  wire _14998 = _12301 < _14997;
  wire _14999 = r1748 ^ _14998;
  wire _15000 = _12298 ? coded_block[1748] : r1748;
  wire _15001 = _12296 ? _14999 : _15000;
  always @ (posedge reset or posedge clock) if (reset) r1748 <= 1'd0; else if (_12300) r1748 <= _15001;
  wire [1:0] _15002 = {_0, _161} + {_0, _3135};
  wire [1:0] _15003 = {_0, _4574} + {_0, _6462};
  wire [2:0] _15004 = {_0, _15002} + {_0, _15003};
  wire [1:0] _15005 = {_0, _8225} + {_0, _10590};
  wire [3:0] _15006 = {_0, _15004} + {_0, _0, _15005};
  wire _15007 = _12301 < _15006;
  wire _15008 = r1747 ^ _15007;
  wire _15009 = _12298 ? coded_block[1747] : r1747;
  wire _15010 = _12296 ? _15008 : _15009;
  always @ (posedge reset or posedge clock) if (reset) r1747 <= 1'd0; else if (_12300) r1747 <= _15010;
  wire [1:0] _15011 = {_0, _1533} + {_0, _3068};
  wire [1:0] _15012 = {_0, _4478} + {_0, _7454};
  wire [2:0] _15013 = {_0, _15011} + {_0, _15012};
  wire [1:0] _15014 = {_0, _9597} + {_0, _11101};
  wire [3:0] _15015 = {_0, _15013} + {_0, _0, _15014};
  wire _15016 = _12301 < _15015;
  wire _15017 = r1746 ^ _15016;
  wire _15018 = _12298 ? coded_block[1746] : r1746;
  wire _15019 = _12296 ? _15017 : _15018;
  always @ (posedge reset or posedge clock) if (reset) r1746 <= 1'd0; else if (_12300) r1746 <= _15019;
  wire [1:0] _15020 = {_0, _1823} + {_0, _3005};
  wire [1:0] _15021 = {_0, _5183} + {_0, _6558};
  wire [2:0] _15022 = {_0, _15020} + {_0, _15021};
  wire [1:0] _15023 = {_0, _9853} + {_0, _11869};
  wire [3:0] _15024 = {_0, _15022} + {_0, _0, _15023};
  wire _15025 = _12301 < _15024;
  wire _15026 = r1745 ^ _15025;
  wire _15027 = _12298 ? coded_block[1745] : r1745;
  wire _15028 = _12296 ? _15026 : _15027;
  always @ (posedge reset or posedge clock) if (reset) r1745 <= 1'd0; else if (_12300) r1745 <= _15028;
  wire [1:0] _15029 = {_0, _1950} + {_0, _2974};
  wire [1:0] _15030 = {_0, _4447} + {_0, _7804};
  wire [2:0] _15031 = {_0, _15029} + {_0, _15030};
  wire [1:0] _15032 = {_0, _9534} + {_0, _11740};
  wire [3:0] _15033 = {_0, _15031} + {_0, _0, _15032};
  wire _15034 = _12301 < _15033;
  wire _15035 = r1744 ^ _15034;
  wire _15036 = _12298 ? coded_block[1744] : r1744;
  wire _15037 = _12296 ? _15035 : _15036;
  always @ (posedge reset or posedge clock) if (reset) r1744 <= 1'd0; else if (_12300) r1744 <= _15037;
  wire [1:0] _15038 = {_0, _1184} + {_0, _2526};
  wire [1:0] _15039 = {_0, _5183} + {_0, _6781};
  wire [2:0] _15040 = {_0, _15038} + {_0, _15039};
  wire [1:0] _15041 = {_0, _8446} + {_0, _11516};
  wire [3:0] _15042 = {_0, _15040} + {_0, _0, _15041};
  wire _15043 = _12301 < _15042;
  wire _15044 = r1743 ^ _15043;
  wire _15045 = _12298 ? coded_block[1743] : r1743;
  wire _15046 = _12296 ? _15044 : _15045;
  always @ (posedge reset or posedge clock) if (reset) r1743 <= 1'd0; else if (_12300) r1743 <= _15046;
  wire [1:0] _15047 = {_0, _1057} + {_0, _2463};
  wire [1:0] _15048 = {_0, _4895} + {_0, _8092};
  wire [2:0] _15049 = {_0, _15047} + {_0, _15048};
  wire [1:0] _15050 = {_0, _9917} + {_0, _10527};
  wire [3:0] _15051 = {_0, _15049} + {_0, _0, _15050};
  wire _15052 = _12301 < _15051;
  wire _15053 = r1742 ^ _15052;
  wire _15054 = _12298 ? coded_block[1742] : r1742;
  wire _15055 = _12296 ? _15053 : _15054;
  always @ (posedge reset or posedge clock) if (reset) r1742 <= 1'd0; else if (_12300) r1742 <= _15055;
  wire [1:0] _15056 = {_0, _1533} + {_0, _2208};
  wire [1:0] _15057 = {_0, _4542} + {_0, _7996};
  wire [2:0] _15058 = {_0, _15056} + {_0, _15057};
  wire [1:0] _15059 = {_0, _9886} + {_0, _10272};
  wire [3:0] _15060 = {_0, _15058} + {_0, _0, _15059};
  wire _15061 = _12301 < _15060;
  wire _15062 = r1741 ^ _15061;
  wire _15063 = _12298 ? coded_block[1741] : r1741;
  wire _15064 = _12296 ? _15062 : _15063;
  always @ (posedge reset or posedge clock) if (reset) r1741 <= 1'd0; else if (_12300) r1741 <= _15064;
  wire [1:0] _15065 = {_0, _1789} + {_0, _2081};
  wire [1:0] _15066 = {_0, _6076} + {_0, _6303};
  wire [2:0] _15067 = {_0, _15065} + {_0, _15066};
  wire [1:0] _15068 = {_0, _8991} + {_0, _10783};
  wire [3:0] _15069 = {_0, _15067} + {_0, _0, _15068};
  wire _15070 = _12301 < _15069;
  wire _15071 = r1740 ^ _15070;
  wire _15072 = _12298 ? coded_block[1740] : r1740;
  wire _15073 = _12296 ? _15071 : _15072;
  always @ (posedge reset or posedge clock) if (reset) r1740 <= 1'd0; else if (_12300) r1740 <= _15073;
  wire [1:0] _15074 = {_0, _1599} + {_0, _2367};
  wire [1:0] _15075 = {_0, _4734} + {_0, _7230};
  wire [2:0] _15076 = {_0, _15074} + {_0, _15075};
  wire [1:0] _15077 = {_0, _8638} + {_0, _11613};
  wire [3:0] _15078 = {_0, _15076} + {_0, _0, _15077};
  wire _15079 = _12301 < _15078;
  wire _15080 = r1739 ^ _15079;
  wire _15081 = _12298 ? coded_block[1739] : r1739;
  wire _15082 = _12296 ? _15080 : _15081;
  always @ (posedge reset or posedge clock) if (reset) r1739 <= 1'd0; else if (_12300) r1739 <= _15082;
  wire [1:0] _15083 = {_0, _1439} + {_0, _4028};
  wire [1:0] _15084 = {_0, _5790} + {_0, _6781};
  wire [2:0] _15085 = {_0, _15083} + {_0, _15084};
  wire [1:0] _15086 = {_0, _8319} + {_0, _11358};
  wire [3:0] _15087 = {_0, _15085} + {_0, _0, _15086};
  wire _15088 = _12301 < _15087;
  wire _15089 = r1738 ^ _15088;
  wire _15090 = _12298 ? coded_block[1738] : r1738;
  wire _15091 = _12296 ? _15089 : _15090;
  always @ (posedge reset or posedge clock) if (reset) r1738 <= 1'd0; else if (_12300) r1738 <= _15091;
  wire [1:0] _15092 = {_0, _1375} + {_0, _3646};
  wire [1:0] _15093 = {_0, _6045} + {_0, _6814};
  wire [2:0] _15094 = {_0, _15092} + {_0, _15093};
  wire [1:0] _15095 = {_0, _9469} + {_0, _11069};
  wire [3:0] _15096 = {_0, _15094} + {_0, _0, _15095};
  wire _15097 = _12301 < _15096;
  wire _15098 = r1737 ^ _15097;
  wire _15099 = _12298 ? coded_block[1737] : r1737;
  wire _15100 = _12296 ? _15098 : _15099;
  always @ (posedge reset or posedge clock) if (reset) r1737 <= 1'd0; else if (_12300) r1737 <= _15100;
  wire [1:0] _15101 = {_0, _1278} + {_0, _3678};
  wire [1:0] _15102 = {_0, _5597} + {_0, _7996};
  wire [2:0] _15103 = {_0, _15101} + {_0, _15102};
  wire [1:0] _15104 = {_0, _8767} + {_0, _11422};
  wire [3:0] _15105 = {_0, _15103} + {_0, _0, _15104};
  wire _15106 = _12301 < _15105;
  wire _15107 = r1736 ^ _15106;
  wire _15108 = _12298 ? coded_block[1736] : r1736;
  wire _15109 = _12296 ? _15107 : _15108;
  always @ (posedge reset or posedge clock) if (reset) r1736 <= 1'd0; else if (_12300) r1736 <= _15109;
  wire [1:0] _15110 = {_0, _1215} + {_0, _3104};
  wire [1:0] _15111 = {_0, _5116} + {_0, _7996};
  wire [2:0] _15112 = {_0, _15110} + {_0, _15111};
  wire [1:0] _15113 = {_0, _8319} + {_0, _11771};
  wire [3:0] _15114 = {_0, _15112} + {_0, _0, _15113};
  wire _15115 = _12301 < _15114;
  wire _15116 = r1735 ^ _15115;
  wire _15117 = _12298 ? coded_block[1735] : r1735;
  wire _15118 = _12296 ? _15116 : _15117;
  always @ (posedge reset or posedge clock) if (reset) r1735 <= 1'd0; else if (_12300) r1735 <= _15118;
  wire [1:0] _15119 = {_0, _1151} + {_0, _3517};
  wire [1:0] _15120 = {_0, _5407} + {_0, _6176};
  wire [2:0] _15121 = {_0, _15119} + {_0, _15120};
  wire [1:0] _15122 = {_0, _9534} + {_0, _11771};
  wire [3:0] _15123 = {_0, _15121} + {_0, _0, _15122};
  wire _15124 = _12301 < _15123;
  wire _15125 = r1734 ^ _15124;
  wire _15126 = _12298 ? coded_block[1734] : r1734;
  wire _15127 = _12296 ? _15125 : _15126;
  always @ (posedge reset or posedge clock) if (reset) r1734 <= 1'd0; else if (_12300) r1734 <= _15127;
  wire [1:0] _15128 = {_0, _1088} + {_0, _2941};
  wire [1:0] _15129 = {_0, _5821} + {_0, _8155};
  wire [2:0] _15130 = {_0, _15128} + {_0, _15129};
  wire [1:0] _15131 = {_0, _9597} + {_0, _11485};
  wire [3:0] _15132 = {_0, _15130} + {_0, _0, _15131};
  wire _15133 = _12301 < _15132;
  wire _15134 = r1733 ^ _15133;
  wire _15135 = _12298 ? coded_block[1733] : r1733;
  wire _15136 = _12296 ? _15134 : _15135;
  always @ (posedge reset or posedge clock) if (reset) r1733 <= 1'd0; else if (_12300) r1733 <= _15136;
  wire [1:0] _15137 = {_0, _927} + {_0, _3517};
  wire [1:0] _15138 = {_0, _5279} + {_0, _6270};
  wire [2:0] _15139 = {_0, _15137} + {_0, _15138};
  wire [1:0] _15140 = {_0, _9822} + {_0, _10846};
  wire [3:0] _15141 = {_0, _15139} + {_0, _0, _15140};
  wire _15142 = _12301 < _15141;
  wire _15143 = r1732 ^ _15142;
  wire _15144 = _12298 ? coded_block[1732] : r1732;
  wire _15145 = _12296 ? _15143 : _15144;
  always @ (posedge reset or posedge clock) if (reset) r1732 <= 1'd0; else if (_12300) r1732 <= _15145;
  wire [1:0] _15146 = {_0, _863} + {_0, _2813};
  wire [1:0] _15147 = {_0, _4415} + {_0, _8092};
  wire [2:0] _15148 = {_0, _15146} + {_0, _15147};
  wire [1:0] _15149 = {_0, _9149} + {_0, _11613};
  wire [3:0] _15150 = {_0, _15148} + {_0, _0, _15149};
  wire _15151 = _12301 < _15150;
  wire _15152 = r1731 ^ _15151;
  wire _15153 = _12298 ? coded_block[1731] : r1731;
  wire _15154 = _12296 ? _15152 : _15153;
  always @ (posedge reset or posedge clock) if (reset) r1731 <= 1'd0; else if (_12300) r1731 <= _15154;
  wire [1:0] _15155 = {_0, _608} + {_0, _2592};
  wire [1:0] _15156 = {_0, _5501} + {_0, _6814};
  wire [2:0] _15157 = {_0, _15155} + {_0, _15156};
  wire [1:0] _15158 = {_0, _9917} + {_0, _10493};
  wire [3:0] _15159 = {_0, _15157} + {_0, _0, _15158};
  wire _15160 = _12301 < _15159;
  wire _15161 = r1730 ^ _15160;
  wire _15162 = _12298 ? coded_block[1730] : r1730;
  wire _15163 = _12296 ? _15161 : _15162;
  always @ (posedge reset or posedge clock) if (reset) r1730 <= 1'd0; else if (_12300) r1730 <= _15163;
  wire [1:0] _15164 = {_0, _416} + {_0, _3453};
  wire [1:0] _15165 = {_0, _4926} + {_0, _6270};
  wire [2:0] _15166 = {_0, _15164} + {_0, _15165};
  wire [1:0] _15167 = {_0, _10014} + {_0, _12219};
  wire [3:0] _15168 = {_0, _15166} + {_0, _0, _15167};
  wire _15169 = _12301 < _15168;
  wire _15170 = r1729 ^ _15169;
  wire _15171 = _12298 ? coded_block[1729] : r1729;
  wire _15172 = _12296 ? _15170 : _15171;
  always @ (posedge reset or posedge clock) if (reset) r1729 <= 1'd0; else if (_12300) r1729 <= _15172;
  wire [1:0] _15173 = {_0, _320} + {_0, _3646};
  wire [1:0] _15174 = {_0, _5022} + {_0, _6303};
  wire [2:0] _15175 = {_0, _15173} + {_0, _15174};
  wire [1:0] _15176 = {_0, _8319} + {_0, _11196};
  wire [3:0] _15177 = {_0, _15175} + {_0, _0, _15176};
  wire _15178 = _12301 < _15177;
  wire _15179 = r1728 ^ _15178;
  wire _15180 = _12298 ? coded_block[1728] : r1728;
  wire _15181 = _12296 ? _15179 : _15180;
  always @ (posedge reset or posedge clock) if (reset) r1728 <= 1'd0; else if (_12300) r1728 <= _15181;
  wire [1:0] _15182 = {_0, _255} + {_0, _2557};
  wire [1:0] _15183 = {_0, _5565} + {_0, _7100};
  wire [2:0] _15184 = {_0, _15182} + {_0, _15183};
  wire [1:0] _15185 = {_0, _10141} + {_0, _10941};
  wire [3:0] _15186 = {_0, _15184} + {_0, _0, _15185};
  wire _15187 = _12301 < _15186;
  wire _15188 = r1727 ^ _15187;
  wire _15189 = _12298 ? coded_block[1727] : r1727;
  wire _15190 = _12296 ? _15188 : _15189;
  always @ (posedge reset or posedge clock) if (reset) r1727 <= 1'd0; else if (_12300) r1727 <= _15190;
  wire [1:0] _15191 = {_0, _224} + {_0, _3870};
  wire [1:0] _15192 = {_0, _4798} + {_0, _6494};
  wire [2:0] _15193 = {_0, _15191} + {_0, _15192};
  wire [1:0] _15194 = {_0, _8767} + {_0, _10685};
  wire [3:0] _15195 = {_0, _15193} + {_0, _0, _15194};
  wire _15196 = _12301 < _15195;
  wire _15197 = r1726 ^ _15196;
  wire _15198 = _12298 ? coded_block[1726] : r1726;
  wire _15199 = _12296 ? _15197 : _15198;
  always @ (posedge reset or posedge clock) if (reset) r1726 <= 1'd0; else if (_12300) r1726 <= _15199;
  wire [1:0] _15200 = {_0, _192} + {_0, _2878};
  wire [1:0] _15201 = {_0, _5215} + {_0, _6652};
  wire [2:0] _15202 = {_0, _15200} + {_0, _15201};
  wire [1:0] _15203 = {_0, _8543} + {_0, _10272};
  wire [3:0] _15204 = {_0, _15202} + {_0, _0, _15203};
  wire _15205 = _12301 < _15204;
  wire _15206 = r1725 ^ _15205;
  wire _15207 = _12298 ? coded_block[1725] : r1725;
  wire _15208 = _12296 ? _15206 : _15207;
  always @ (posedge reset or posedge clock) if (reset) r1725 <= 1'd0; else if (_12300) r1725 <= _15208;
  wire [1:0] _15209 = {_0, _34} + {_0, _2336};
  wire [1:0] _15210 = {_0, _4415} + {_0, _6494};
  wire [2:0] _15211 = {_0, _15209} + {_0, _15210};
  wire [1:0] _15212 = {_0, _8574} + {_0, _10654};
  wire [3:0] _15213 = {_0, _15211} + {_0, _0, _15212};
  wire _15214 = _12301 < _15213;
  wire _15215 = r1724 ^ _15214;
  wire _15216 = _12298 ? coded_block[1724] : r1724;
  wire _15217 = _12296 ? _15215 : _15216;
  always @ (posedge reset or posedge clock) if (reset) r1724 <= 1'd0; else if (_12300) r1724 <= _15217;
  wire [1:0] _15218 = {_0, _1854} + {_0, _3901};
  wire [1:0] _15219 = {_0, _5949} + {_0, _7996};
  wire [2:0] _15220 = {_0, _15218} + {_0, _15219};
  wire [1:0] _15221 = {_0, _10045} + {_0, _12092};
  wire [3:0] _15222 = {_0, _15220} + {_0, _0, _15221};
  wire _15223 = _12301 < _15222;
  wire _15224 = r1723 ^ _15223;
  wire _15225 = _12298 ? coded_block[1723] : r1723;
  wire _15226 = _12296 ? _15224 : _15225;
  always @ (posedge reset or posedge clock) if (reset) r1723 <= 1'd0; else if (_12300) r1723 <= _15226;
  wire [1:0] _15227 = {_0, _1917} + {_0, _3964};
  wire [1:0] _15228 = {_0, _6012} + {_0, _8059};
  wire [2:0] _15229 = {_0, _15227} + {_0, _15228};
  wire [1:0] _15230 = {_0, _10108} + {_0, _12155};
  wire [3:0] _15231 = {_0, _15229} + {_0, _0, _15230};
  wire _15232 = _12301 < _15231;
  wire _15233 = r1722 ^ _15232;
  wire _15234 = _12298 ? coded_block[1722] : r1722;
  wire _15235 = _12296 ? _15233 : _15234;
  always @ (posedge reset or posedge clock) if (reset) r1722 <= 1'd0; else if (_12300) r1722 <= _15235;
  wire [1:0] _15236 = {_0, _1950} + {_0, _3997};
  wire [1:0] _15237 = {_0, _6045} + {_0, _8092};
  wire [2:0] _15238 = {_0, _15236} + {_0, _15237};
  wire [1:0] _15239 = {_0, _10141} + {_0, _12188};
  wire [3:0] _15240 = {_0, _15238} + {_0, _0, _15239};
  wire _15241 = _12301 < _15240;
  wire _15242 = r1721 ^ _15241;
  wire _15243 = _12298 ? coded_block[1721] : r1721;
  wire _15244 = _12296 ? _15242 : _15243;
  always @ (posedge reset or posedge clock) if (reset) r1721 <= 1'd0; else if (_12300) r1721 <= _15244;
  wire [1:0] _15245 = {_0, _2013} + {_0, _4060};
  wire [1:0] _15246 = {_0, _6108} + {_0, _8155};
  wire [2:0] _15247 = {_0, _15245} + {_0, _15246};
  wire [1:0] _15248 = {_0, _10204} + {_0, _12251};
  wire [3:0] _15249 = {_0, _15247} + {_0, _0, _15248};
  wire _15250 = _12301 < _15249;
  wire _15251 = r1720 ^ _15250;
  wire _15252 = _12298 ? coded_block[1720] : r1720;
  wire _15253 = _12296 ? _15251 : _15252;
  always @ (posedge reset or posedge clock) if (reset) r1720 <= 1'd0; else if (_12300) r1720 <= _15253;
  wire [1:0] _15254 = {_0, _1981} + {_0, _4028};
  wire [1:0] _15255 = {_0, _6076} + {_0, _8123};
  wire [2:0] _15256 = {_0, _15254} + {_0, _15255};
  wire [1:0] _15257 = {_0, _10172} + {_0, _12219};
  wire [3:0] _15258 = {_0, _15256} + {_0, _0, _15257};
  wire _15259 = _12301 < _15258;
  wire _15260 = r1719 ^ _15259;
  wire _15261 = _12298 ? coded_block[1719] : r1719;
  wire _15262 = _12296 ? _15260 : _15261;
  always @ (posedge reset or posedge clock) if (reset) r1719 <= 1'd0; else if (_12300) r1719 <= _15262;
  wire [1:0] _15263 = {_0, _34} + {_0, _2112};
  wire [1:0] _15264 = {_0, _4192} + {_0, _6270};
  wire [2:0] _15265 = {_0, _15263} + {_0, _15264};
  wire [1:0] _15266 = {_0, _8352} + {_0, _10430};
  wire [3:0] _15267 = {_0, _15265} + {_0, _0, _15266};
  wire _15268 = _12301 < _15267;
  wire _15269 = r1718 ^ _15268;
  wire _15270 = _12298 ? coded_block[1718] : r1718;
  wire _15271 = _12296 ? _15269 : _15270;
  always @ (posedge reset or posedge clock) if (reset) r1718 <= 1'd0; else if (_12300) r1718 <= _15271;
  wire [1:0] _15272 = {_0, _1312} + {_0, _3486};
  wire [1:0] _15273 = {_0, _5757} + {_0, _7675};
  wire [2:0] _15274 = {_0, _15272} + {_0, _15273};
  wire [1:0] _15275 = {_0, _10077} + {_0, _10846};
  wire [3:0] _15276 = {_0, _15274} + {_0, _0, _15275};
  wire _15277 = _12301 < _15276;
  wire _15278 = r1717 ^ _15277;
  wire _15279 = _12298 ? coded_block[1717] : r1717;
  wire _15280 = _12296 ? _15278 : _15279;
  always @ (posedge reset or posedge clock) if (reset) r1717 <= 1'd0; else if (_12300) r1717 <= _15280;
  wire [1:0] _15281 = {_0, _1343} + {_0, _3870};
  wire [1:0] _15282 = {_0, _5565} + {_0, _7837};
  wire [2:0] _15283 = {_0, _15281} + {_0, _15282};
  wire [1:0] _15284 = {_0, _9759} + {_0, _12155};
  wire [3:0] _15285 = {_0, _15283} + {_0, _0, _15284};
  wire _15286 = _12301 < _15285;
  wire _15287 = r1716 ^ _15286;
  wire _15288 = _12298 ? coded_block[1716] : r1716;
  wire _15289 = _12296 ? _15287 : _15288;
  always @ (posedge reset or posedge clock) if (reset) r1716 <= 1'd0; else if (_12300) r1716 <= _15289;
  wire [1:0] _15290 = {_0, _1375} + {_0, _3005};
  wire [1:0] _15291 = {_0, _5949} + {_0, _7644};
  wire [2:0] _15292 = {_0, _15290} + {_0, _15291};
  wire [1:0] _15293 = {_0, _9917} + {_0, _11837};
  wire [3:0] _15294 = {_0, _15292} + {_0, _0, _15293};
  wire _15295 = _12301 < _15294;
  wire _15296 = r1715 ^ _15295;
  wire _15297 = _12298 ? coded_block[1715] : r1715;
  wire _15298 = _12296 ? _15296 : _15297;
  always @ (posedge reset or posedge clock) if (reset) r1715 <= 1'd0; else if (_12300) r1715 <= _15298;
  wire [1:0] _15299 = {_0, _1439} + {_0, _3359};
  wire [1:0] _15300 = {_0, _4861} + {_0, _7163};
  wire [2:0] _15301 = {_0, _15299} + {_0, _15300};
  wire [1:0] _15302 = {_0, _10108} + {_0, _11806};
  wire [3:0] _15303 = {_0, _15301} + {_0, _0, _15302};
  wire _15304 = _12301 < _15303;
  wire _15305 = r1714 ^ _15304;
  wire _15306 = _12298 ? coded_block[1714] : r1714;
  wire _15307 = _12296 ? _15305 : _15306;
  always @ (posedge reset or posedge clock) if (reset) r1714 <= 1'd0; else if (_12300) r1714 <= _15307;
  wire [1:0] _15308 = {_0, _1470} + {_0, _3294};
  wire [1:0] _15309 = {_0, _5438} + {_0, _6942};
  wire [2:0] _15310 = {_0, _15308} + {_0, _15309};
  wire [1:0] _15311 = {_0, _9248} + {_0, _12188};
  wire [3:0] _15312 = {_0, _15310} + {_0, _0, _15311};
  wire _15313 = _12301 < _15312;
  wire _15314 = r1713 ^ _15313;
  wire _15315 = _12298 ? coded_block[1713] : r1713;
  wire _15316 = _12296 ? _15314 : _15315;
  always @ (posedge reset or posedge clock) if (reset) r1713 <= 1'd0; else if (_12300) r1713 <= _15316;
  wire [1:0] _15317 = {_0, _1631} + {_0, _3325};
  wire [1:0] _15318 = {_0, _4447} + {_0, _6814};
  wire [2:0] _15319 = {_0, _15317} + {_0, _15318};
  wire [1:0] _15320 = {_0, _9311} + {_0, _10717};
  wire [3:0] _15321 = {_0, _15319} + {_0, _0, _15320};
  wire _15322 = _12301 < _15321;
  wire _15323 = r1712 ^ _15322;
  wire _15324 = _12298 ? coded_block[1712] : r1712;
  wire _15325 = _12296 ? _15323 : _15324;
  always @ (posedge reset or posedge clock) if (reset) r1712 <= 1'd0; else if (_12300) r1712 <= _15325;
  wire [1:0] _15326 = {_0, _1695} + {_0, _3805};
  wire [1:0] _15327 = {_0, _4895} + {_0, _7485};
  wire [2:0] _15328 = {_0, _15326} + {_0, _15327};
  wire [1:0] _15329 = {_0, _8607} + {_0, _10973};
  wire [3:0] _15330 = {_0, _15328} + {_0, _0, _15329};
  wire _15331 = _12301 < _15330;
  wire _15332 = r1711 ^ _15331;
  wire _15333 = _12298 ? coded_block[1711] : r1711;
  wire _15334 = _12296 ? _15332 : _15333;
  always @ (posedge reset or posedge clock) if (reset) r1711 <= 1'd0; else if (_12300) r1711 <= _15334;
  wire [1:0] _15335 = {_0, _1789} + {_0, _3262};
  wire [1:0] _15336 = {_0, _5821} + {_0, _6718};
  wire [2:0] _15337 = {_0, _15335} + {_0, _15336};
  wire [1:0] _15338 = {_0, _10045} + {_0, _11132};
  wire [3:0] _15339 = {_0, _15337} + {_0, _0, _15338};
  wire _15340 = _12301 < _15339;
  wire _15341 = r1710 ^ _15340;
  wire _15342 = _12298 ? coded_block[1710] : r1710;
  wire _15343 = _12296 ? _15341 : _15342;
  always @ (posedge reset or posedge clock) if (reset) r1710 <= 1'd0; else if (_12300) r1710 <= _15343;
  wire [1:0] _15344 = {_0, _1823} + {_0, _3390};
  wire [1:0] _15345 = {_0, _5342} + {_0, _7900};
  wire [2:0] _15346 = {_0, _15344} + {_0, _15345};
  wire [1:0] _15347 = {_0, _8799} + {_0, _12124};
  wire [3:0] _15348 = {_0, _15346} + {_0, _0, _15347};
  wire _15349 = _12301 < _15348;
  wire _15350 = r1709 ^ _15349;
  wire _15351 = _12298 ? coded_block[1709] : r1709;
  wire _15352 = _12296 ? _15350 : _15351;
  always @ (posedge reset or posedge clock) if (reset) r1709 <= 1'd0; else if (_12300) r1709 <= _15352;
  wire [1:0] _15353 = {_0, _2044} + {_0, _2271};
  wire [1:0] _15354 = {_0, _4511} + {_0, _7199};
  wire [2:0] _15355 = {_0, _15353} + {_0, _15354};
  wire [1:0] _15356 = {_0, _8991} + {_0, _12251};
  wire [3:0] _15357 = {_0, _15355} + {_0, _0, _15356};
  wire _15358 = _12301 < _15357;
  wire _15359 = r1708 ^ _15358;
  wire _15360 = _12298 ? coded_block[1708] : r1708;
  wire _15361 = _12296 ? _15359 : _15360;
  always @ (posedge reset or posedge clock) if (reset) r1708 <= 1'd0; else if (_12300) r1708 <= _15361;
  wire [1:0] _15362 = {_0, _97} + {_0, _2302};
  wire [1:0] _15363 = {_0, _4129} + {_0, _6431};
  wire [2:0] _15364 = {_0, _15362} + {_0, _15363};
  wire [1:0] _15365 = {_0, _8670} + {_0, _11358};
  wire [3:0] _15366 = {_0, _15364} + {_0, _0, _15365};
  wire _15367 = _12301 < _15366;
  wire _15368 = r1707 ^ _15367;
  wire _15369 = _12298 ? coded_block[1707] : r1707;
  wire _15370 = _12296 ? _15368 : _15369;
  always @ (posedge reset or posedge clock) if (reset) r1707 <= 1'd0; else if (_12300) r1707 <= _15370;
  wire [1:0] _15371 = {_0, _224} + {_0, _4091};
  wire [1:0] _15372 = {_0, _4958} + {_0, _7293};
  wire [2:0] _15373 = {_0, _15371} + {_0, _15372};
  wire [1:0] _15374 = {_0, _8736} + {_0, _10621};
  wire [3:0] _15375 = {_0, _15373} + {_0, _0, _15374};
  wire _15376 = _12301 < _15375;
  wire _15377 = r1706 ^ _15376;
  wire _15378 = _12298 ? coded_block[1706] : r1706;
  wire _15379 = _12296 ? _15377 : _15378;
  always @ (posedge reset or posedge clock) if (reset) r1706 <= 1'd0; else if (_12300) r1706 <= _15379;
  wire [1:0] _15380 = {_0, _255} + {_0, _2144};
  wire [1:0] _15381 = {_0, _4160} + {_0, _7036};
  wire [2:0] _15382 = {_0, _15380} + {_0, _15381};
  wire [1:0] _15383 = {_0, _9375} + {_0, _10814};
  wire [3:0] _15384 = {_0, _15382} + {_0, _0, _15383};
  wire _15385 = _12301 < _15384;
  wire _15386 = r1705 ^ _15385;
  wire _15387 = _12298 ? coded_block[1705] : r1705;
  wire _15388 = _12296 ? _15386 : _15387;
  always @ (posedge reset or posedge clock) if (reset) r1705 <= 1'd0; else if (_12300) r1705 <= _15388;
  wire [1:0] _15389 = {_0, _352} + {_0, _3549};
  wire [1:0] _15390 = {_0, _5726} + {_0, _7100};
  wire [2:0] _15391 = {_0, _15389} + {_0, _15390};
  wire [1:0] _15392 = {_0, _8383} + {_0, _10399};
  wire [3:0] _15393 = {_0, _15391} + {_0, _0, _15392};
  wire _15394 = _12301 < _15393;
  wire _15395 = r1704 ^ _15394;
  wire _15396 = _12298 ? coded_block[1704] : r1704;
  wire _15397 = _12296 ? _15395 : _15396;
  always @ (posedge reset or posedge clock) if (reset) r1704 <= 1'd0; else if (_12300) r1704 <= _15397;
  wire [1:0] _15398 = {_0, _416} + {_0, _2910};
  wire [1:0] _15399 = {_0, _6139} + {_0, _7710};
  wire [2:0] _15400 = {_0, _15398} + {_0, _15399};
  wire [1:0] _15401 = {_0, _9886} + {_0, _11259};
  wire [3:0] _15402 = {_0, _15400} + {_0, _0, _15401};
  wire _15403 = _12301 < _15402;
  wire _15404 = r1703 ^ _15403;
  wire _15405 = _12298 ? coded_block[1703] : r1703;
  wire _15406 = _12296 ? _15404 : _15405;
  always @ (posedge reset or posedge clock) if (reset) r1703 <= 1'd0; else if (_12300) r1703 <= _15406;
  wire [1:0] _15407 = {_0, _447} + {_0, _2175};
  wire [1:0] _15408 = {_0, _4989} + {_0, _6207};
  wire [2:0] _15409 = {_0, _15407} + {_0, _15408};
  wire [1:0] _15410 = {_0, _9790} + {_0, _11964};
  wire [3:0] _15411 = {_0, _15409} + {_0, _0, _15410};
  wire _15412 = _12301 < _15411;
  wire _15413 = r1702 ^ _15412;
  wire _15414 = _12298 ? coded_block[1702] : r1702;
  wire _15415 = _12296 ? _15413 : _15414;
  always @ (posedge reset or posedge clock) if (reset) r1702 <= 1'd0; else if (_12300) r1702 <= _15415;
  wire [1:0] _15416 = {_0, _510} + {_0, _3773};
  wire [1:0] _15417 = {_0, _5310} + {_0, _6334};
  wire [2:0] _15418 = {_0, _15416} + {_0, _15417};
  wire [1:0] _15419 = {_0, _9149} + {_0, _10366};
  wire [3:0] _15420 = {_0, _15418} + {_0, _0, _15419};
  wire _15421 = _12301 < _15420;
  wire _15422 = r1701 ^ _15421;
  wire _15423 = _12298 ? coded_block[1701] : r1701;
  wire _15424 = _12296 ? _15422 : _15423;
  always @ (posedge reset or posedge clock) if (reset) r1701 <= 1'd0; else if (_12300) r1701 <= _15424;
  wire [1:0] _15425 = {_0, _545} + {_0, _2847};
  wire [1:0] _15426 = {_0, _5853} + {_0, _7389};
  wire [2:0] _15427 = {_0, _15425} + {_0, _15426};
  wire [1:0] _15428 = {_0, _8415} + {_0, _11228};
  wire [3:0] _15429 = {_0, _15427} + {_0, _0, _15428};
  wire _15430 = _12301 < _15429;
  wire _15431 = r1700 ^ _15430;
  wire _15432 = _12298 ? coded_block[1700] : r1700;
  wire _15433 = _12296 ? _15431 : _15432;
  always @ (posedge reset or posedge clock) if (reset) r1700 <= 1'd0; else if (_12300) r1700 <= _15433;
  wire [1:0] _15434 = {_0, _576} + {_0, _3167};
  wire [1:0] _15435 = {_0, _4926} + {_0, _7931};
  wire [2:0] _15436 = {_0, _15434} + {_0, _15435};
  wire [1:0] _15437 = {_0, _9469} + {_0, _10493};
  wire [3:0] _15438 = {_0, _15436} + {_0, _0, _15437};
  wire _15439 = _12301 < _15438;
  wire _15440 = r1699 ^ _15439;
  wire _15441 = _12298 ? coded_block[1699] : r1699;
  wire _15442 = _12296 ? _15440 : _15441;
  always @ (posedge reset or posedge clock) if (reset) r1699 <= 1'd0; else if (_12300) r1699 <= _15442;
  wire [1:0] _15443 = {_0, _608} + {_0, _3615};
  wire [1:0] _15444 = {_0, _5246} + {_0, _7005};
  wire [2:0] _15445 = {_0, _15443} + {_0, _15444};
  wire [1:0] _15446 = {_0, _10014} + {_0, _11550};
  wire [3:0] _15447 = {_0, _15445} + {_0, _0, _15446};
  wire _15448 = _12301 < _15447;
  wire _15449 = r1698 ^ _15448;
  wire _15450 = _12298 ? coded_block[1698] : r1698;
  wire _15451 = _12296 ? _15449 : _15450;
  always @ (posedge reset or posedge clock) if (reset) r1698 <= 1'd0; else if (_12300) r1698 <= _15451;
  wire [1:0] _15452 = {_0, _639} + {_0, _2974};
  wire [1:0] _15453 = {_0, _5694} + {_0, _7326};
  wire [2:0] _15454 = {_0, _15452} + {_0, _15453};
  wire [1:0] _15455 = {_0, _9085} + {_0, _12092};
  wire [3:0] _15456 = {_0, _15454} + {_0, _0, _15455};
  wire _15457 = _12301 < _15456;
  wire _15458 = r1697 ^ _15457;
  wire _15459 = _12298 ? coded_block[1697] : r1697;
  wire _15460 = _12296 ? _15458 : _15459;
  always @ (posedge reset or posedge clock) if (reset) r1697 <= 1'd0; else if (_12300) r1697 <= _15460;
  wire [1:0] _15461 = {_0, _672} + {_0, _3901};
  wire [1:0] _15462 = {_0, _5053} + {_0, _7773};
  wire [2:0] _15463 = {_0, _15461} + {_0, _15462};
  wire [1:0] _15464 = {_0, _9406} + {_0, _11165};
  wire [3:0] _15465 = {_0, _15463} + {_0, _0, _15464};
  wire _15466 = _12301 < _15465;
  wire _15467 = r1696 ^ _15466;
  wire _15468 = _12298 ? coded_block[1696] : r1696;
  wire _15469 = _12296 ? _15467 : _15468;
  always @ (posedge reset or posedge clock) if (reset) r1696 <= 1'd0; else if (_12300) r1696 <= _15469;
  wire [1:0] _15470 = {_0, _800} + {_0, _2592};
  wire [1:0] _15471 = {_0, _5790} + {_0, _7612};
  wire [2:0] _15472 = {_0, _15470} + {_0, _15471};
  wire [1:0] _15473 = {_0, _10235} + {_0, _12219};
  wire [3:0] _15474 = {_0, _15472} + {_0, _0, _15473};
  wire _15475 = _12301 < _15474;
  wire _15476 = r1695 ^ _15475;
  wire _15477 = _12298 ? coded_block[1695] : r1695;
  wire _15478 = _12296 ? _15476 : _15477;
  always @ (posedge reset or posedge clock) if (reset) r1695 <= 1'd0; else if (_12300) r1695 <= _15478;
  wire [1:0] _15479 = {_0, _863} + {_0, _2463};
  wire [1:0] _15480 = {_0, _4319} + {_0, _6750};
  wire [2:0] _15481 = {_0, _15479} + {_0, _15480};
  wire [1:0] _15482 = {_0, _9949} + {_0, _11771};
  wire [3:0] _15483 = {_0, _15481} + {_0, _0, _15482};
  wire _15484 = _12301 < _15483;
  wire _15485 = r1694 ^ _15484;
  wire _15486 = _12298 ? coded_block[1694] : r1694;
  wire _15487 = _12296 ? _15485 : _15486;
  always @ (posedge reset or posedge clock) if (reset) r1694 <= 1'd0; else if (_12300) r1694 <= _15487;
  wire [1:0] _15488 = {_0, _927} + {_0, _2686};
  wire [1:0] _15489 = {_0, _4415} + {_0, _6621};
  wire [2:0] _15490 = {_0, _15488} + {_0, _15489};
  wire [1:0] _15491 = {_0, _8480} + {_0, _10910};
  wire [3:0] _15492 = {_0, _15490} + {_0, _0, _15491};
  wire _15493 = _12301 < _15492;
  wire _15494 = r1693 ^ _15493;
  wire _15495 = _12298 ? coded_block[1693] : r1693;
  wire _15496 = _12296 ? _15494 : _15495;
  always @ (posedge reset or posedge clock) if (reset) r1693 <= 1'd0; else if (_12300) r1693 <= _15496;
  wire [1:0] _15497 = {_0, _990} + {_0, _4028};
  wire [1:0] _15498 = {_0, _5501} + {_0, _6845};
  wire [2:0] _15499 = {_0, _15497} + {_0, _15498};
  wire [1:0] _15500 = {_0, _8574} + {_0, _10783};
  wire [3:0] _15501 = {_0, _15499} + {_0, _0, _15500};
  wire _15502 = _12301 < _15501;
  wire _15503 = r1692 ^ _15502;
  wire _15504 = _12298 ? coded_block[1692] : r1692;
  wire _15505 = _12296 ? _15503 : _15504;
  always @ (posedge reset or posedge clock) if (reset) r1692 <= 1'd0; else if (_12300) r1692 <= _15505;
  wire [1:0] _15506 = {_0, _1057} + {_0, _3198};
  wire [1:0] _15507 = {_0, _5663} + {_0, _8186};
  wire [2:0] _15508 = {_0, _15506} + {_0, _15507};
  wire [1:0] _15509 = {_0, _9661} + {_0, _11004};
  wire [3:0] _15510 = {_0, _15508} + {_0, _0, _15509};
  wire _15511 = _12301 < _15510;
  wire _15512 = r1691 ^ _15511;
  wire _15513 = _12298 ? coded_block[1691] : r1691;
  wire _15514 = _12296 ? _15512 : _15513;
  always @ (posedge reset or posedge clock) if (reset) r1691 <= 1'd0; else if (_12300) r1691 <= _15514;
  wire [1:0] _15515 = {_0, _1088} + {_0, _2208};
  wire [1:0] _15516 = {_0, _5279} + {_0, _7741};
  wire [2:0] _15517 = {_0, _15515} + {_0, _15516};
  wire [1:0] _15518 = {_0, _8256} + {_0, _11740};
  wire [3:0] _15519 = {_0, _15517} + {_0, _0, _15518};
  wire _15520 = _12301 < _15519;
  wire _15521 = r1690 ^ _15520;
  wire _15522 = _12298 ? coded_block[1690] : r1690;
  wire _15523 = _12296 ? _15521 : _15522;
  always @ (posedge reset or posedge clock) if (reset) r1690 <= 1'd0; else if (_12300) r1690 <= _15523;
  wire [1:0] _15524 = {_0, _1151} + {_0, _3104};
  wire [1:0] _15525 = {_0, _4703} + {_0, _6366};
  wire [2:0] _15526 = {_0, _15524} + {_0, _15525};
  wire [1:0] _15527 = {_0, _9438} + {_0, _11900};
  wire [3:0] _15528 = {_0, _15526} + {_0, _0, _15527};
  wire _15529 = _12301 < _15528;
  wire _15530 = r1689 ^ _15529;
  wire _15531 = _12298 ? coded_block[1689] : r1689;
  wire _15532 = _12296 ? _15530 : _15531;
  always @ (posedge reset or posedge clock) if (reset) r1689 <= 1'd0; else if (_12300) r1689 <= _15532;
  wire [1:0] _15533 = {_0, _1215} + {_0, _3836};
  wire [1:0] _15534 = {_0, _4605} + {_0, _7262};
  wire [2:0] _15535 = {_0, _15533} + {_0, _15534};
  wire [1:0] _15536 = {_0, _8863} + {_0, _10527};
  wire [3:0] _15537 = {_0, _15535} + {_0, _0, _15536};
  wire _15538 = _12301 < _15537;
  wire _15539 = r1688 ^ _15538;
  wire _15540 = _12298 ? coded_block[1688] : r1688;
  wire _15541 = _12296 ? _15539 : _15540;
  always @ (posedge reset or posedge clock) if (reset) r1688 <= 1'd0; else if (_12300) r1688 <= _15541;
  wire [1:0] _15542 = {_0, _34} + {_0, _2974};
  wire [1:0] _15543 = {_0, _5053} + {_0, _7132};
  wire [2:0] _15544 = {_0, _15542} + {_0, _15543};
  wire [1:0] _15545 = {_0, _9212} + {_0, _11295};
  wire [3:0] _15546 = {_0, _15544} + {_0, _0, _15545};
  wire _15547 = _12301 < _15546;
  wire _15548 = r1687 ^ _15547;
  wire _15549 = _12298 ? coded_block[1687] : r1687;
  wire _15550 = _12296 ? _15548 : _15549;
  always @ (posedge reset or posedge clock) if (reset) r1687 <= 1'd0; else if (_12300) r1687 <= _15550;
  wire [1:0] _15551 = {_0, _1854} + {_0, _2878};
  wire [1:0] _15552 = {_0, _4350} + {_0, _7710};
  wire [2:0] _15553 = {_0, _15551} + {_0, _15552};
  wire [1:0] _15554 = {_0, _9438} + {_0, _11644};
  wire [3:0] _15555 = {_0, _15553} + {_0, _0, _15554};
  wire _15556 = _12301 < _15555;
  wire _15557 = r1686 ^ _15556;
  wire _15558 = _12298 ? coded_block[1686] : r1686;
  wire _15559 = _12296 ? _15557 : _15558;
  always @ (posedge reset or posedge clock) if (reset) r1686 <= 1'd0; else if (_12300) r1686 <= _15559;
  wire [1:0] _15560 = {_0, _1886} + {_0, _2430};
  wire [1:0] _15561 = {_0, _4958} + {_0, _6431};
  wire [2:0] _15562 = {_0, _15560} + {_0, _15561};
  wire [1:0] _15563 = {_0, _9790} + {_0, _11516};
  wire [3:0] _15564 = {_0, _15562} + {_0, _0, _15563};
  wire _15565 = _12301 < _15564;
  wire _15566 = r1685 ^ _15565;
  wire _15567 = _12298 ? coded_block[1685] : r1685;
  wire _15568 = _12296 ? _15566 : _15567;
  always @ (posedge reset or posedge clock) if (reset) r1685 <= 1'd0; else if (_12300) r1685 <= _15568;
  wire [1:0] _15569 = {_0, _1950} + {_0, _3068};
  wire [1:0] _15570 = {_0, _6139} + {_0, _6589};
  wire [2:0] _15571 = {_0, _15569} + {_0, _15570};
  wire [1:0] _15572 = {_0, _9118} + {_0, _10590};
  wire [3:0] _15573 = {_0, _15571} + {_0, _0, _15572};
  wire _15574 = _12301 < _15573;
  wire _15575 = r1684 ^ _15574;
  wire _15576 = _12298 ? coded_block[1684] : r1684;
  wire _15577 = _12296 ? _15575 : _15576;
  always @ (posedge reset or posedge clock) if (reset) r1684 <= 1'd0; else if (_12300) r1684 <= _15577;
  wire [1:0] _15578 = {_0, _1981} + {_0, _3486};
  wire [1:0] _15579 = {_0, _5152} + {_0, _6207};
  wire [2:0] _15580 = {_0, _15578} + {_0, _15579};
  wire [1:0] _15581 = {_0, _8670} + {_0, _11196};
  wire [3:0] _15582 = {_0, _15580} + {_0, _0, _15581};
  wire _15583 = _12301 < _15582;
  wire _15584 = r1683 ^ _15583;
  wire _15585 = _12298 ? coded_block[1683] : r1683;
  wire _15586 = _12296 ? _15584 : _15585;
  always @ (posedge reset or posedge clock) if (reset) r1683 <= 1'd0; else if (_12300) r1683 <= _15586;
  wire [1:0] _15587 = {_0, _2013} + {_0, _3964};
  wire [1:0] _15588 = {_0, _5565} + {_0, _7230};
  wire [2:0] _15589 = {_0, _15587} + {_0, _15588};
  wire [1:0] _15590 = {_0, _8288} + {_0, _10748};
  wire [3:0] _15591 = {_0, _15589} + {_0, _0, _15590};
  wire _15592 = _12301 < _15591;
  wire _15593 = r1682 ^ _15592;
  wire _15594 = _12298 ? coded_block[1682] : r1682;
  wire _15595 = _12296 ? _15593 : _15594;
  always @ (posedge reset or posedge clock) if (reset) r1682 <= 1'd0; else if (_12300) r1682 <= _15595;
  wire [1:0] _15596 = {_0, _65} + {_0, _2686};
  wire [1:0] _15597 = {_0, _5470} + {_0, _8123};
  wire [2:0] _15598 = {_0, _15596} + {_0, _15597};
  wire [1:0] _15599 = {_0, _9724} + {_0, _11389};
  wire [3:0] _15600 = {_0, _15598} + {_0, _0, _15599};
  wire _15601 = _12301 < _15600;
  wire _15602 = r1681 ^ _15601;
  wire _15603 = _12298 ? coded_block[1681] : r1681;
  wire _15604 = _12296 ? _15602 : _15603;
  always @ (posedge reset or posedge clock) if (reset) r1681 <= 1'd0; else if (_12300) r1681 <= _15604;
  wire [1:0] _15605 = {_0, _128} + {_0, _2526};
  wire [1:0] _15606 = {_0, _4447} + {_0, _6845};
  wire [2:0] _15607 = {_0, _15605} + {_0, _15606};
  wire [1:0] _15608 = {_0, _9630} + {_0, _12282};
  wire [3:0] _15609 = {_0, _15607} + {_0, _0, _15608};
  wire _15610 = _12301 < _15609;
  wire _15611 = r1680 ^ _15610;
  wire _15612 = _12298 ? coded_block[1680] : r1680;
  wire _15613 = _12296 ? _15611 : _15612;
  always @ (posedge reset or posedge clock) if (reset) r1680 <= 1'd0; else if (_12300) r1680 <= _15613;
  wire [1:0] _15614 = {_0, _161} + {_0, _2336};
  wire [1:0] _15615 = {_0, _4605} + {_0, _6525};
  wire [2:0] _15616 = {_0, _15614} + {_0, _15615};
  wire [1:0] _15617 = {_0, _8926} + {_0, _11708};
  wire [3:0] _15618 = {_0, _15616} + {_0, _0, _15617};
  wire _15619 = _12301 < _15618;
  wire _15620 = r1679 ^ _15619;
  wire _15621 = _12298 ? coded_block[1679] : r1679;
  wire _15622 = _12296 ? _15620 : _15621;
  always @ (posedge reset or posedge clock) if (reset) r1679 <= 1'd0; else if (_12300) r1679 <= _15622;
  wire [1:0] _15623 = {_0, _192} + {_0, _2719};
  wire [1:0] _15624 = {_0, _4415} + {_0, _6687};
  wire [2:0] _15625 = {_0, _15623} + {_0, _15624};
  wire [1:0] _15626 = {_0, _8607} + {_0, _11004};
  wire [3:0] _15627 = {_0, _15625} + {_0, _0, _15626};
  wire _15628 = _12301 < _15627;
  wire _15629 = r1678 ^ _15628;
  wire _15630 = _12298 ? coded_block[1678] : r1678;
  wire _15631 = _12296 ? _15629 : _15630;
  always @ (posedge reset or posedge clock) if (reset) r1678 <= 1'd0; else if (_12300) r1678 <= _15631;
  wire [1:0] _15632 = {_0, _255} + {_0, _3646};
  wire [1:0] _15633 = {_0, _5949} + {_0, _6877};
  wire [2:0] _15634 = {_0, _15632} + {_0, _15633};
  wire [1:0] _15635 = {_0, _8574} + {_0, _10846};
  wire [3:0] _15636 = {_0, _15634} + {_0, _0, _15635};
  wire _15637 = _12301 < _15636;
  wire _15638 = r1677 ^ _15637;
  wire _15639 = _12298 ? coded_block[1677] : r1677;
  wire _15640 = _12296 ? _15638 : _15639;
  always @ (posedge reset or posedge clock) if (reset) r1677 <= 1'd0; else if (_12300) r1677 <= _15640;
  wire [1:0] _15641 = {_0, _289} + {_0, _2208};
  wire [1:0] _15642 = {_0, _5726} + {_0, _8028};
  wire [2:0] _15643 = {_0, _15641} + {_0, _15642};
  wire [1:0] _15644 = {_0, _8957} + {_0, _10654};
  wire [3:0] _15645 = {_0, _15643} + {_0, _0, _15644};
  wire _15646 = _12301 < _15645;
  wire _15647 = r1676 ^ _15646;
  wire _15648 = _12298 ? coded_block[1676] : r1676;
  wire _15649 = _12296 ? _15647 : _15648;
  always @ (posedge reset or posedge clock) if (reset) r1676 <= 1'd0; else if (_12300) r1676 <= _15649;
  wire [1:0] _15650 = {_0, _320} + {_0, _2144};
  wire [1:0] _15651 = {_0, _4287} + {_0, _7804};
  wire [2:0] _15652 = {_0, _15650} + {_0, _15651};
  wire [1:0] _15653 = {_0, _10108} + {_0, _11038};
  wire [3:0] _15654 = {_0, _15652} + {_0, _0, _15653};
  wire _15655 = _12301 < _15654;
  wire _15656 = r1675 ^ _15655;
  wire _15657 = _12298 ? coded_block[1675] : r1675;
  wire _15658 = _12296 ? _15656 : _15657;
  always @ (posedge reset or posedge clock) if (reset) r1675 <= 1'd0; else if (_12300) r1675 <= _15658;
  wire [1:0] _15659 = {_0, _352} + {_0, _3262};
  wire [1:0] _15660 = {_0, _4223} + {_0, _6366};
  wire [2:0] _15661 = {_0, _15659} + {_0, _15660};
  wire [1:0] _15662 = {_0, _9886} + {_0, _12188};
  wire [3:0] _15663 = {_0, _15661} + {_0, _0, _15662};
  wire _15664 = _12301 < _15663;
  wire _15665 = r1674 ^ _15664;
  wire _15666 = _12298 ? coded_block[1674] : r1674;
  wire _15667 = _12296 ? _15665 : _15666;
  always @ (posedge reset or posedge clock) if (reset) r1674 <= 1'd0; else if (_12300) r1674 <= _15667;
  wire [1:0] _15668 = {_0, _383} + {_0, _3933};
  wire [1:0] _15669 = {_0, _5342} + {_0, _6303};
  wire [2:0] _15670 = {_0, _15668} + {_0, _15669};
  wire [1:0] _15671 = {_0, _8446} + {_0, _11964};
  wire [3:0] _15672 = {_0, _15670} + {_0, _0, _15671};
  wire _15673 = _12301 < _15672;
  wire _15674 = r1673 ^ _15673;
  wire _15675 = _12298 ? coded_block[1673] : r1673;
  wire _15676 = _12296 ? _15674 : _15675;
  always @ (posedge reset or posedge clock) if (reset) r1673 <= 1'd0; else if (_12300) r1673 <= _15676;
  wire [1:0] _15677 = {_0, _416} + {_0, _3517};
  wire [1:0] _15678 = {_0, _6012} + {_0, _7420};
  wire [2:0] _15679 = {_0, _15677} + {_0, _15678};
  wire [1:0] _15680 = {_0, _8383} + {_0, _10527};
  wire [3:0] _15681 = {_0, _15679} + {_0, _0, _15680};
  wire _15682 = _12301 < _15681;
  wire _15683 = r1672 ^ _15682;
  wire _15684 = _12298 ? coded_block[1672] : r1672;
  wire _15685 = _12296 ? _15683 : _15684;
  always @ (posedge reset or posedge clock) if (reset) r1672 <= 1'd0; else if (_12300) r1672 <= _15685;
  wire [1:0] _15686 = {_0, _447} + {_0, _3231};
  wire [1:0] _15687 = {_0, _5597} + {_0, _8092};
  wire [2:0] _15688 = {_0, _15686} + {_0, _15687};
  wire [1:0] _15689 = {_0, _9503} + {_0, _10462};
  wire [3:0] _15690 = {_0, _15688} + {_0, _0, _15689};
  wire _15691 = _12301 < _15690;
  wire _15692 = r1671 ^ _15691;
  wire _15693 = _12298 ? coded_block[1671] : r1671;
  wire _15694 = _12296 ? _15692 : _15693;
  always @ (posedge reset or posedge clock) if (reset) r1671 <= 1'd0; else if (_12300) r1671 <= _15694;
  wire [1:0] _15695 = {_0, _545} + {_0, _2655};
  wire [1:0] _15696 = {_0, _5757} + {_0, _6334};
  wire [2:0] _15697 = {_0, _15695} + {_0, _15696};
  wire [1:0] _15698 = {_0, _9469} + {_0, _11837};
  wire [3:0] _15699 = {_0, _15697} + {_0, _0, _15698};
  wire _15700 = _12301 < _15699;
  wire _15701 = r1670 ^ _15700;
  wire _15702 = _12298 ? coded_block[1670] : r1670;
  wire _15703 = _12296 ? _15701 : _15702;
  always @ (posedge reset or posedge clock) if (reset) r1670 <= 1'd0; else if (_12300) r1670 <= _15703;
  wire [1:0] _15704 = {_0, _639} + {_0, _2112};
  wire [1:0] _15705 = {_0, _4671} + {_0, _7581};
  wire [2:0] _15706 = {_0, _15704} + {_0, _15705};
  wire [1:0] _15707 = {_0, _8894} + {_0, _11996};
  wire [3:0] _15708 = {_0, _15706} + {_0, _0, _15707};
  wire _15709 = _12301 < _15708;
  wire _15710 = r1669 ^ _15709;
  wire _15711 = _12298 ? coded_block[1669] : r1669;
  wire _15712 = _12296 ? _15710 : _15711;
  always @ (posedge reset or posedge clock) if (reset) r1669 <= 1'd0; else if (_12300) r1669 <= _15712;
  wire [1:0] _15713 = {_0, _703} + {_0, _3580};
  wire [1:0] _15714 = {_0, _4319} + {_0, _6270};
  wire [2:0] _15715 = {_0, _15713} + {_0, _15714};
  wire [1:0] _15716 = {_0, _8830} + {_0, _11740};
  wire [3:0] _15717 = {_0, _15715} + {_0, _0, _15716};
  wire _15718 = _12301 < _15717;
  wire _15719 = r1668 ^ _15718;
  wire _15720 = _12298 ? coded_block[1668] : r1668;
  wire _15721 = _12296 ? _15719 : _15720;
  always @ (posedge reset or posedge clock) if (reset) r1668 <= 1'd0; else if (_12300) r1668 <= _15721;
  wire [1:0] _15722 = {_0, _800} + {_0, _3615};
  wire [1:0] _15723 = {_0, _4861} + {_0, _6973};
  wire [2:0] _15724 = {_0, _15722} + {_0, _15723};
  wire [1:0] _15725 = {_0, _9822} + {_0, _10558};
  wire [3:0] _15726 = {_0, _15724} + {_0, _0, _15725};
  wire _15727 = _12301 < _15726;
  wire _15728 = r1667 ^ _15727;
  wire _15729 = _12298 ? coded_block[1667] : r1667;
  wire _15730 = _12296 ? _15728 : _15729;
  always @ (posedge reset or posedge clock) if (reset) r1667 <= 1'd0; else if (_12300) r1667 <= _15730;
  wire [1:0] _15731 = {_0, _863} + {_0, _3294};
  wire [1:0] _15732 = {_0, _5981} + {_0, _7773};
  wire [2:0] _15733 = {_0, _15731} + {_0, _15732};
  wire [1:0] _15734 = {_0, _9022} + {_0, _11132};
  wire [3:0] _15735 = {_0, _15733} + {_0, _0, _15734};
  wire _15736 = _12301 < _15735;
  wire _15737 = r1666 ^ _15736;
  wire _15738 = _12298 ? coded_block[1666] : r1666;
  wire _15739 = _12296 ? _15737 : _15738;
  always @ (posedge reset or posedge clock) if (reset) r1666 <= 1'd0; else if (_12300) r1666 <= _15739;
  wire [1:0] _15740 = {_0, _894} + {_0, _3135};
  wire [1:0] _15741 = {_0, _5373} + {_0, _8059};
  wire [2:0] _15742 = {_0, _15740} + {_0, _15741};
  wire [1:0] _15743 = {_0, _9853} + {_0, _11101};
  wire [3:0] _15744 = {_0, _15742} + {_0, _0, _15743};
  wire _15745 = _12301 < _15744;
  wire _15746 = r1665 ^ _15745;
  wire _15747 = _12298 ? coded_block[1665] : r1665;
  wire _15748 = _12296 ? _15746 : _15747;
  always @ (posedge reset or posedge clock) if (reset) r1665 <= 1'd0; else if (_12300) r1665 <= _15748;
  wire [1:0] _15749 = {_0, _927} + {_0, _2081};
  wire [1:0] _15750 = {_0, _5215} + {_0, _7454};
  wire [2:0] _15751 = {_0, _15749} + {_0, _15750};
  wire [1:0] _15752 = {_0, _10141} + {_0, _11933};
  wire [3:0] _15753 = {_0, _15751} + {_0, _0, _15752};
  wire _15754 = _12301 < _15753;
  wire _15755 = r1664 ^ _15754;
  wire _15756 = _12298 ? coded_block[1664] : r1664;
  wire _15757 = _12296 ? _15755 : _15756;
  always @ (posedge reset or posedge clock) if (reset) r1664 <= 1'd0; else if (_12300) r1664 <= _15757;
  wire [1:0] _15758 = {_0, _990} + {_0, _3359};
  wire [1:0] _15759 = {_0, _5246} + {_0, _6176};
  wire [2:0] _15760 = {_0, _15758} + {_0, _15759};
  wire [1:0] _15761 = {_0, _9375} + {_0, _11613};
  wire [3:0] _15762 = {_0, _15760} + {_0, _0, _15761};
  wire _15763 = _12301 < _15762;
  wire _15764 = r1663 ^ _15763;
  wire _15765 = _12298 ? coded_block[1663] : r1663;
  wire _15766 = _12296 ? _15764 : _15765;
  always @ (posedge reset or posedge clock) if (reset) r1663 <= 1'd0; else if (_12300) r1663 <= _15766;
  wire [1:0] _15767 = {_0, _1057} + {_0, _3742};
  wire [1:0] _15768 = {_0, _6076} + {_0, _7517};
  wire [2:0] _15769 = {_0, _15767} + {_0, _15768};
  wire [1:0] _15770 = {_0, _9406} + {_0, _10272};
  wire [3:0] _15771 = {_0, _15769} + {_0, _0, _15770};
  wire _15772 = _12301 < _15771;
  wire _15773 = r1662 ^ _15772;
  wire _15774 = _12298 ? coded_block[1662] : r1662;
  wire _15775 = _12296 ? _15773 : _15774;
  always @ (posedge reset or posedge clock) if (reset) r1662 <= 1'd0; else if (_12300) r1662 <= _15775;
  wire [1:0] _15776 = {_0, _1120} + {_0, _3005};
  wire [1:0] _15777 = {_0, _5022} + {_0, _7900};
  wire [2:0] _15778 = {_0, _15776} + {_0, _15777};
  wire [1:0] _15779 = {_0, _10235} + {_0, _11677};
  wire [3:0] _15780 = {_0, _15778} + {_0, _0, _15779};
  wire _15781 = _12301 < _15780;
  wire _15782 = r1661 ^ _15781;
  wire _15783 = _12298 ? coded_block[1661] : r1661;
  wire _15784 = _12296 ? _15782 : _15783;
  always @ (posedge reset or posedge clock) if (reset) r1661 <= 1'd0; else if (_12300) r1661 <= _15784;
  wire [1:0] _15785 = {_0, _1151} + {_0, _3805};
  wire [1:0] _15786 = {_0, _5085} + {_0, _7100};
  wire [2:0] _15787 = {_0, _15785} + {_0, _15786};
  wire [1:0] _15788 = {_0, _9980} + {_0, _10303};
  wire [3:0] _15789 = {_0, _15787} + {_0, _0, _15788};
  wire _15790 = _12301 < _15789;
  wire _15791 = r1660 ^ _15790;
  wire _15792 = _12298 ? coded_block[1660] : r1660;
  wire _15793 = _12296 ? _15791 : _15792;
  always @ (posedge reset or posedge clock) if (reset) r1660 <= 1'd0; else if (_12300) r1660 <= _15793;
  wire [1:0] _15794 = {_0, _1184} + {_0, _2494};
  wire [1:0] _15795 = {_0, _5884} + {_0, _7163};
  wire [2:0] _15796 = {_0, _15794} + {_0, _15795};
  wire [1:0] _15797 = {_0, _9181} + {_0, _12061};
  wire [3:0] _15798 = {_0, _15796} + {_0, _0, _15797};
  wire _15799 = _12301 < _15798;
  wire _15800 = r1659 ^ _15799;
  wire _15801 = _12298 ? coded_block[1659] : r1659;
  wire _15802 = _12296 ? _15800 : _15801;
  always @ (posedge reset or posedge clock) if (reset) r1659 <= 1'd0; else if (_12300) r1659 <= _15802;
  wire [1:0] _15803 = {_0, _1215} + {_0, _2399};
  wire [1:0] _15804 = {_0, _4574} + {_0, _7965};
  wire [2:0] _15805 = {_0, _15803} + {_0, _15804};
  wire [1:0] _15806 = {_0, _9248} + {_0, _11259};
  wire [3:0] _15807 = {_0, _15805} + {_0, _0, _15806};
  wire _15808 = _12301 < _15807;
  wire _15809 = r1658 ^ _15808;
  wire _15810 = _12298 ? coded_block[1658] : r1658;
  wire _15811 = _12296 ? _15809 : _15810;
  always @ (posedge reset or posedge clock) if (reset) r1658 <= 1'd0; else if (_12300) r1658 <= _15811;
  wire [1:0] _15812 = {_0, _1278} + {_0, _3773};
  wire [1:0] _15813 = {_0, _4989} + {_0, _6558};
  wire [2:0] _15814 = {_0, _15812} + {_0, _15813};
  wire [1:0] _15815 = {_0, _8736} + {_0, _12124};
  wire [3:0] _15816 = {_0, _15814} + {_0, _0, _15815};
  wire _15817 = _12301 < _15816;
  wire _15818 = r1657 ^ _15817;
  wire _15819 = _12298 ? coded_block[1657] : r1657;
  wire _15820 = _12296 ? _15818 : _15819;
  always @ (posedge reset or posedge clock) if (reset) r1657 <= 1'd0; else if (_12300) r1657 <= _15820;
  wire [1:0] _15821 = {_0, _1312} + {_0, _3037};
  wire [1:0] _15822 = {_0, _5853} + {_0, _7069};
  wire [2:0] _15823 = {_0, _15821} + {_0, _15822};
  wire [1:0] _15824 = {_0, _8638} + {_0, _10814};
  wire [3:0] _15825 = {_0, _15823} + {_0, _0, _15824};
  wire _15826 = _12301 < _15825;
  wire _15827 = r1656 ^ _15826;
  wire _15828 = _12298 ? coded_block[1656] : r1656;
  wire _15829 = _12296 ? _15827 : _15828;
  always @ (posedge reset or posedge clock) if (reset) r1656 <= 1'd0; else if (_12300) r1656 <= _15829;
  wire [1:0] _15830 = {_0, _1375} + {_0, _2623};
  wire [1:0] _15831 = {_0, _4160} + {_0, _7199};
  wire [2:0] _15832 = {_0, _15830} + {_0, _15831};
  wire [1:0] _15833 = {_0, _10014} + {_0, _11228};
  wire [3:0] _15834 = {_0, _15832} + {_0, _0, _15833};
  wire _15835 = _12301 < _15834;
  wire _15836 = r1655 ^ _15835;
  wire _15837 = _12298 ? coded_block[1655] : r1655;
  wire _15838 = _12296 ? _15836 : _15837;
  always @ (posedge reset or posedge clock) if (reset) r1655 <= 1'd0; else if (_12300) r1655 <= _15838;
  wire [1:0] _15839 = {_0, _1406} + {_0, _3709};
  wire [1:0] _15840 = {_0, _4703} + {_0, _6239};
  wire [2:0] _15841 = {_0, _15839} + {_0, _15840};
  wire [1:0] _15842 = {_0, _9279} + {_0, _12092};
  wire [3:0] _15843 = {_0, _15841} + {_0, _0, _15842};
  wire _15844 = _12301 < _15843;
  wire _15845 = r1654 ^ _15844;
  wire _15846 = _12298 ? coded_block[1654] : r1654;
  wire _15847 = _12296 ? _15845 : _15846;
  always @ (posedge reset or posedge clock) if (reset) r1654 <= 1'd0; else if (_12300) r1654 <= _15847;
  wire [1:0] _15848 = {_0, _1470} + {_0, _2463};
  wire [1:0] _15849 = {_0, _6108} + {_0, _7868};
  wire [2:0] _15850 = {_0, _15848} + {_0, _15849};
  wire [1:0] _15851 = {_0, _8863} + {_0, _10399};
  wire [3:0] _15852 = {_0, _15850} + {_0, _0, _15851};
  wire _15853 = _12301 < _15852;
  wire _15854 = r1653 ^ _15853;
  wire _15855 = _12298 ? coded_block[1653] : r1653;
  wire _15856 = _12296 ? _15854 : _15855;
  always @ (posedge reset or posedge clock) if (reset) r1653 <= 1'd0; else if (_12300) r1653 <= _15856;
  wire [1:0] _15857 = {_0, _1533} + {_0, _2750};
  wire [1:0] _15858 = {_0, _5918} + {_0, _6621};
  wire [2:0] _15859 = {_0, _15857} + {_0, _15858};
  wire [1:0] _15860 = {_0, _8256} + {_0, _12027};
  wire [3:0] _15861 = {_0, _15859} + {_0, _0, _15860};
  wire _15862 = _12301 < _15861;
  wire _15863 = r1652 ^ _15862;
  wire _15864 = _12298 ? coded_block[1652] : r1652;
  wire _15865 = _12296 ? _15863 : _15864;
  always @ (posedge reset or posedge clock) if (reset) r1652 <= 1'd0; else if (_12300) r1652 <= _15865;
  wire [1:0] _15866 = {_0, _1599} + {_0, _2302};
  wire [1:0] _15867 = {_0, _4926} + {_0, _6908};
  wire [2:0] _15868 = {_0, _15866} + {_0, _15867};
  wire [1:0] _15869 = {_0, _10077} + {_0, _10783};
  wire [3:0] _15870 = {_0, _15868} + {_0, _0, _15869};
  wire _15871 = _12301 < _15870;
  wire _15872 = r1651 ^ _15871;
  wire _15873 = _12298 ? coded_block[1651] : r1651;
  wire _15874 = _12296 ? _15872 : _15873;
  always @ (posedge reset or posedge clock) if (reset) r1651 <= 1'd0; else if (_12300) r1651 <= _15874;
  wire [1:0] _15875 = {_0, _1726} + {_0, _3325};
  wire [1:0] _15876 = {_0, _5183} + {_0, _7612};
  wire [2:0] _15877 = {_0, _15875} + {_0, _15876};
  wire [1:0] _15878 = {_0, _8799} + {_0, _10621};
  wire [3:0] _15879 = {_0, _15877} + {_0, _0, _15878};
  wire _15880 = _12301 < _15879;
  wire _15881 = r1650 ^ _15880;
  wire _15882 = _12298 ? coded_block[1650] : r1650;
  wire _15883 = _12296 ? _15881 : _15882;
  always @ (posedge reset or posedge clock) if (reset) r1650 <= 1'd0; else if (_12300) r1650 <= _15883;
  wire [1:0] _15884 = {_0, _1758} + {_0, _3198};
  wire [1:0] _15885 = {_0, _5407} + {_0, _7262};
  wire [2:0] _15886 = {_0, _15884} + {_0, _15885};
  wire [1:0] _15887 = {_0, _9693} + {_0, _10877};
  wire [3:0] _15888 = {_0, _15886} + {_0, _0, _15887};
  wire _15889 = _12301 < _15888;
  wire _15890 = r1649 ^ _15889;
  wire _15891 = _12298 ? coded_block[1649] : r1649;
  wire _15892 = _12296 ? _15890 : _15891;
  always @ (posedge reset or posedge clock) if (reset) r1649 <= 1'd0; else if (_12300) r1649 <= _15892;
  wire [1:0] _15893 = {_0, _34} + {_0, _3836};
  wire [1:0] _15894 = {_0, _5918} + {_0, _7996};
  wire [2:0] _15895 = {_0, _15893} + {_0, _15894};
  wire [1:0] _15896 = {_0, _10077} + {_0, _12155};
  wire [3:0] _15897 = {_0, _15895} + {_0, _0, _15896};
  wire _15898 = _12301 < _15897;
  wire _15899 = r1648 ^ _15898;
  wire _15900 = _12298 ? coded_block[1648] : r1648;
  wire _15901 = _12296 ? _15899 : _15900;
  always @ (posedge reset or posedge clock) if (reset) r1648 <= 1'd0; else if (_12300) r1648 <= _15901;
  wire [1:0] _15902 = {_0, _128} + {_0, _2623};
  wire [1:0] _15903 = {_0, _5853} + {_0, _7420};
  wire [2:0] _15904 = {_0, _15902} + {_0, _15903};
  wire [1:0] _15905 = {_0, _9597} + {_0, _10973};
  wire [3:0] _15906 = {_0, _15904} + {_0, _0, _15905};
  wire _15907 = _12301 < _15906;
  wire _15908 = r1647 ^ _15907;
  wire _15909 = _12298 ? coded_block[1647] : r1647;
  wire _15910 = _12296 ? _15908 : _15909;
  always @ (posedge reset or posedge clock) if (reset) r1647 <= 1'd0; else if (_12300) r1647 <= _15910;
  wire [1:0] _15911 = {_0, _161} + {_0, _3901};
  wire [1:0] _15912 = {_0, _4703} + {_0, _7931};
  wire [2:0] _15913 = {_0, _15911} + {_0, _15912};
  wire [1:0] _15914 = {_0, _9503} + {_0, _11677};
  wire [3:0] _15915 = {_0, _15913} + {_0, _0, _15914};
  wire _15916 = _12301 < _15915;
  wire _15917 = r1646 ^ _15916;
  wire _15918 = _12298 ? coded_block[1646] : r1646;
  wire _15919 = _12296 ? _15917 : _15918;
  always @ (posedge reset or posedge clock) if (reset) r1646 <= 1'd0; else if (_12300) r1646 <= _15919;
  wire [1:0] _15920 = {_0, _192} + {_0, _2941};
  wire [1:0] _15921 = {_0, _5981} + {_0, _6781};
  wire [2:0] _15922 = {_0, _15920} + {_0, _15921};
  wire [1:0] _15923 = {_0, _10014} + {_0, _11581};
  wire [3:0] _15924 = {_0, _15922} + {_0, _0, _15923};
  wire _15925 = _12301 < _15924;
  wire _15926 = r1645 ^ _15925;
  wire _15927 = _12298 ? coded_block[1645] : r1645;
  wire _15928 = _12296 ? _15926 : _15927;
  always @ (posedge reset or posedge clock) if (reset) r1645 <= 1'd0; else if (_12300) r1645 <= _15928;
  wire [1:0] _15929 = {_0, _224} + {_0, _3486};
  wire [1:0] _15930 = {_0, _5022} + {_0, _8059};
  wire [2:0] _15931 = {_0, _15929} + {_0, _15930};
  wire [1:0] _15932 = {_0, _8863} + {_0, _12092};
  wire [3:0] _15933 = {_0, _15931} + {_0, _0, _15932};
  wire _15934 = _12301 < _15933;
  wire _15935 = r1644 ^ _15934;
  wire _15936 = _12298 ? coded_block[1644] : r1644;
  wire _15937 = _12296 ? _15935 : _15936;
  always @ (posedge reset or posedge clock) if (reset) r1644 <= 1'd0; else if (_12300) r1644 <= _15937;
  wire [1:0] _15938 = {_0, _289} + {_0, _2878};
  wire [1:0] _15939 = {_0, _4640} + {_0, _7644};
  wire [2:0] _15940 = {_0, _15938} + {_0, _15939};
  wire [1:0] _15941 = {_0, _9181} + {_0, _12219};
  wire [3:0] _15942 = {_0, _15940} + {_0, _0, _15941};
  wire _15943 = _12301 < _15942;
  wire _15944 = r1643 ^ _15943;
  wire _15945 = _12298 ? coded_block[1643] : r1643;
  wire _15946 = _12296 ? _15944 : _15945;
  always @ (posedge reset or posedge clock) if (reset) r1643 <= 1'd0; else if (_12300) r1643 <= _15946;
  wire [1:0] _15947 = {_0, _320} + {_0, _3325};
  wire [1:0] _15948 = {_0, _4958} + {_0, _6718};
  wire [2:0] _15949 = {_0, _15947} + {_0, _15948};
  wire [1:0] _15950 = {_0, _9724} + {_0, _11259};
  wire [3:0] _15951 = {_0, _15949} + {_0, _0, _15950};
  wire _15952 = _12301 < _15951;
  wire _15953 = r1642 ^ _15952;
  wire _15954 = _12298 ? coded_block[1642] : r1642;
  wire _15955 = _12296 ? _15953 : _15954;
  always @ (posedge reset or posedge clock) if (reset) r1642 <= 1'd0; else if (_12300) r1642 <= _15955;
  wire [1:0] _15956 = {_0, _352} + {_0, _2686};
  wire [1:0] _15957 = {_0, _5407} + {_0, _7036};
  wire [2:0] _15958 = {_0, _15956} + {_0, _15957};
  wire [1:0] _15959 = {_0, _8799} + {_0, _11806};
  wire [3:0] _15960 = {_0, _15958} + {_0, _0, _15959};
  wire _15961 = _12301 < _15960;
  wire _15962 = r1641 ^ _15961;
  wire _15963 = _12298 ? coded_block[1641] : r1641;
  wire _15964 = _12296 ? _15962 : _15963;
  always @ (posedge reset or posedge clock) if (reset) r1641 <= 1'd0; else if (_12300) r1641 <= _15964;
  wire [1:0] _15965 = {_0, _383} + {_0, _3615};
  wire [1:0] _15966 = {_0, _4767} + {_0, _7485};
  wire [2:0] _15967 = {_0, _15965} + {_0, _15966};
  wire [1:0] _15968 = {_0, _9118} + {_0, _10877};
  wire [3:0] _15969 = {_0, _15967} + {_0, _0, _15968};
  wire _15970 = _12301 < _15969;
  wire _15971 = r1640 ^ _15970;
  wire _15972 = _12298 ? coded_block[1640] : r1640;
  wire _15973 = _12296 ? _15971 : _15972;
  always @ (posedge reset or posedge clock) if (reset) r1640 <= 1'd0; else if (_12300) r1640 <= _15973;
  wire [1:0] _15974 = {_0, _416} + {_0, _3709};
  wire [1:0] _15975 = {_0, _5694} + {_0, _6845};
  wire [2:0] _15976 = {_0, _15974} + {_0, _15975};
  wire [1:0] _15977 = {_0, _9566} + {_0, _11196};
  wire [3:0] _15978 = {_0, _15976} + {_0, _0, _15977};
  wire _15979 = _12301 < _15978;
  wire _15980 = r1639 ^ _15979;
  wire _15981 = _12298 ? coded_block[1639] : r1639;
  wire _15982 = _12296 ? _15980 : _15981;
  always @ (posedge reset or posedge clock) if (reset) r1639 <= 1'd0; else if (_12300) r1639 <= _15982;
  wire [1:0] _15983 = {_0, _447} + {_0, _3167};
  wire [1:0] _15984 = {_0, _5790} + {_0, _7773};
  wire [2:0] _15985 = {_0, _15983} + {_0, _15984};
  wire [1:0] _15986 = {_0, _8926} + {_0, _11644};
  wire [3:0] _15987 = {_0, _15985} + {_0, _0, _15986};
  wire _15988 = _12301 < _15987;
  wire _15989 = r1638 ^ _15988;
  wire _15990 = _12298 ? coded_block[1638] : r1638;
  wire _15991 = _12296 ? _15989 : _15990;
  always @ (posedge reset or posedge clock) if (reset) r1638 <= 1'd0; else if (_12300) r1638 <= _15991;
  wire [1:0] _15992 = {_0, _479} + {_0, _3422};
  wire [1:0] _15993 = {_0, _5246} + {_0, _7868};
  wire [2:0] _15994 = {_0, _15992} + {_0, _15993};
  wire [1:0] _15995 = {_0, _9853} + {_0, _11004};
  wire [3:0] _15996 = {_0, _15994} + {_0, _0, _15995};
  wire _15997 = _12301 < _15996;
  wire _15998 = r1637 ^ _15997;
  wire _15999 = _12298 ? coded_block[1637] : r1637;
  wire _16000 = _12296 ? _15998 : _15999;
  always @ (posedge reset or posedge clock) if (reset) r1637 <= 1'd0; else if (_12300) r1637 <= _16000;
  wire [1:0] _16001 = {_0, _545} + {_0, _3964};
  wire [1:0] _16002 = {_0, _4384} + {_0, _7581};
  wire [2:0] _16003 = {_0, _16001} + {_0, _16002};
  wire [1:0] _16004 = {_0, _9406} + {_0, _12027};
  wire [3:0] _16005 = {_0, _16003} + {_0, _0, _16004};
  wire _16006 = _12301 < _16005;
  wire _16007 = r1636 ^ _16006;
  wire _16008 = _12298 ? coded_block[1636] : r1636;
  wire _16009 = _12296 ? _16007 : _16008;
  always @ (posedge reset or posedge clock) if (reset) r1636 <= 1'd0; else if (_12300) r1636 <= _16009;
  wire [1:0] _16010 = {_0, _608} + {_0, _4060};
  wire [1:0] _16011 = {_0, _4256} + {_0, _8123};
  wire [2:0] _16012 = {_0, _16010} + {_0, _16011};
  wire [1:0] _16013 = {_0, _8543} + {_0, _11740};
  wire [3:0] _16014 = {_0, _16012} + {_0, _0, _16013};
  wire _16015 = _12301 < _16014;
  wire _16016 = r1635 ^ _16015;
  wire _16017 = _12298 ? coded_block[1635] : r1635;
  wire _16018 = _12296 ? _16016 : _16017;
  always @ (posedge reset or posedge clock) if (reset) r1635 <= 1'd0; else if (_12300) r1635 <= _16018;
  wire [1:0] _16019 = {_0, _639} + {_0, _2399};
  wire [1:0] _16020 = {_0, _6139} + {_0, _6334};
  wire [2:0] _16021 = {_0, _16019} + {_0, _16020};
  wire [1:0] _16022 = {_0, _10204} + {_0, _10621};
  wire [3:0] _16023 = {_0, _16021} + {_0, _0, _16022};
  wire _16024 = _12301 < _16023;
  wire _16025 = r1634 ^ _16024;
  wire _16026 = _12298 ? coded_block[1634] : r1634;
  wire _16027 = _12296 ? _16025 : _16026;
  always @ (posedge reset or posedge clock) if (reset) r1634 <= 1'd0; else if (_12300) r1634 <= _16027;
  wire [1:0] _16028 = {_0, _672} + {_0, _3135};
  wire [1:0] _16029 = {_0, _4478} + {_0, _6207};
  wire [2:0] _16030 = {_0, _16028} + {_0, _16029};
  wire [1:0] _16031 = {_0, _8415} + {_0, _12282};
  wire [3:0] _16032 = {_0, _16030} + {_0, _0, _16031};
  wire _16033 = _12301 < _16032;
  wire _16034 = r1633 ^ _16033;
  wire _16035 = _12298 ? coded_block[1633] : r1633;
  wire _16036 = _12296 ? _16034 : _16035;
  always @ (posedge reset or posedge clock) if (reset) r1633 <= 1'd0; else if (_12300) r1633 <= _16036;
  wire [1:0] _16037 = {_0, _703} + {_0, _3742};
  wire [1:0] _16038 = {_0, _5215} + {_0, _6558};
  wire [2:0] _16039 = {_0, _16037} + {_0, _16038};
  wire [1:0] _16040 = {_0, _8288} + {_0, _10493};
  wire [3:0] _16041 = {_0, _16039} + {_0, _0, _16040};
  wire _16042 = _12301 < _16041;
  wire _16043 = r1632 ^ _16042;
  wire _16044 = _12298 ? coded_block[1632] : r1632;
  wire _16045 = _12296 ? _16043 : _16044;
  always @ (posedge reset or posedge clock) if (reset) r1632 <= 1'd0; else if (_12300) r1632 <= _16045;
  wire [1:0] _16046 = {_0, _735} + {_0, _3294};
  wire [1:0] _16047 = {_0, _5821} + {_0, _7293};
  wire [2:0] _16048 = {_0, _16046} + {_0, _16047};
  wire [1:0] _16049 = {_0, _8638} + {_0, _10366};
  wire [3:0] _16050 = {_0, _16048} + {_0, _0, _16049};
  wire _16051 = _12301 < _16050;
  wire _16052 = r1631 ^ _16051;
  wire _16053 = _12298 ? coded_block[1631] : r1631;
  wire _16054 = _12296 ? _16052 : _16053;
  always @ (posedge reset or posedge clock) if (reset) r1631 <= 1'd0; else if (_12300) r1631 <= _16054;
  wire [1:0] _16055 = {_0, _766} + {_0, _2910};
  wire [1:0] _16056 = {_0, _5373} + {_0, _7900};
  wire [2:0] _16057 = {_0, _16055} + {_0, _16056};
  wire [1:0] _16058 = {_0, _9375} + {_0, _10717};
  wire [3:0] _16059 = {_0, _16057} + {_0, _0, _16058};
  wire _16060 = _12301 < _16059;
  wire _16061 = r1630 ^ _16060;
  wire _16062 = _12298 ? coded_block[1630] : r1630;
  wire _16063 = _12296 ? _16061 : _16062;
  always @ (posedge reset or posedge clock) if (reset) r1630 <= 1'd0; else if (_12300) r1630 <= _16063;
  wire [1:0] _16064 = {_0, _831} + {_0, _2336};
  wire [1:0] _16065 = {_0, _6012} + {_0, _7069};
  wire [2:0] _16066 = {_0, _16064} + {_0, _16065};
  wire [1:0] _16067 = {_0, _9534} + {_0, _12061};
  wire [3:0] _16068 = {_0, _16066} + {_0, _0, _16067};
  wire _16069 = _12301 < _16068;
  wire _16070 = r1629 ^ _16069;
  wire _16071 = _12298 ? coded_block[1629] : r1629;
  wire _16072 = _12296 ? _16070 : _16071;
  always @ (posedge reset or posedge clock) if (reset) r1629 <= 1'd0; else if (_12300) r1629 <= _16072;
  wire [1:0] _16073 = {_0, _927} + {_0, _3549};
  wire [1:0] _16074 = {_0, _4319} + {_0, _6973};
  wire [2:0] _16075 = {_0, _16073} + {_0, _16074};
  wire [1:0] _16076 = {_0, _8574} + {_0, _12251};
  wire [3:0] _16077 = {_0, _16075} + {_0, _0, _16076};
  wire _16078 = _12301 < _16077;
  wire _16079 = r1628 ^ _16078;
  wire _16080 = _12298 ? coded_block[1628] : r1628;
  wire _16081 = _12296 ? _16079 : _16080;
  always @ (posedge reset or posedge clock) if (reset) r1628 <= 1'd0; else if (_12300) r1628 <= _16081;
  wire [1:0] _16082 = {_0, _958} + {_0, _3231};
  wire [1:0] _16083 = {_0, _5628} + {_0, _6397};
  wire [2:0] _16084 = {_0, _16082} + {_0, _16083};
  wire [1:0] _16085 = {_0, _9054} + {_0, _10654};
  wire [3:0] _16086 = {_0, _16084} + {_0, _0, _16085};
  wire _16087 = _12301 < _16086;
  wire _16088 = r1627 ^ _16087;
  wire _16089 = _12298 ? coded_block[1627] : r1627;
  wire _16090 = _12296 ? _16088 : _16089;
  always @ (posedge reset or posedge clock) if (reset) r1627 <= 1'd0; else if (_12300) r1627 <= _16090;
  wire [1:0] _16091 = {_0, _1021} + {_0, _3198};
  wire [1:0] _16092 = {_0, _5470} + {_0, _7389};
  wire [2:0] _16093 = {_0, _16091} + {_0, _16092};
  wire [1:0] _16094 = {_0, _9790} + {_0, _10558};
  wire [3:0] _16095 = {_0, _16093} + {_0, _0, _16094};
  wire _16096 = _12301 < _16095;
  wire _16097 = r1626 ^ _16096;
  wire _16098 = _12298 ? coded_block[1626] : r1626;
  wire _16099 = _12296 ? _16097 : _16098;
  always @ (posedge reset or posedge clock) if (reset) r1626 <= 1'd0; else if (_12300) r1626 <= _16099;
  wire [1:0] _16100 = {_0, _1088} + {_0, _2719};
  wire [1:0] _16101 = {_0, _5663} + {_0, _7357};
  wire [2:0] _16102 = {_0, _16100} + {_0, _16101};
  wire [1:0] _16103 = {_0, _9630} + {_0, _11550};
  wire [3:0] _16104 = {_0, _16102} + {_0, _0, _16103};
  wire _16105 = _12301 < _16104;
  wire _16106 = r1625 ^ _16105;
  wire _16107 = _12298 ? coded_block[1625] : r1625;
  wire _16108 = _12296 ? _16106 : _16107;
  always @ (posedge reset or posedge clock) if (reset) r1625 <= 1'd0; else if (_12300) r1625 <= _16108;
  wire [1:0] _16109 = {_0, _1120} + {_0, _2494};
  wire [1:0] _16110 = {_0, _4798} + {_0, _7741};
  wire [2:0] _16111 = {_0, _16109} + {_0, _16110};
  wire [1:0] _16112 = {_0, _9438} + {_0, _11708};
  wire [3:0] _16113 = {_0, _16111} + {_0, _0, _16112};
  wire _16114 = _12301 < _16113;
  wire _16115 = r1624 ^ _16114;
  wire _16116 = _12298 ? coded_block[1624] : r1624;
  wire _16117 = _12296 ? _16115 : _16116;
  always @ (posedge reset or posedge clock) if (reset) r1624 <= 1'd0; else if (_12300) r1624 <= _16117;
  wire [1:0] _16118 = {_0, _1151} + {_0, _3068};
  wire [1:0] _16119 = {_0, _4574} + {_0, _6877};
  wire [2:0] _16120 = {_0, _16118} + {_0, _16119};
  wire [1:0] _16121 = {_0, _9822} + {_0, _11516};
  wire [3:0] _16122 = {_0, _16120} + {_0, _0, _16121};
  wire _16123 = _12301 < _16122;
  wire _16124 = r1623 ^ _16123;
  wire _16125 = _12298 ? coded_block[1623] : r1623;
  wire _16126 = _12296 ? _16124 : _16125;
  always @ (posedge reset or posedge clock) if (reset) r1623 <= 1'd0; else if (_12300) r1623 <= _16126;
  wire [1:0] _16127 = {_0, _1184} + {_0, _3005};
  wire [1:0] _16128 = {_0, _5152} + {_0, _6652};
  wire [2:0] _16129 = {_0, _16127} + {_0, _16128};
  wire [1:0] _16130 = {_0, _8957} + {_0, _11900};
  wire [3:0] _16131 = {_0, _16129} + {_0, _0, _16130};
  wire _16132 = _12301 < _16131;
  wire _16133 = r1622 ^ _16132;
  wire _16134 = _12298 ? coded_block[1622] : r1622;
  wire _16135 = _12296 ? _16133 : _16134;
  always @ (posedge reset or posedge clock) if (reset) r1622 <= 1'd0; else if (_12300) r1622 <= _16135;
  wire [1:0] _16136 = {_0, _1215} + {_0, _2112};
  wire [1:0] _16137 = {_0, _5085} + {_0, _7230};
  wire [2:0] _16138 = {_0, _16136} + {_0, _16137};
  wire [1:0] _16139 = {_0, _8736} + {_0, _11038};
  wire [3:0] _16140 = {_0, _16138} + {_0, _0, _16139};
  wire _16141 = _12301 < _16140;
  wire _16142 = r1621 ^ _16141;
  wire _16143 = _12298 ? coded_block[1621] : r1621;
  wire _16144 = _12296 ? _16142 : _16143;
  always @ (posedge reset or posedge clock) if (reset) r1621 <= 1'd0; else if (_12300) r1621 <= _16144;
  wire [1:0] _16145 = {_0, _1247} + {_0, _2782};
  wire [1:0] _16146 = {_0, _4192} + {_0, _7163};
  wire [2:0] _16147 = {_0, _16145} + {_0, _16146};
  wire [1:0] _16148 = {_0, _9311} + {_0, _10814};
  wire [3:0] _16149 = {_0, _16147} + {_0, _0, _16148};
  wire _16150 = _12301 < _16149;
  wire _16151 = r1620 ^ _16150;
  wire _16152 = _12298 ? coded_block[1620] : r1620;
  wire _16153 = _12296 ? _16151 : _16152;
  always @ (posedge reset or posedge clock) if (reset) r1620 <= 1'd0; else if (_12300) r1620 <= _16153;
  wire [1:0] _16154 = {_0, _1278} + {_0, _2367};
  wire [1:0] _16155 = {_0, _4861} + {_0, _6270};
  wire [2:0] _16156 = {_0, _16154} + {_0, _16155};
  wire [1:0] _16157 = {_0, _9248} + {_0, _11389};
  wire [3:0] _16158 = {_0, _16156} + {_0, _0, _16157};
  wire _16159 = _12301 < _16158;
  wire _16160 = r1619 ^ _16159;
  wire _16161 = _12298 ? coded_block[1619] : r1619;
  wire _16162 = _12296 ? _16160 : _16161;
  always @ (posedge reset or posedge clock) if (reset) r1619 <= 1'd0; else if (_12300) r1619 <= _16162;
  wire [1:0] _16163 = {_0, _1312} + {_0, _4091};
  wire [1:0] _16164 = {_0, _4447} + {_0, _6942};
  wire [2:0] _16165 = {_0, _16163} + {_0, _16164};
  wire [1:0] _16166 = {_0, _8352} + {_0, _11326};
  wire [3:0] _16167 = {_0, _16165} + {_0, _0, _16166};
  wire _16168 = _12301 < _16167;
  wire _16169 = r1618 ^ _16168;
  wire _16170 = _12298 ? coded_block[1618] : r1618;
  wire _16171 = _12296 ? _16169 : _16170;
  always @ (posedge reset or posedge clock) if (reset) r1618 <= 1'd0; else if (_12300) r1618 <= _16171;
  wire [1:0] _16172 = {_0, _1343} + {_0, _3037};
  wire [1:0] _16173 = {_0, _4160} + {_0, _6525};
  wire [2:0] _16174 = {_0, _16172} + {_0, _16173};
  wire [1:0] _16175 = {_0, _9022} + {_0, _10430};
  wire [3:0] _16176 = {_0, _16174} + {_0, _0, _16175};
  wire _16177 = _12301 < _16176;
  wire _16178 = r1617 ^ _16177;
  wire _16179 = _12298 ? coded_block[1617] : r1617;
  wire _16180 = _12296 ? _16178 : _16179;
  always @ (posedge reset or posedge clock) if (reset) r1617 <= 1'd0; else if (_12300) r1617 <= _16180;
  wire [1:0] _16181 = {_0, _1375} + {_0, _2526};
  wire [1:0] _16182 = {_0, _5116} + {_0, _6239};
  wire [2:0] _16183 = {_0, _16181} + {_0, _16182};
  wire [1:0] _16184 = {_0, _8607} + {_0, _11101};
  wire [3:0] _16185 = {_0, _16183} + {_0, _0, _16184};
  wire _16186 = _12301 < _16185;
  wire _16187 = r1616 ^ _16186;
  wire _16188 = _12298 ? coded_block[1616] : r1616;
  wire _16189 = _12296 ? _16187 : _16188;
  always @ (posedge reset or posedge clock) if (reset) r1616 <= 1'd0; else if (_12300) r1616 <= _16189;
  wire [1:0] _16190 = {_0, _1406} + {_0, _3517};
  wire [1:0] _16191 = {_0, _4605} + {_0, _7199};
  wire [2:0] _16192 = {_0, _16190} + {_0, _16191};
  wire [1:0] _16193 = {_0, _8319} + {_0, _10685};
  wire [3:0] _16194 = {_0, _16192} + {_0, _0, _16193};
  wire _16195 = _12301 < _16194;
  wire _16196 = r1615 ^ _16195;
  wire _16197 = _12298 ? coded_block[1615] : r1615;
  wire _16198 = _12296 ? _16196 : _16197;
  always @ (posedge reset or posedge clock) if (reset) r1615 <= 1'd0; else if (_12300) r1615 <= _16198;
  wire [1:0] _16199 = {_0, _1439} + {_0, _2271};
  wire [1:0] _16200 = {_0, _5597} + {_0, _6687};
  wire [2:0] _16201 = {_0, _16199} + {_0, _16200};
  wire [1:0] _16202 = {_0, _9279} + {_0, _10399};
  wire [3:0] _16203 = {_0, _16201} + {_0, _0, _16202};
  wire _16204 = _12301 < _16203;
  wire _16205 = r1614 ^ _16204;
  wire _16206 = _12298 ? coded_block[1614] : r1614;
  wire _16207 = _12296 ? _16205 : _16206;
  always @ (posedge reset or posedge clock) if (reset) r1614 <= 1'd0; else if (_12300) r1614 <= _16207;
  wire [1:0] _16208 = {_0, _1502} + {_0, _2974};
  wire [1:0] _16209 = {_0, _5534} + {_0, _6431};
  wire [2:0] _16210 = {_0, _16208} + {_0, _16209};
  wire [1:0] _16211 = {_0, _9759} + {_0, _10846};
  wire [3:0] _16212 = {_0, _16210} + {_0, _0, _16211};
  wire _16213 = _12301 < _16212;
  wire _16214 = r1613 ^ _16213;
  wire _16215 = _12298 ? coded_block[1613] : r1613;
  wire _16216 = _12296 ? _16214 : _16215;
  always @ (posedge reset or posedge clock) if (reset) r1613 <= 1'd0; else if (_12300) r1613 <= _16216;
  wire [1:0] _16217 = {_0, _1533} + {_0, _3104};
  wire [1:0] _16218 = {_0, _5053} + {_0, _7612};
  wire [2:0] _16219 = {_0, _16217} + {_0, _16218};
  wire [1:0] _16220 = {_0, _8511} + {_0, _11837};
  wire [3:0] _16221 = {_0, _16219} + {_0, _0, _16220};
  wire _16222 = _12301 < _16221;
  wire _16223 = r1612 ^ _16222;
  wire _16224 = _12298 ? coded_block[1612] : r1612;
  wire _16225 = _12296 ? _16223 : _16224;
  always @ (posedge reset or posedge clock) if (reset) r1612 <= 1'd0; else if (_12300) r1612 <= _16225;
  wire [1:0] _16226 = {_0, _1599} + {_0, _3678};
  wire [1:0] _16227 = {_0, _4511} + {_0, _7262};
  wire [2:0] _16228 = {_0, _16226} + {_0, _16227};
  wire [1:0] _16229 = {_0, _9212} + {_0, _11771};
  wire [3:0] _16230 = {_0, _16228} + {_0, _0, _16229};
  wire _16231 = _12301 < _16230;
  wire _16232 = r1611 ^ _16231;
  wire _16233 = _12298 ? coded_block[1611] : r1611;
  wire _16234 = _12296 ? _16232 : _16233;
  always @ (posedge reset or posedge clock) if (reset) r1611 <= 1'd0; else if (_12300) r1611 <= _16234;
  wire [1:0] _16235 = {_0, _1631} + {_0, _3646};
  wire [1:0] _16236 = {_0, _5757} + {_0, _6589};
  wire [2:0] _16237 = {_0, _16235} + {_0, _16236};
  wire [1:0] _16238 = {_0, _9342} + {_0, _11295};
  wire [3:0] _16239 = {_0, _16237} + {_0, _0, _16238};
  wire _16240 = _12301 < _16239;
  wire _16241 = r1610 ^ _16240;
  wire _16242 = _12298 ? coded_block[1610] : r1610;
  wire _16243 = _12296 ? _16241 : _16242;
  always @ (posedge reset or posedge clock) if (reset) r1610 <= 1'd0; else if (_12300) r1610 <= _16243;
  wire [1:0] _16244 = {_0, _1662} + {_0, _2463};
  wire [1:0] _16245 = {_0, _5726} + {_0, _7837};
  wire [2:0] _16246 = {_0, _16244} + {_0, _16245};
  wire [1:0] _16247 = {_0, _8670} + {_0, _11422};
  wire [3:0] _16248 = {_0, _16246} + {_0, _0, _16247};
  wire _16249 = _12301 < _16248;
  wire _16250 = r1609 ^ _16249;
  wire _16251 = _12298 ? coded_block[1609] : r1609;
  wire _16252 = _12296 ? _16250 : _16251;
  always @ (posedge reset or posedge clock) if (reset) r1609 <= 1'd0; else if (_12300) r1609 <= _16252;
  wire [1:0] _16253 = {_0, _1758} + {_0, _3997};
  wire [1:0] _16254 = {_0, _4223} + {_0, _6908};
  wire [2:0] _16255 = {_0, _16253} + {_0, _16254};
  wire [1:0] _16256 = {_0, _8701} + {_0, _11964};
  wire [3:0] _16257 = {_0, _16255} + {_0, _0, _16256};
  wire _16258 = _12301 < _16257;
  wire _16259 = r1608 ^ _16258;
  wire _16260 = _12298 ? coded_block[1608] : r1608;
  wire _16261 = _12296 ? _16259 : _16260;
  always @ (posedge reset or posedge clock) if (reset) r1608 <= 1'd0; else if (_12300) r1608 <= _16261;
  wire [1:0] _16262 = {_0, _34} + {_0, _2239};
  wire [1:0] _16263 = {_0, _4319} + {_0, _6397};
  wire [2:0] _16264 = {_0, _16262} + {_0, _16263};
  wire [1:0] _16265 = {_0, _8480} + {_0, _10558};
  wire [3:0] _16266 = {_0, _16264} + {_0, _0, _16265};
  wire _16267 = _12301 < _16266;
  wire _16268 = r1607 ^ _16267;
  wire _16269 = _12298 ? coded_block[1607] : r1607;
  wire _16270 = _12296 ? _16268 : _16269;
  always @ (posedge reset or posedge clock) if (reset) r1607 <= 1'd0; else if (_12300) r1607 <= _16270;
  wire [1:0] _16271 = {_0, _1120} + {_0, _2144};
  wire [1:0] _16272 = {_0, _5628} + {_0, _6973};
  wire [2:0] _16273 = {_0, _16271} + {_0, _16272};
  wire [1:0] _16274 = {_0, _8701} + {_0, _10910};
  wire [3:0] _16275 = {_0, _16273} + {_0, _0, _16274};
  wire _16276 = _12301 < _16275;
  wire _16277 = r1606 ^ _16276;
  wire _16278 = _12298 ? coded_block[1606] : r1606;
  wire _16279 = _12296 ? _16277 : _16278;
  always @ (posedge reset or posedge clock) if (reset) r1606 <= 1'd0; else if (_12300) r1606 <= _16279;
  wire [1:0] _16280 = {_0, _1151} + {_0, _3709};
  wire [1:0] _16281 = {_0, _4223} + {_0, _7710};
  wire [2:0] _16282 = {_0, _16280} + {_0, _16281};
  wire [1:0] _16283 = {_0, _9054} + {_0, _10783};
  wire [3:0] _16284 = {_0, _16282} + {_0, _0, _16283};
  wire _16285 = _12301 < _16284;
  wire _16286 = r1605 ^ _16285;
  wire _16287 = _12298 ? coded_block[1605] : r1605;
  wire _16288 = _12296 ? _16286 : _16287;
  always @ (posedge reset or posedge clock) if (reset) r1605 <= 1'd0; else if (_12300) r1605 <= _16288;
  wire [1:0] _16289 = {_0, _1184} + {_0, _3325};
  wire [1:0] _16290 = {_0, _5790} + {_0, _6303};
  wire [2:0] _16291 = {_0, _16289} + {_0, _16290};
  wire [1:0] _16292 = {_0, _9790} + {_0, _11132};
  wire [3:0] _16293 = {_0, _16291} + {_0, _0, _16292};
  wire _16294 = _12301 < _16293;
  wire _16295 = r1604 ^ _16294;
  wire _16296 = _12298 ? coded_block[1604] : r1604;
  wire _16297 = _12296 ? _16295 : _16296;
  always @ (posedge reset or posedge clock) if (reset) r1604 <= 1'd0; else if (_12300) r1604 <= _16297;
  wire [1:0] _16298 = {_0, _1215} + {_0, _2336};
  wire [1:0] _16299 = {_0, _5407} + {_0, _7868};
  wire [2:0] _16300 = {_0, _16298} + {_0, _16299};
  wire [1:0] _16301 = {_0, _8383} + {_0, _11869};
  wire [3:0] _16302 = {_0, _16300} + {_0, _0, _16301};
  wire _16303 = _12301 < _16302;
  wire _16304 = r1603 ^ _16303;
  wire _16305 = _12298 ? coded_block[1603] : r1603;
  wire _16306 = _12296 ? _16304 : _16305;
  always @ (posedge reset or posedge clock) if (reset) r1603 <= 1'd0; else if (_12300) r1603 <= _16306;
  wire [1:0] _16307 = {_0, _1278} + {_0, _3231};
  wire [1:0] _16308 = {_0, _4830} + {_0, _6494};
  wire [2:0] _16309 = {_0, _16307} + {_0, _16308};
  wire [1:0] _16310 = {_0, _9566} + {_0, _12027};
  wire [3:0] _16311 = {_0, _16309} + {_0, _0, _16310};
  wire _16312 = _12301 < _16311;
  wire _16313 = r1602 ^ _16312;
  wire _16314 = _12298 ? coded_block[1602] : r1602;
  wire _16315 = _12296 ? _16313 : _16314;
  always @ (posedge reset or posedge clock) if (reset) r1602 <= 1'd0; else if (_12300) r1602 <= _16315;
  wire [1:0] _16316 = {_0, _1312} + {_0, _2655};
  wire [1:0] _16317 = {_0, _5310} + {_0, _6908};
  wire [2:0] _16318 = {_0, _16316} + {_0, _16317};
  wire [1:0] _16319 = {_0, _8574} + {_0, _11644};
  wire [3:0] _16320 = {_0, _16318} + {_0, _0, _16319};
  wire _16321 = _12301 < _16320;
  wire _16322 = r1601 ^ _16321;
  wire _16323 = _12298 ? coded_block[1601] : r1601;
  wire _16324 = _12296 ? _16322 : _16323;
  always @ (posedge reset or posedge clock) if (reset) r1601 <= 1'd0; else if (_12300) r1601 <= _16324;
  wire [1:0] _16325 = {_0, _1343} + {_0, _3964};
  wire [1:0] _16326 = {_0, _4734} + {_0, _7389};
  wire [2:0] _16327 = {_0, _16325} + {_0, _16326};
  wire [1:0] _16328 = {_0, _8991} + {_0, _10654};
  wire [3:0] _16329 = {_0, _16327} + {_0, _0, _16328};
  wire _16330 = _12301 < _16329;
  wire _16331 = r1600 ^ _16330;
  wire _16332 = _12298 ? coded_block[1600] : r1600;
  wire _16333 = _12296 ? _16331 : _16332;
  always @ (posedge reset or posedge clock) if (reset) r1600 <= 1'd0; else if (_12300) r1600 <= _16333;
  wire [1:0] _16334 = {_0, _1406} + {_0, _3805};
  wire [1:0] _16335 = {_0, _5726} + {_0, _8123};
  wire [2:0] _16336 = {_0, _16334} + {_0, _16335};
  wire [1:0] _16337 = {_0, _8894} + {_0, _11550};
  wire [3:0] _16338 = {_0, _16336} + {_0, _0, _16337};
  wire _16339 = _12301 < _16338;
  wire _16340 = r1599 ^ _16339;
  wire _16341 = _12298 ? coded_block[1599] : r1599;
  wire _16342 = _12296 ? _16340 : _16341;
  always @ (posedge reset or posedge clock) if (reset) r1599 <= 1'd0; else if (_12300) r1599 <= _16342;
  wire [1:0] _16343 = {_0, _1439} + {_0, _3615};
  wire [1:0] _16344 = {_0, _5884} + {_0, _7804};
  wire [2:0] _16345 = {_0, _16343} + {_0, _16344};
  wire [1:0] _16346 = {_0, _10204} + {_0, _10973};
  wire [3:0] _16347 = {_0, _16345} + {_0, _0, _16346};
  wire _16348 = _12301 < _16347;
  wire _16349 = r1598 ^ _16348;
  wire _16350 = _12298 ? coded_block[1598] : r1598;
  wire _16351 = _12296 ? _16349 : _16350;
  always @ (posedge reset or posedge clock) if (reset) r1598 <= 1'd0; else if (_12300) r1598 <= _16351;
  wire [1:0] _16352 = {_0, _1470} + {_0, _3997};
  wire [1:0] _16353 = {_0, _5694} + {_0, _7965};
  wire [2:0] _16354 = {_0, _16352} + {_0, _16353};
  wire [1:0] _16355 = {_0, _9886} + {_0, _12282};
  wire [3:0] _16356 = {_0, _16354} + {_0, _0, _16355};
  wire _16357 = _12301 < _16356;
  wire _16358 = r1597 ^ _16357;
  wire _16359 = _12298 ? coded_block[1597] : r1597;
  wire _16360 = _12296 ? _16358 : _16359;
  always @ (posedge reset or posedge clock) if (reset) r1597 <= 1'd0; else if (_12300) r1597 <= _16360;
  wire [1:0] _16361 = {_0, _1502} + {_0, _3135};
  wire [1:0] _16362 = {_0, _6076} + {_0, _7773};
  wire [2:0] _16363 = {_0, _16361} + {_0, _16362};
  wire [1:0] _16364 = {_0, _10045} + {_0, _11964};
  wire [3:0] _16365 = {_0, _16363} + {_0, _0, _16364};
  wire _16366 = _12301 < _16365;
  wire _16367 = r1596 ^ _16366;
  wire _16368 = _12298 ? coded_block[1596] : r1596;
  wire _16369 = _12296 ? _16367 : _16368;
  always @ (posedge reset or posedge clock) if (reset) r1596 <= 1'd0; else if (_12300) r1596 <= _16369;
  wire [1:0] _16370 = {_0, _1568} + {_0, _3486};
  wire [1:0] _16371 = {_0, _4989} + {_0, _7293};
  wire [2:0] _16372 = {_0, _16370} + {_0, _16371};
  wire [1:0] _16373 = {_0, _10235} + {_0, _11933};
  wire [3:0] _16374 = {_0, _16372} + {_0, _0, _16373};
  wire _16375 = _12301 < _16374;
  wire _16376 = r1595 ^ _16375;
  wire _16377 = _12298 ? coded_block[1595] : r1595;
  wire _16378 = _12296 ? _16376 : _16377;
  always @ (posedge reset or posedge clock) if (reset) r1595 <= 1'd0; else if (_12300) r1595 <= _16378;
  wire [1:0] _16379 = {_0, _1599} + {_0, _3422};
  wire [1:0] _16380 = {_0, _5565} + {_0, _7069};
  wire [2:0] _16381 = {_0, _16379} + {_0, _16380};
  wire [1:0] _16382 = {_0, _9375} + {_0, _10303};
  wire [3:0] _16383 = {_0, _16381} + {_0, _0, _16382};
  wire _16384 = _12301 < _16383;
  wire _16385 = r1594 ^ _16384;
  wire _16386 = _12298 ? coded_block[1594] : r1594;
  wire _16387 = _12296 ? _16385 : _16386;
  always @ (posedge reset or posedge clock) if (reset) r1594 <= 1'd0; else if (_12300) r1594 <= _16387;
  wire [1:0] _16388 = {_0, _1631} + {_0, _2526};
  wire [1:0] _16389 = {_0, _5501} + {_0, _7644};
  wire [2:0] _16390 = {_0, _16388} + {_0, _16389};
  wire [1:0] _16391 = {_0, _9149} + {_0, _11453};
  wire [3:0] _16392 = {_0, _16390} + {_0, _0, _16391};
  wire _16393 = _12301 < _16392;
  wire _16394 = r1593 ^ _16393;
  wire _16395 = _12298 ? coded_block[1593] : r1593;
  wire _16396 = _12296 ? _16394 : _16395;
  always @ (posedge reset or posedge clock) if (reset) r1593 <= 1'd0; else if (_12300) r1593 <= _16396;
  wire [1:0] _16397 = {_0, _1662} + {_0, _3198};
  wire [1:0] _16398 = {_0, _4605} + {_0, _7581};
  wire [2:0] _16399 = {_0, _16397} + {_0, _16398};
  wire [1:0] _16400 = {_0, _9724} + {_0, _11228};
  wire [3:0] _16401 = {_0, _16399} + {_0, _0, _16400};
  wire _16402 = _12301 < _16401;
  wire _16403 = r1592 ^ _16402;
  wire _16404 = _12298 ? coded_block[1592] : r1592;
  wire _16405 = _12296 ? _16403 : _16404;
  always @ (posedge reset or posedge clock) if (reset) r1592 <= 1'd0; else if (_12300) r1592 <= _16405;
  wire [1:0] _16406 = {_0, _1789} + {_0, _2941};
  wire [1:0] _16407 = {_0, _5534} + {_0, _6652};
  wire [2:0] _16408 = {_0, _16406} + {_0, _16407};
  wire [1:0] _16409 = {_0, _9022} + {_0, _11516};
  wire [3:0] _16410 = {_0, _16408} + {_0, _0, _16409};
  wire _16411 = _12301 < _16410;
  wire _16412 = r1591 ^ _16411;
  wire _16413 = _12298 ? coded_block[1591] : r1591;
  wire _16414 = _12296 ? _16412 : _16413;
  always @ (posedge reset or posedge clock) if (reset) r1591 <= 1'd0; else if (_12300) r1591 <= _16414;
  wire [1:0] _16415 = {_0, _1854} + {_0, _2686};
  wire [1:0] _16416 = {_0, _6012} + {_0, _7100};
  wire [2:0] _16417 = {_0, _16415} + {_0, _16416};
  wire [1:0] _16418 = {_0, _9693} + {_0, _10814};
  wire [3:0] _16419 = {_0, _16417} + {_0, _0, _16418};
  wire _16420 = _12301 < _16419;
  wire _16421 = r1590 ^ _16420;
  wire _16422 = _12298 ? coded_block[1590] : r1590;
  wire _16423 = _12296 ? _16421 : _16422;
  always @ (posedge reset or posedge clock) if (reset) r1590 <= 1'd0; else if (_12300) r1590 <= _16423;
  wire [1:0] _16424 = {_0, _1886} + {_0, _3870};
  wire [1:0] _16425 = {_0, _4767} + {_0, _8092};
  wire [2:0] _16426 = {_0, _16424} + {_0, _16425};
  wire [1:0] _16427 = {_0, _9181} + {_0, _11771};
  wire [3:0] _16428 = {_0, _16426} + {_0, _0, _16427};
  wire _16429 = _12301 < _16428;
  wire _16430 = r1589 ^ _16429;
  wire _16431 = _12298 ? coded_block[1589] : r1589;
  wire _16432 = _12296 ? _16430 : _16431;
  always @ (posedge reset or posedge clock) if (reset) r1589 <= 1'd0; else if (_12300) r1589 <= _16432;
  wire [1:0] _16433 = {_0, _1950} + {_0, _3517};
  wire [1:0] _16434 = {_0, _5470} + {_0, _8028};
  wire [2:0] _16435 = {_0, _16433} + {_0, _16434};
  wire [1:0] _16436 = {_0, _8926} + {_0, _12251};
  wire [3:0] _16437 = {_0, _16435} + {_0, _0, _16436};
  wire _16438 = _12301 < _16437;
  wire _16439 = r1588 ^ _16438;
  wire _16440 = _12298 ? coded_block[1588] : r1588;
  wire _16441 = _12296 ? _16439 : _16440;
  always @ (posedge reset or posedge clock) if (reset) r1588 <= 1'd0; else if (_12300) r1588 <= _16441;
  wire [1:0] _16442 = {_0, _2013} + {_0, _4091};
  wire [1:0] _16443 = {_0, _4926} + {_0, _7675};
  wire [2:0] _16444 = {_0, _16442} + {_0, _16443};
  wire [1:0] _16445 = {_0, _9630} + {_0, _12188};
  wire [3:0] _16446 = {_0, _16444} + {_0, _0, _16445};
  wire _16447 = _12301 < _16446;
  wire _16448 = r1587 ^ _16447;
  wire _16449 = _12298 ? coded_block[1587] : r1587;
  wire _16450 = _12296 ? _16448 : _16449;
  always @ (posedge reset or posedge clock) if (reset) r1587 <= 1'd0; else if (_12300) r1587 <= _16450;
  wire [1:0] _16451 = {_0, _2044} + {_0, _4060};
  wire [1:0] _16452 = {_0, _4160} + {_0, _7005};
  wire [2:0] _16453 = {_0, _16451} + {_0, _16452};
  wire [1:0] _16454 = {_0, _9759} + {_0, _11708};
  wire [3:0] _16455 = {_0, _16453} + {_0, _0, _16454};
  wire _16456 = _12301 < _16455;
  wire _16457 = r1586 ^ _16456;
  wire _16458 = _12298 ? coded_block[1586] : r1586;
  wire _16459 = _12296 ? _16457 : _16458;
  always @ (posedge reset or posedge clock) if (reset) r1586 <= 1'd0; else if (_12300) r1586 <= _16459;
  wire [1:0] _16460 = {_0, _65} + {_0, _2878};
  wire [1:0] _16461 = {_0, _6139} + {_0, _6239};
  wire [2:0] _16462 = {_0, _16460} + {_0, _16461};
  wire [1:0] _16463 = {_0, _9085} + {_0, _11837};
  wire [3:0] _16464 = {_0, _16462} + {_0, _0, _16463};
  wire _16465 = _12301 < _16464;
  wire _16466 = r1585 ^ _16465;
  wire _16467 = _12298 ? coded_block[1585] : r1585;
  wire _16468 = _12296 ? _16466 : _16467;
  always @ (posedge reset or posedge clock) if (reset) r1585 <= 1'd0; else if (_12300) r1585 <= _16468;
  wire [1:0] _16469 = {_0, _97} + {_0, _3167};
  wire [1:0] _16470 = {_0, _4958} + {_0, _6207};
  wire [2:0] _16471 = {_0, _16469} + {_0, _16470};
  wire [1:0] _16472 = {_0, _8319} + {_0, _11165};
  wire [3:0] _16473 = {_0, _16471} + {_0, _0, _16472};
  wire _16474 = _12301 < _16473;
  wire _16475 = r1584 ^ _16474;
  wire _16476 = _12298 ? coded_block[1584] : r1584;
  wire _16477 = _12296 ? _16475 : _16476;
  always @ (posedge reset or posedge clock) if (reset) r1584 <= 1'd0; else if (_12300) r1584 <= _16477;
  wire [1:0] _16478 = {_0, _161} + {_0, _2399};
  wire [1:0] _16479 = {_0, _4640} + {_0, _7326};
  wire [2:0] _16480 = {_0, _16478} + {_0, _16479};
  wire [1:0] _16481 = {_0, _9118} + {_0, _10366};
  wire [3:0] _16482 = {_0, _16480} + {_0, _0, _16481};
  wire _16483 = _12301 < _16482;
  wire _16484 = r1583 ^ _16483;
  wire _16485 = _12298 ? coded_block[1583] : r1583;
  wire _16486 = _12296 ? _16484 : _16485;
  always @ (posedge reset or posedge clock) if (reset) r1583 <= 1'd0; else if (_12300) r1583 <= _16486;
  wire [1:0] _16487 = {_0, _192} + {_0, _2081};
  wire [1:0] _16488 = {_0, _4478} + {_0, _6718};
  wire [2:0] _16489 = {_0, _16487} + {_0, _16488};
  wire [1:0] _16490 = {_0, _9406} + {_0, _11196};
  wire [3:0] _16491 = {_0, _16489} + {_0, _0, _16490};
  wire _16492 = _12301 < _16491;
  wire _16493 = r1582 ^ _16492;
  wire _16494 = _12298 ? coded_block[1582] : r1582;
  wire _16495 = _12296 ? _16493 : _16494;
  always @ (posedge reset or posedge clock) if (reset) r1582 <= 1'd0; else if (_12300) r1582 <= _16495;
  wire [1:0] _16496 = {_0, _224} + {_0, _2430};
  wire [1:0] _16497 = {_0, _4129} + {_0, _6558};
  wire [2:0] _16498 = {_0, _16496} + {_0, _16497};
  wire [1:0] _16499 = {_0, _8799} + {_0, _11485};
  wire [3:0] _16500 = {_0, _16498} + {_0, _0, _16499};
  wire _16501 = _12301 < _16500;
  wire _16502 = r1581 ^ _16501;
  wire _16503 = _12298 ? coded_block[1581] : r1581;
  wire _16504 = _12296 ? _16502 : _16503;
  always @ (posedge reset or posedge clock) if (reset) r1581 <= 1'd0; else if (_12300) r1581 <= _16504;
  wire [1:0] _16505 = {_0, _255} + {_0, _2623};
  wire [1:0] _16506 = {_0, _4511} + {_0, _6176};
  wire [2:0] _16507 = {_0, _16505} + {_0, _16506};
  wire [1:0] _16508 = {_0, _8638} + {_0, _10877};
  wire [3:0] _16509 = {_0, _16507} + {_0, _0, _16508};
  wire _16510 = _12301 < _16509;
  wire _16511 = r1580 ^ _16510;
  wire _16512 = _12298 ? coded_block[1580] : r1580;
  wire _16513 = _12296 ? _16511 : _16512;
  always @ (posedge reset or posedge clock) if (reset) r1580 <= 1'd0; else if (_12300) r1580 <= _16513;
  wire [1:0] _16514 = {_0, _320} + {_0, _3005};
  wire [1:0] _16515 = {_0, _5342} + {_0, _6781};
  wire [2:0] _16516 = {_0, _16514} + {_0, _16515};
  wire [1:0] _16517 = {_0, _8670} + {_0, _10272};
  wire [3:0] _16518 = {_0, _16516} + {_0, _0, _16517};
  wire _16519 = _12301 < _16518;
  wire _16520 = r1579 ^ _16519;
  wire _16521 = _12298 ? coded_block[1579] : r1579;
  wire _16522 = _12296 ? _16520 : _16521;
  always @ (posedge reset or posedge clock) if (reset) r1579 <= 1'd0; else if (_12300) r1579 <= _16522;
  wire [1:0] _16523 = {_0, _352} + {_0, _2208};
  wire [1:0] _16524 = {_0, _5085} + {_0, _7420};
  wire [2:0] _16525 = {_0, _16523} + {_0, _16524};
  wire [1:0] _16526 = {_0, _8863} + {_0, _10748};
  wire [3:0] _16527 = {_0, _16525} + {_0, _0, _16526};
  wire _16528 = _12301 < _16527;
  wire _16529 = r1578 ^ _16528;
  wire _16530 = _12298 ? coded_block[1578] : r1578;
  wire _16531 = _12296 ? _16529 : _16530;
  always @ (posedge reset or posedge clock) if (reset) r1578 <= 1'd0; else if (_12300) r1578 <= _16531;
  wire [1:0] _16532 = {_0, _383} + {_0, _2271};
  wire [1:0] _16533 = {_0, _4287} + {_0, _7163};
  wire [2:0] _16534 = {_0, _16532} + {_0, _16533};
  wire [1:0] _16535 = {_0, _9503} + {_0, _10941};
  wire [3:0] _16536 = {_0, _16534} + {_0, _0, _16535};
  wire _16537 = _12301 < _16536;
  wire _16538 = r1577 ^ _16537;
  wire _16539 = _12298 ? coded_block[1577] : r1577;
  wire _16540 = _12296 ? _16538 : _16539;
  always @ (posedge reset or posedge clock) if (reset) r1577 <= 1'd0; else if (_12300) r1577 <= _16540;
  wire [1:0] _16541 = {_0, _447} + {_0, _3773};
  wire [1:0] _16542 = {_0, _5152} + {_0, _6431};
  wire [2:0] _16543 = {_0, _16541} + {_0, _16542};
  wire [1:0] _16544 = {_0, _8446} + {_0, _11326};
  wire [3:0] _16545 = {_0, _16543} + {_0, _0, _16544};
  wire _16546 = _12301 < _16545;
  wire _16547 = r1576 ^ _16546;
  wire _16548 = _12298 ? coded_block[1576] : r1576;
  wire _16549 = _12296 ? _16547 : _16548;
  always @ (posedge reset or posedge clock) if (reset) r1576 <= 1'd0; else if (_12300) r1576 <= _16549;
  wire [1:0] _16550 = {_0, _34} + {_0, _3135};
  wire [1:0] _16551 = {_0, _5215} + {_0, _7293};
  wire [2:0] _16552 = {_0, _16550} + {_0, _16551};
  wire [1:0] _16553 = {_0, _9375} + {_0, _11453};
  wire [3:0] _16554 = {_0, _16552} + {_0, _0, _16553};
  wire _16555 = _12301 < _16554;
  wire _16556 = r1575 ^ _16555;
  wire _16557 = _12298 ? coded_block[1575] : r1575;
  wire _16558 = _12296 ? _16556 : _16557;
  always @ (posedge reset or posedge clock) if (reset) r1575 <= 1'd0; else if (_12300) r1575 <= _16558;
  wire [1:0] _16559 = {_0, _1088} + {_0, _2081};
  wire [1:0] _16560 = {_0, _5373} + {_0, _7612};
  wire [2:0] _16561 = {_0, _16559} + {_0, _16560};
  wire [1:0] _16562 = {_0, _8288} + {_0, _12092};
  wire [3:0] _16563 = {_0, _16561} + {_0, _0, _16562};
  wire _16564 = _12301 < _16563;
  wire _16565 = r1574 ^ _16564;
  wire _16566 = _12298 ? coded_block[1574] : r1574;
  wire _16567 = _12296 ? _16565 : _16566;
  always @ (posedge reset or posedge clock) if (reset) r1574 <= 1'd0; else if (_12300) r1574 <= _16567;
  wire [1:0] _16568 = {_0, _1120} + {_0, _3325};
  wire [1:0] _16569 = {_0, _4129} + {_0, _7454};
  wire [2:0] _16570 = {_0, _16568} + {_0, _16569};
  wire [1:0] _16571 = {_0, _9693} + {_0, _10366};
  wire [3:0] _16572 = {_0, _16570} + {_0, _0, _16571};
  wire _16573 = _12301 < _16572;
  wire _16574 = r1573 ^ _16573;
  wire _16575 = _12298 ? coded_block[1573] : r1573;
  wire _16576 = _12296 ? _16574 : _16575;
  always @ (posedge reset or posedge clock) if (reset) r1573 <= 1'd0; else if (_12300) r1573 <= _16576;
  wire [1:0] _16577 = {_0, _1215} + {_0, _3901};
  wire [1:0] _16578 = {_0, _4223} + {_0, _7675};
  wire [2:0] _16579 = {_0, _16577} + {_0, _16578};
  wire [1:0] _16580 = {_0, _9566} + {_0, _10272};
  wire [3:0] _16581 = {_0, _16579} + {_0, _0, _16580};
  wire _16582 = _12301 < _16581;
  wire _16583 = r1572 ^ _16582;
  wire _16584 = _12298 ? coded_block[1572] : r1572;
  wire _16585 = _12296 ? _16583 : _16584;
  always @ (posedge reset or posedge clock) if (reset) r1572 <= 1'd0; else if (_12300) r1572 <= _16585;
  wire [1:0] _16586 = {_0, _1247} + {_0, _3104};
  wire [1:0] _16587 = {_0, _5981} + {_0, _6303};
  wire [2:0] _16588 = {_0, _16586} + {_0, _16587};
  wire [1:0] _16589 = {_0, _9759} + {_0, _11644};
  wire [3:0] _16590 = {_0, _16588} + {_0, _0, _16589};
  wire _16591 = _12301 < _16590;
  wire _16592 = r1571 ^ _16591;
  wire _16593 = _12298 ? coded_block[1571] : r1571;
  wire _16594 = _12296 ? _16592 : _16593;
  always @ (posedge reset or posedge clock) if (reset) r1571 <= 1'd0; else if (_12300) r1571 <= _16594;
  wire [1:0] _16595 = {_0, _1278} + {_0, _3167};
  wire [1:0] _16596 = {_0, _5183} + {_0, _8059};
  wire [2:0] _16597 = {_0, _16595} + {_0, _16596};
  wire [1:0] _16598 = {_0, _8383} + {_0, _11837};
  wire [3:0] _16599 = {_0, _16597} + {_0, _0, _16598};
  wire _16600 = _12301 < _16599;
  wire _16601 = r1570 ^ _16600;
  wire _16602 = _12298 ? coded_block[1570] : r1570;
  wire _16603 = _12296 ? _16601 : _16602;
  always @ (posedge reset or posedge clock) if (reset) r1570 <= 1'd0; else if (_12300) r1570 <= _16603;
  wire [1:0] _16604 = {_0, _1312} + {_0, _3964};
  wire [1:0] _16605 = {_0, _5246} + {_0, _7262};
  wire [2:0] _16606 = {_0, _16604} + {_0, _16605};
  wire [1:0] _16607 = {_0, _10141} + {_0, _10462};
  wire [3:0] _16608 = {_0, _16606} + {_0, _0, _16607};
  wire _16609 = _12301 < _16608;
  wire _16610 = r1569 ^ _16609;
  wire _16611 = _12298 ? coded_block[1569] : r1569;
  wire _16612 = _12296 ? _16610 : _16611;
  always @ (posedge reset or posedge clock) if (reset) r1569 <= 1'd0; else if (_12300) r1569 <= _16612;
  wire [1:0] _16613 = {_0, _1343} + {_0, _2655};
  wire [1:0] _16614 = {_0, _6045} + {_0, _7326};
  wire [2:0] _16615 = {_0, _16613} + {_0, _16614};
  wire [1:0] _16616 = {_0, _9342} + {_0, _12219};
  wire [3:0] _16617 = {_0, _16615} + {_0, _0, _16616};
  wire _16618 = _12301 < _16617;
  wire _16619 = r1568 ^ _16618;
  wire _16620 = _12298 ? coded_block[1568] : r1568;
  wire _16621 = _12296 ? _16619 : _16620;
  always @ (posedge reset or posedge clock) if (reset) r1568 <= 1'd0; else if (_12300) r1568 <= _16621;
  wire [1:0] _16622 = {_0, _1375} + {_0, _2557};
  wire [1:0] _16623 = {_0, _4734} + {_0, _8123};
  wire [2:0] _16624 = {_0, _16622} + {_0, _16623};
  wire [1:0] _16625 = {_0, _9406} + {_0, _11422};
  wire [3:0] _16626 = {_0, _16624} + {_0, _0, _16625};
  wire _16627 = _12301 < _16626;
  wire _16628 = r1567 ^ _16627;
  wire _16629 = _12298 ? coded_block[1567] : r1567;
  wire _16630 = _12296 ? _16628 : _16629;
  always @ (posedge reset or posedge clock) if (reset) r1567 <= 1'd0; else if (_12300) r1567 <= _16630;
  wire [1:0] _16631 = {_0, _1406} + {_0, _3068};
  wire [1:0] _16632 = {_0, _4640} + {_0, _6814};
  wire [2:0] _16633 = {_0, _16631} + {_0, _16632};
  wire [1:0] _16634 = {_0, _10204} + {_0, _11485};
  wire [3:0] _16635 = {_0, _16633} + {_0, _0, _16634};
  wire _16636 = _12301 < _16635;
  wire _16637 = r1566 ^ _16636;
  wire _16638 = _12298 ? coded_block[1566] : r1566;
  wire _16639 = _12296 ? _16637 : _16638;
  always @ (posedge reset or posedge clock) if (reset) r1566 <= 1'd0; else if (_12300) r1566 <= _16639;
  wire [1:0] _16640 = {_0, _1439} + {_0, _3933};
  wire [1:0] _16641 = {_0, _5152} + {_0, _6718};
  wire [2:0] _16642 = {_0, _16640} + {_0, _16641};
  wire [1:0] _16643 = {_0, _8894} + {_0, _12282};
  wire [3:0] _16644 = {_0, _16642} + {_0, _0, _16643};
  wire _16645 = _12301 < _16644;
  wire _16646 = r1565 ^ _16645;
  wire _16647 = _12298 ? coded_block[1565] : r1565;
  wire _16648 = _12296 ? _16646 : _16647;
  always @ (posedge reset or posedge clock) if (reset) r1565 <= 1'd0; else if (_12300) r1565 <= _16648;
  wire [1:0] _16649 = {_0, _1470} + {_0, _3198};
  wire [1:0] _16650 = {_0, _6012} + {_0, _7230};
  wire [2:0] _16651 = {_0, _16649} + {_0, _16650};
  wire [1:0] _16652 = {_0, _8799} + {_0, _10973};
  wire [3:0] _16653 = {_0, _16651} + {_0, _0, _16652};
  wire _16654 = _12301 < _16653;
  wire _16655 = r1564 ^ _16654;
  wire _16656 = _12298 ? coded_block[1564] : r1564;
  wire _16657 = _12296 ? _16655 : _16656;
  always @ (posedge reset or posedge clock) if (reset) r1564 <= 1'd0; else if (_12300) r1564 <= _16657;
  wire [1:0] _16658 = {_0, _1502} + {_0, _2239};
  wire [1:0] _16659 = {_0, _5279} + {_0, _8092};
  wire [2:0] _16660 = {_0, _16658} + {_0, _16659};
  wire [1:0] _16661 = {_0, _9311} + {_0, _10877};
  wire [3:0] _16662 = {_0, _16660} + {_0, _0, _16661};
  wire _16663 = _12301 < _16662;
  wire _16664 = r1563 ^ _16663;
  wire _16665 = _12298 ? coded_block[1563] : r1563;
  wire _16666 = _12296 ? _16664 : _16665;
  always @ (posedge reset or posedge clock) if (reset) r1563 <= 1'd0; else if (_12300) r1563 <= _16666;
  wire [1:0] _16667 = {_0, _1568} + {_0, _3870};
  wire [1:0] _16668 = {_0, _4861} + {_0, _6397};
  wire [2:0] _16669 = {_0, _16667} + {_0, _16668};
  wire [1:0] _16670 = {_0, _9438} + {_0, _12251};
  wire [3:0] _16671 = {_0, _16669} + {_0, _0, _16670};
  wire _16672 = _12301 < _16671;
  wire _16673 = r1562 ^ _16672;
  wire _16674 = _12298 ? coded_block[1562] : r1562;
  wire _16675 = _12296 ? _16673 : _16674;
  always @ (posedge reset or posedge clock) if (reset) r1562 <= 1'd0; else if (_12300) r1562 <= _16675;
  wire [1:0] _16676 = {_0, _1599} + {_0, _2175};
  wire [1:0] _16677 = {_0, _5949} + {_0, _6942};
  wire [2:0] _16678 = {_0, _16676} + {_0, _16677};
  wire [1:0] _16679 = {_0, _8480} + {_0, _11516};
  wire [3:0] _16680 = {_0, _16678} + {_0, _0, _16679};
  wire _16681 = _12301 < _16680;
  wire _16682 = r1561 ^ _16681;
  wire _16683 = _12298 ? coded_block[1561] : r1561;
  wire _16684 = _12296 ? _16682 : _16683;
  always @ (posedge reset or posedge clock) if (reset) r1561 <= 1'd0; else if (_12300) r1561 <= _16684;
  wire [1:0] _16685 = {_0, _1631} + {_0, _2623};
  wire [1:0] _16686 = {_0, _4256} + {_0, _8028};
  wire [2:0] _16687 = {_0, _16685} + {_0, _16686};
  wire [1:0] _16688 = {_0, _9022} + {_0, _10558};
  wire [3:0] _16689 = {_0, _16687} + {_0, _0, _16688};
  wire _16690 = _12301 < _16689;
  wire _16691 = r1560 ^ _16690;
  wire _16692 = _12298 ? coded_block[1560] : r1560;
  wire _16693 = _12296 ? _16691 : _16692;
  always @ (posedge reset or posedge clock) if (reset) r1560 <= 1'd0; else if (_12300) r1560 <= _16693;
  wire [1:0] _16694 = {_0, _1695} + {_0, _2910};
  wire [1:0] _16695 = {_0, _6076} + {_0, _6781};
  wire [2:0] _16696 = {_0, _16694} + {_0, _16695};
  wire [1:0] _16697 = {_0, _8415} + {_0, _12188};
  wire [3:0] _16698 = {_0, _16696} + {_0, _0, _16697};
  wire _16699 = _12301 < _16698;
  wire _16700 = r1559 ^ _16699;
  wire _16701 = _12298 ? coded_block[1559] : r1559;
  wire _16702 = _12296 ? _16700 : _16701;
  always @ (posedge reset or posedge clock) if (reset) r1559 <= 1'd0; else if (_12300) r1559 <= _16702;
  wire [1:0] _16703 = {_0, _863} + {_0, _3198};
  wire [1:0] _16704 = {_0, _5918} + {_0, _7548};
  wire [2:0] _16705 = {_0, _16703} + {_0, _16704};
  wire [1:0] _16706 = {_0, _9311} + {_0, _10303};
  wire [3:0] _16707 = {_0, _16705} + {_0, _0, _16706};
  wire _16708 = _12301 < _16707;
  wire _16709 = r1558 ^ _16708;
  wire _16710 = _12298 ? coded_block[1558] : r1558;
  wire _16711 = _12296 ? _16709 : _16710;
  always @ (posedge reset or posedge clock) if (reset) r1558 <= 1'd0; else if (_12300) r1558 <= _16711;
  wire [1:0] _16712 = {_0, _894} + {_0, _2112};
  wire [1:0] _16713 = {_0, _5279} + {_0, _7996};
  wire [2:0] _16714 = {_0, _16712} + {_0, _16713};
  wire [1:0] _16715 = {_0, _9630} + {_0, _11389};
  wire [3:0] _16716 = {_0, _16714} + {_0, _0, _16715};
  wire _16717 = _12301 < _16716;
  wire _16718 = r1557 ^ _16717;
  wire _16719 = _12298 ? coded_block[1557] : r1557;
  wire _16720 = _12296 ? _16718 : _16719;
  always @ (posedge reset or posedge clock) if (reset) r1557 <= 1'd0; else if (_12300) r1557 <= _16720;
  wire [1:0] _16721 = {_0, _927} + {_0, _2208};
  wire [1:0] _16722 = {_0, _4192} + {_0, _7357};
  wire [2:0] _16723 = {_0, _16721} + {_0, _16722};
  wire [1:0] _16724 = {_0, _10077} + {_0, _11708};
  wire [3:0] _16725 = {_0, _16723} + {_0, _0, _16724};
  wire _16726 = _12301 < _16725;
  wire _16727 = r1556 ^ _16726;
  wire _16728 = _12298 ? coded_block[1556] : r1556;
  wire _16729 = _12296 ? _16727 : _16728;
  always @ (posedge reset or posedge clock) if (reset) r1556 <= 1'd0; else if (_12300) r1556 <= _16729;
  wire [1:0] _16730 = {_0, _958} + {_0, _3678};
  wire [1:0] _16731 = {_0, _4287} + {_0, _6270};
  wire [2:0] _16732 = {_0, _16730} + {_0, _16731};
  wire [1:0] _16733 = {_0, _9438} + {_0, _12155};
  wire [3:0] _16734 = {_0, _16732} + {_0, _0, _16733};
  wire _16735 = _12301 < _16734;
  wire _16736 = r1555 ^ _16735;
  wire _16737 = _12298 ? coded_block[1555] : r1555;
  wire _16738 = _12296 ? _16736 : _16737;
  always @ (posedge reset or posedge clock) if (reset) r1555 <= 1'd0; else if (_12300) r1555 <= _16738;
  wire [1:0] _16739 = {_0, _1021} + {_0, _2813};
  wire [1:0] _16740 = {_0, _6012} + {_0, _7837};
  wire [2:0] _16741 = {_0, _16739} + {_0, _16740};
  wire [1:0] _16742 = {_0, _8446} + {_0, _10430};
  wire [3:0] _16743 = {_0, _16741} + {_0, _0, _16742};
  wire _16744 = _12301 < _16743;
  wire _16745 = r1554 ^ _16744;
  wire _16746 = _12298 ? coded_block[1554] : r1554;
  wire _16747 = _12296 ? _16745 : _16746;
  always @ (posedge reset or posedge clock) if (reset) r1554 <= 1'd0; else if (_12300) r1554 <= _16747;
  wire [1:0] _16748 = {_0, _1375} + {_0, _3325};
  wire [1:0] _16749 = {_0, _4926} + {_0, _6589};
  wire [2:0] _16750 = {_0, _16748} + {_0, _16749};
  wire [1:0] _16751 = {_0, _9661} + {_0, _12124};
  wire [3:0] _16752 = {_0, _16750} + {_0, _0, _16751};
  wire _16753 = _12301 < _16752;
  wire _16754 = r1553 ^ _16753;
  wire _16755 = _12298 ? coded_block[1553] : r1553;
  wire _16756 = _12296 ? _16754 : _16755;
  always @ (posedge reset or posedge clock) if (reset) r1553 <= 1'd0; else if (_12300) r1553 <= _16756;
  wire [1:0] _16757 = {_0, _34} + {_0, _3068};
  wire [1:0] _16758 = {_0, _5152} + {_0, _7230};
  wire [2:0] _16759 = {_0, _16757} + {_0, _16758};
  wire [1:0] _16760 = {_0, _9311} + {_0, _11389};
  wire [3:0] _16761 = {_0, _16759} + {_0, _0, _16760};
  wire _16762 = _12301 < _16761;
  wire _16763 = r1552 ^ _16762;
  wire _16764 = _12298 ? coded_block[1552] : r1552;
  wire _16765 = _12296 ? _16763 : _16764;
  always @ (posedge reset or posedge clock) if (reset) r1552 <= 1'd0; else if (_12300) r1552 <= _16765;
  wire [1:0] _16766 = {_0, _2044} + {_0, _3167};
  wire [1:0] _16767 = {_0, _4223} + {_0, _6687};
  wire [2:0] _16768 = {_0, _16766} + {_0, _16767};
  wire [1:0] _16769 = {_0, _9212} + {_0, _10685};
  wire [3:0] _16770 = {_0, _16768} + {_0, _0, _16769};
  wire _16771 = _12301 < _16770;
  wire _16772 = r1551 ^ _16771;
  wire _16773 = _12298 ? coded_block[1551] : r1551;
  wire _16774 = _12296 ? _16772 : _16773;
  always @ (posedge reset or posedge clock) if (reset) r1551 <= 1'd0; else if (_12300) r1551 <= _16774;
  wire [1:0] _16775 = {_0, _65} + {_0, _3580};
  wire [1:0] _16776 = {_0, _5246} + {_0, _6303};
  wire [2:0] _16777 = {_0, _16775} + {_0, _16776};
  wire [1:0] _16778 = {_0, _8767} + {_0, _11295};
  wire [3:0] _16779 = {_0, _16777} + {_0, _0, _16778};
  wire _16780 = _12301 < _16779;
  wire _16781 = r1550 ^ _16780;
  wire _16782 = _12298 ? coded_block[1550] : r1550;
  wire _16783 = _12296 ? _16781 : _16782;
  always @ (posedge reset or posedge clock) if (reset) r1550 <= 1'd0; else if (_12300) r1550 <= _16783;
  wire [1:0] _16784 = {_0, _97} + {_0, _4060};
  wire [1:0] _16785 = {_0, _5663} + {_0, _7326};
  wire [2:0] _16786 = {_0, _16784} + {_0, _16785};
  wire [1:0] _16787 = {_0, _8383} + {_0, _10846};
  wire [3:0] _16788 = {_0, _16786} + {_0, _0, _16787};
  wire _16789 = _12301 < _16788;
  wire _16790 = r1549 ^ _16789;
  wire _16791 = _12298 ? coded_block[1549] : r1549;
  wire _16792 = _12296 ? _16790 : _16791;
  always @ (posedge reset or posedge clock) if (reset) r1549 <= 1'd0; else if (_12300) r1549 <= _16792;
  wire [1:0] _16793 = {_0, _128} + {_0, _3486};
  wire [1:0] _16794 = {_0, _6139} + {_0, _7741};
  wire [2:0] _16795 = {_0, _16793} + {_0, _16794};
  wire [1:0] _16796 = {_0, _9406} + {_0, _10462};
  wire [3:0] _16797 = {_0, _16795} + {_0, _0, _16796};
  wire _16798 = _12301 < _16797;
  wire _16799 = r1548 ^ _16798;
  wire _16800 = _12298 ? coded_block[1548] : r1548;
  wire _16801 = _12296 ? _16799 : _16800;
  always @ (posedge reset or posedge clock) if (reset) r1548 <= 1'd0; else if (_12300) r1548 <= _16801;
  wire [1:0] _16802 = {_0, _192} + {_0, _2463};
  wire [1:0] _16803 = {_0, _4861} + {_0, _7644};
  wire [2:0] _16804 = {_0, _16802} + {_0, _16803};
  wire [1:0] _16805 = {_0, _8288} + {_0, _11900};
  wire [3:0] _16806 = {_0, _16804} + {_0, _0, _16805};
  wire _16807 = _12301 < _16806;
  wire _16808 = r1547 ^ _16807;
  wire _16809 = _12298 ? coded_block[1547] : r1547;
  wire _16810 = _12296 ? _16808 : _16809;
  always @ (posedge reset or posedge clock) if (reset) r1547 <= 1'd0; else if (_12300) r1547 <= _16810;
  wire [1:0] _16811 = {_0, _224} + {_0, _2623};
  wire [1:0] _16812 = {_0, _4542} + {_0, _6942};
  wire [2:0] _16813 = {_0, _16811} + {_0, _16812};
  wire [1:0] _16814 = {_0, _9724} + {_0, _10366};
  wire [3:0] _16815 = {_0, _16813} + {_0, _0, _16814};
  wire _16816 = _12301 < _16815;
  wire _16817 = r1546 ^ _16816;
  wire _16818 = _12298 ? coded_block[1546] : r1546;
  wire _16819 = _12296 ? _16817 : _16818;
  always @ (posedge reset or posedge clock) if (reset) r1546 <= 1'd0; else if (_12300) r1546 <= _16819;
  wire [1:0] _16820 = {_0, _255} + {_0, _2430};
  wire [1:0] _16821 = {_0, _4703} + {_0, _6621};
  wire [2:0] _16822 = {_0, _16820} + {_0, _16821};
  wire [1:0] _16823 = {_0, _9022} + {_0, _11806};
  wire [3:0] _16824 = {_0, _16822} + {_0, _0, _16823};
  wire _16825 = _12301 < _16824;
  wire _16826 = r1545 ^ _16825;
  wire _16827 = _12298 ? coded_block[1545] : r1545;
  wire _16828 = _12296 ? _16826 : _16827;
  always @ (posedge reset or posedge clock) if (reset) r1545 <= 1'd0; else if (_12300) r1545 <= _16828;
  wire [1:0] _16829 = {_0, _289} + {_0, _2813};
  wire [1:0] _16830 = {_0, _4511} + {_0, _6781};
  wire [2:0] _16831 = {_0, _16829} + {_0, _16830};
  wire [1:0] _16832 = {_0, _8701} + {_0, _11101};
  wire [3:0] _16833 = {_0, _16831} + {_0, _0, _16832};
  wire _16834 = _12301 < _16833;
  wire _16835 = r1544 ^ _16834;
  wire _16836 = _12298 ? coded_block[1544] : r1544;
  wire _16837 = _12296 ? _16835 : _16836;
  always @ (posedge reset or posedge clock) if (reset) r1544 <= 1'd0; else if (_12300) r1544 <= _16837;
  wire [1:0] _16838 = {_0, _320} + {_0, _3964};
  wire [1:0] _16839 = {_0, _4895} + {_0, _6589};
  wire [2:0] _16840 = {_0, _16838} + {_0, _16839};
  wire [1:0] _16841 = {_0, _8863} + {_0, _10783};
  wire [3:0] _16842 = {_0, _16840} + {_0, _0, _16841};
  wire _16843 = _12301 < _16842;
  wire _16844 = r1543 ^ _16843;
  wire _16845 = _12298 ? coded_block[1543] : r1543;
  wire _16846 = _12296 ? _16844 : _16845;
  always @ (posedge reset or posedge clock) if (reset) r1543 <= 1'd0; else if (_12300) r1543 <= _16846;
  wire [1:0] _16847 = {_0, _352} + {_0, _3742};
  wire [1:0] _16848 = {_0, _6045} + {_0, _6973};
  wire [2:0] _16849 = {_0, _16847} + {_0, _16848};
  wire [1:0] _16850 = {_0, _8670} + {_0, _10941};
  wire [3:0] _16851 = {_0, _16849} + {_0, _0, _16850};
  wire _16852 = _12301 < _16851;
  wire _16853 = r1542 ^ _16852;
  wire _16854 = _12298 ? coded_block[1542] : r1542;
  wire _16855 = _12296 ? _16853 : _16854;
  always @ (posedge reset or posedge clock) if (reset) r1542 <= 1'd0; else if (_12300) r1542 <= _16855;
  wire [1:0] _16856 = {_0, _383} + {_0, _2302};
  wire [1:0] _16857 = {_0, _5821} + {_0, _8123};
  wire [2:0] _16858 = {_0, _16856} + {_0, _16857};
  wire [1:0] _16859 = {_0, _9054} + {_0, _10748};
  wire [3:0] _16860 = {_0, _16858} + {_0, _0, _16859};
  wire _16861 = _12301 < _16860;
  wire _16862 = r1541 ^ _16861;
  wire _16863 = _12298 ? coded_block[1541] : r1541;
  wire _16864 = _12296 ? _16862 : _16863;
  always @ (posedge reset or posedge clock) if (reset) r1541 <= 1'd0; else if (_12300) r1541 <= _16864;
  wire [1:0] _16865 = {_0, _416} + {_0, _2239};
  wire [1:0] _16866 = {_0, _4384} + {_0, _7900};
  wire [2:0] _16867 = {_0, _16865} + {_0, _16866};
  wire [1:0] _16868 = {_0, _10204} + {_0, _11132};
  wire [3:0] _16869 = {_0, _16867} + {_0, _0, _16868};
  wire _16870 = _12301 < _16869;
  wire _16871 = r1540 ^ _16870;
  wire _16872 = _12298 ? coded_block[1540] : r1540;
  wire _16873 = _12296 ? _16871 : _16872;
  always @ (posedge reset or posedge clock) if (reset) r1540 <= 1'd0; else if (_12300) r1540 <= _16873;
  wire [1:0] _16874 = {_0, _479} + {_0, _4028};
  wire [1:0] _16875 = {_0, _5438} + {_0, _6397};
  wire [2:0] _16876 = {_0, _16874} + {_0, _16875};
  wire [1:0] _16877 = {_0, _8543} + {_0, _12061};
  wire [3:0] _16878 = {_0, _16876} + {_0, _0, _16877};
  wire _16879 = _12301 < _16878;
  wire _16880 = r1539 ^ _16879;
  wire _16881 = _12298 ? coded_block[1539] : r1539;
  wire _16882 = _12296 ? _16880 : _16881;
  always @ (posedge reset or posedge clock) if (reset) r1539 <= 1'd0; else if (_12300) r1539 <= _16882;
  wire [1:0] _16883 = {_0, _545} + {_0, _3325};
  wire [1:0] _16884 = {_0, _5694} + {_0, _8186};
  wire [2:0] _16885 = {_0, _16883} + {_0, _16884};
  wire [1:0] _16886 = {_0, _9597} + {_0, _10558};
  wire [3:0] _16887 = {_0, _16885} + {_0, _0, _16886};
  wire _16888 = _12301 < _16887;
  wire _16889 = r1538 ^ _16888;
  wire _16890 = _12298 ? coded_block[1538] : r1538;
  wire _16891 = _12296 ? _16889 : _16890;
  always @ (posedge reset or posedge clock) if (reset) r1538 <= 1'd0; else if (_12300) r1538 <= _16891;
  wire [1:0] _16892 = {_0, _608} + {_0, _3773};
  wire [1:0] _16893 = {_0, _4350} + {_0, _7485};
  wire [2:0] _16894 = {_0, _16892} + {_0, _16893};
  wire [1:0] _16895 = {_0, _9853} + {_0, _10335};
  wire [3:0] _16896 = {_0, _16894} + {_0, _0, _16895};
  wire _16897 = _12301 < _16896;
  wire _16898 = r1537 ^ _16897;
  wire _16899 = _12298 ? coded_block[1537] : r1537;
  wire _16900 = _12296 ? _16898 : _16899;
  always @ (posedge reset or posedge clock) if (reset) r1537 <= 1'd0; else if (_12300) r1537 <= _16900;
  wire [1:0] _16901 = {_0, _34} + {_0, _3580};
  wire [1:0] _16902 = {_0, _5663} + {_0, _7741};
  wire [2:0] _16903 = {_0, _16901} + {_0, _16902};
  wire [1:0] _16904 = {_0, _9822} + {_0, _11900};
  wire [3:0] _16905 = {_0, _16903} + {_0, _0, _16904};
  wire _16906 = _12301 < _16905;
  wire _16907 = r1536 ^ _16906;
  wire _16908 = _12298 ? coded_block[1536] : r1536;
  wire _16909 = _12296 ? _16907 : _16908;
  always @ (posedge reset or posedge clock) if (reset) r1536 <= 1'd0; else if (_12300) r1536 <= _16909;
  wire [1:0] _16910 = {_0, _65} + {_0, _3068};
  wire [1:0] _16911 = {_0, _4703} + {_0, _6462};
  wire [2:0] _16912 = {_0, _16910} + {_0, _16911};
  wire [1:0] _16913 = {_0, _9469} + {_0, _11004};
  wire [3:0] _16914 = {_0, _16912} + {_0, _0, _16913};
  wire _16915 = _12301 < _16914;
  wire _16916 = r1535 ^ _16915;
  wire _16917 = _12298 ? coded_block[1535] : r1535;
  wire _16918 = _12296 ? _16916 : _16917;
  always @ (posedge reset or posedge clock) if (reset) r1535 <= 1'd0; else if (_12300) r1535 <= _16918;
  wire [1:0] _16919 = {_0, _97} + {_0, _2430};
  wire [1:0] _16920 = {_0, _5152} + {_0, _6781};
  wire [2:0] _16921 = {_0, _16919} + {_0, _16920};
  wire [1:0] _16922 = {_0, _8543} + {_0, _11550};
  wire [3:0] _16923 = {_0, _16921} + {_0, _0, _16922};
  wire _16924 = _12301 < _16923;
  wire _16925 = r1534 ^ _16924;
  wire _16926 = _12298 ? coded_block[1534] : r1534;
  wire _16927 = _12296 ? _16925 : _16926;
  always @ (posedge reset or posedge clock) if (reset) r1534 <= 1'd0; else if (_12300) r1534 <= _16927;
  wire [1:0] _16928 = {_0, _128} + {_0, _3359};
  wire [1:0] _16929 = {_0, _4511} + {_0, _7230};
  wire [2:0] _16930 = {_0, _16928} + {_0, _16929};
  wire [1:0] _16931 = {_0, _8863} + {_0, _10621};
  wire [3:0] _16932 = {_0, _16930} + {_0, _0, _16931};
  wire _16933 = _12301 < _16932;
  wire _16934 = r1533 ^ _16933;
  wire _16935 = _12298 ? coded_block[1533] : r1533;
  wire _16936 = _12296 ? _16934 : _16935;
  always @ (posedge reset or posedge clock) if (reset) r1533 <= 1'd0; else if (_12300) r1533 <= _16936;
  wire [1:0] _16937 = {_0, _34} + {_0, _2271};
  wire [1:0] _16938 = {_0, _4350} + {_0, _6431};
  wire [2:0] _16939 = {_0, _16937} + {_0, _16938};
  wire [1:0] _16940 = {_0, _8511} + {_0, _10590};
  wire [3:0] _16941 = {_0, _16939} + {_0, _0, _16940};
  wire _16942 = _12301 < _16941;
  wire _16943 = r1532 ^ _16942;
  wire _16944 = _12298 ? coded_block[1532] : r1532;
  wire _16945 = _12296 ? _16943 : _16944;
  always @ (posedge reset or posedge clock) if (reset) r1532 <= 1'd0; else if (_12300) r1532 <= _16945;
  wire [1:0] _16946 = {_0, _479} + {_0, _3805};
  wire [1:0] _16947 = {_0, _5183} + {_0, _6462};
  wire [2:0] _16948 = {_0, _16946} + {_0, _16947};
  wire [1:0] _16949 = {_0, _8480} + {_0, _11358};
  wire [3:0] _16950 = {_0, _16948} + {_0, _0, _16949};
  wire _16951 = _12301 < _16950;
  wire _16952 = r1531 ^ _16951;
  wire _16953 = _12298 ? coded_block[1531] : r1531;
  wire _16954 = _12296 ? _16952 : _16953;
  always @ (posedge reset or posedge clock) if (reset) r1531 <= 1'd0; else if (_12300) r1531 <= _16954;
  wire [1:0] _16955 = {_0, _510} + {_0, _3709};
  wire [1:0] _16956 = {_0, _5884} + {_0, _7262};
  wire [2:0] _16957 = {_0, _16955} + {_0, _16956};
  wire [1:0] _16958 = {_0, _8543} + {_0, _10558};
  wire [3:0] _16959 = {_0, _16957} + {_0, _0, _16958};
  wire _16960 = _12301 < _16959;
  wire _16961 = r1530 ^ _16960;
  wire _16962 = _12298 ? coded_block[1530] : r1530;
  wire _16963 = _12296 ? _16961 : _16962;
  always @ (posedge reset or posedge clock) if (reset) r1530 <= 1'd0; else if (_12300) r1530 <= _16963;
  wire [1:0] _16964 = {_0, _545} + {_0, _2208};
  wire [1:0] _16965 = {_0, _5790} + {_0, _7965};
  wire [2:0] _16966 = {_0, _16964} + {_0, _16965};
  wire [1:0] _16967 = {_0, _9342} + {_0, _10621};
  wire [3:0] _16968 = {_0, _16966} + {_0, _0, _16967};
  wire _16969 = _12301 < _16968;
  wire _16970 = r1529 ^ _16969;
  wire _16971 = _12298 ? coded_block[1529] : r1529;
  wire _16972 = _12296 ? _16970 : _16971;
  always @ (posedge reset or posedge clock) if (reset) r1529 <= 1'd0; else if (_12300) r1529 <= _16972;
  wire [1:0] _16973 = {_0, _576} + {_0, _3068};
  wire [1:0] _16974 = {_0, _4287} + {_0, _7868};
  wire [2:0] _16975 = {_0, _16973} + {_0, _16974};
  wire [1:0] _16976 = {_0, _10045} + {_0, _11422};
  wire [3:0] _16977 = {_0, _16975} + {_0, _0, _16976};
  wire _16978 = _12301 < _16977;
  wire _16979 = r1528 ^ _16978;
  wire _16980 = _12298 ? coded_block[1528] : r1528;
  wire _16981 = _12296 ? _16979 : _16980;
  always @ (posedge reset or posedge clock) if (reset) r1528 <= 1'd0; else if (_12300) r1528 <= _16981;
  wire [1:0] _16982 = {_0, _608} + {_0, _2336};
  wire [1:0] _16983 = {_0, _5152} + {_0, _6366};
  wire [2:0] _16984 = {_0, _16982} + {_0, _16983};
  wire [1:0] _16985 = {_0, _9949} + {_0, _12124};
  wire [3:0] _16986 = {_0, _16984} + {_0, _0, _16985};
  wire _16987 = _12301 < _16986;
  wire _16988 = r1527 ^ _16987;
  wire _16989 = _12298 ? coded_block[1527] : r1527;
  wire _16990 = _12296 ? _16988 : _16989;
  always @ (posedge reset or posedge clock) if (reset) r1527 <= 1'd0; else if (_12300) r1527 <= _16990;
  wire [1:0] _16991 = {_0, _639} + {_0, _3390};
  wire [1:0] _16992 = {_0, _4415} + {_0, _7230};
  wire [2:0] _16993 = {_0, _16991} + {_0, _16992};
  wire [1:0] _16994 = {_0, _8446} + {_0, _12027};
  wire [3:0] _16995 = {_0, _16993} + {_0, _0, _16994};
  wire _16996 = _12301 < _16995;
  wire _16997 = r1526 ^ _16996;
  wire _16998 = _12298 ? coded_block[1526] : r1526;
  wire _16999 = _12296 ? _16997 : _16998;
  always @ (posedge reset or posedge clock) if (reset) r1526 <= 1'd0; else if (_12300) r1526 <= _16999;
  wire [1:0] _17000 = {_0, _34} + {_0, _3262};
  wire [1:0] _17001 = {_0, _5342} + {_0, _7420};
  wire [2:0] _17002 = {_0, _17000} + {_0, _17001};
  wire [1:0] _17003 = {_0, _9503} + {_0, _11581};
  wire [3:0] _17004 = {_0, _17002} + {_0, _0, _17003};
  wire _17005 = _12301 < _17004;
  wire _17006 = r1525 ^ _17005;
  wire _17007 = _12298 ? coded_block[1525] : r1525;
  wire _17008 = _12296 ? _17006 : _17007;
  always @ (posedge reset or posedge clock) if (reset) r1525 <= 1'd0; else if (_12300) r1525 <= _17008;
  wire [1:0] _17009 = {_0, _2013} + {_0, _3615};
  wire [1:0] _17010 = {_0, _5470} + {_0, _7900};
  wire [2:0] _17011 = {_0, _17009} + {_0, _17010};
  wire [1:0] _17012 = {_0, _9085} + {_0, _10910};
  wire [3:0] _17013 = {_0, _17011} + {_0, _0, _17012};
  wire _17014 = _12301 < _17013;
  wire _17015 = r1524 ^ _17014;
  wire _17016 = _12298 ? coded_block[1524] : r1524;
  wire _17017 = _12296 ? _17015 : _17016;
  always @ (posedge reset or posedge clock) if (reset) r1524 <= 1'd0; else if (_12300) r1524 <= _17017;
  wire [1:0] _17018 = {_0, _2044} + {_0, _3486};
  wire [1:0] _17019 = {_0, _5694} + {_0, _7548};
  wire [2:0] _17020 = {_0, _17018} + {_0, _17019};
  wire [1:0] _17021 = {_0, _9980} + {_0, _11165};
  wire [3:0] _17022 = {_0, _17020} + {_0, _0, _17021};
  wire _17023 = _12301 < _17022;
  wire _17024 = r1523 ^ _17023;
  wire _17025 = _12298 ? coded_block[1523] : r1523;
  wire _17026 = _12296 ? _17024 : _17025;
  always @ (posedge reset or posedge clock) if (reset) r1523 <= 1'd0; else if (_12300) r1523 <= _17026;
  wire [1:0] _17027 = {_0, _65} + {_0, _3836};
  wire [1:0] _17028 = {_0, _5565} + {_0, _7773};
  wire [2:0] _17029 = {_0, _17027} + {_0, _17028};
  wire [1:0] _17030 = {_0, _9630} + {_0, _12061};
  wire [3:0] _17031 = {_0, _17029} + {_0, _0, _17030};
  wire _17032 = _12301 < _17031;
  wire _17033 = r1522 ^ _17032;
  wire _17034 = _12298 ? coded_block[1522] : r1522;
  wire _17035 = _12296 ? _17033 : _17034;
  always @ (posedge reset or posedge clock) if (reset) r1522 <= 1'd0; else if (_12300) r1522 <= _17035;
  wire [1:0] _17036 = {_0, _97} + {_0, _2557};
  wire [1:0] _17037 = {_0, _5918} + {_0, _7644};
  wire [2:0] _17038 = {_0, _17036} + {_0, _17037};
  wire [1:0] _17039 = {_0, _9853} + {_0, _11708};
  wire [3:0] _17040 = {_0, _17038} + {_0, _0, _17039};
  wire _17041 = _12301 < _17040;
  wire _17042 = r1521 ^ _17041;
  wire _17043 = _12298 ? coded_block[1521] : r1521;
  wire _17044 = _12296 ? _17042 : _17043;
  always @ (posedge reset or posedge clock) if (reset) r1521 <= 1'd0; else if (_12300) r1521 <= _17044;
  wire [1:0] _17045 = {_0, _128} + {_0, _3167};
  wire [1:0] _17046 = {_0, _4640} + {_0, _7996};
  wire [2:0] _17047 = {_0, _17045} + {_0, _17046};
  wire [1:0] _17048 = {_0, _9724} + {_0, _11933};
  wire [3:0] _17049 = {_0, _17047} + {_0, _0, _17048};
  wire _17050 = _12301 < _17049;
  wire _17051 = r1520 ^ _17050;
  wire _17052 = _12298 ? coded_block[1520] : r1520;
  wire _17053 = _12296 ? _17051 : _17052;
  always @ (posedge reset or posedge clock) if (reset) r1520 <= 1'd0; else if (_12300) r1520 <= _17053;
  wire [1:0] _17054 = {_0, _34} + {_0, _3231};
  wire [1:0] _17055 = {_0, _5310} + {_0, _7389};
  wire [2:0] _17056 = {_0, _17054} + {_0, _17055};
  wire [1:0] _17057 = {_0, _9469} + {_0, _11550};
  wire [3:0] _17058 = {_0, _17056} + {_0, _0, _17057};
  wire _17059 = _12301 < _17058;
  wire _17060 = r1519 ^ _17059;
  wire _17061 = _12298 ? coded_block[1519] : r1519;
  wire _17062 = _12296 ? _17060 : _17061;
  always @ (posedge reset or posedge clock) if (reset) r1519 <= 1'd0; else if (_12300) r1519 <= _17062;
  wire [1:0] _17063 = {_0, _1247} + {_0, _3615};
  wire [1:0] _17064 = {_0, _5501} + {_0, _6176};
  wire [2:0] _17065 = {_0, _17063} + {_0, _17064};
  wire [1:0] _17066 = {_0, _9630} + {_0, _11869};
  wire [3:0] _17067 = {_0, _17065} + {_0, _0, _17066};
  wire _17068 = _12301 < _17067;
  wire _17069 = r1518 ^ _17068;
  wire _17070 = _12298 ? coded_block[1518] : r1518;
  wire _17071 = _12296 ? _17069 : _17070;
  always @ (posedge reset or posedge clock) if (reset) r1518 <= 1'd0; else if (_12300) r1518 <= _17071;
  wire [1:0] _17072 = {_0, _1278} + {_0, _2239};
  wire [1:0] _17073 = {_0, _5694} + {_0, _7581};
  wire [2:0] _17074 = {_0, _17072} + {_0, _17073};
  wire [1:0] _17075 = {_0, _8225} + {_0, _11708};
  wire [3:0] _17076 = {_0, _17074} + {_0, _0, _17075};
  wire _17077 = _12301 < _17076;
  wire _17078 = r1517 ^ _17077;
  wire _17079 = _12298 ? coded_block[1517] : r1517;
  wire _17080 = _12296 ? _17078 : _17079;
  always @ (posedge reset or posedge clock) if (reset) r1517 <= 1'd0; else if (_12300) r1517 <= _17080;
  wire [1:0] _17081 = {_0, _1375} + {_0, _3262};
  wire [1:0] _17082 = {_0, _5279} + {_0, _8155};
  wire [2:0] _17083 = {_0, _17081} + {_0, _17082};
  wire [1:0] _17084 = {_0, _8480} + {_0, _11933};
  wire [3:0] _17085 = {_0, _17083} + {_0, _0, _17084};
  wire _17086 = _12301 < _17085;
  wire _17087 = r1516 ^ _17086;
  wire _17088 = _12298 ? coded_block[1516] : r1516;
  wire _17089 = _12296 ? _17087 : _17088;
  always @ (posedge reset or posedge clock) if (reset) r1516 <= 1'd0; else if (_12300) r1516 <= _17089;
  wire [1:0] _17090 = {_0, _1406} + {_0, _4060};
  wire [1:0] _17091 = {_0, _5342} + {_0, _7357};
  wire [2:0] _17092 = {_0, _17090} + {_0, _17091};
  wire [1:0] _17093 = {_0, _10235} + {_0, _10558};
  wire [3:0] _17094 = {_0, _17092} + {_0, _0, _17093};
  wire _17095 = _12301 < _17094;
  wire _17096 = r1515 ^ _17095;
  wire _17097 = _12298 ? coded_block[1515] : r1515;
  wire _17098 = _12296 ? _17096 : _17097;
  always @ (posedge reset or posedge clock) if (reset) r1515 <= 1'd0; else if (_12300) r1515 <= _17098;
  wire [1:0] _17099 = {_0, _34} + {_0, _3422};
  wire [1:0] _17100 = {_0, _5501} + {_0, _7581};
  wire [2:0] _17101 = {_0, _17099} + {_0, _17100};
  wire [1:0] _17102 = {_0, _9661} + {_0, _11740};
  wire [3:0] _17103 = {_0, _17101} + {_0, _0, _17102};
  wire _17104 = _12301 < _17103;
  wire _17105 = r1514 ^ _17104;
  wire _17106 = _12298 ? coded_block[1514] : r1514;
  wire _17107 = _12296 ? _17105 : _17106;
  always @ (posedge reset or posedge clock) if (reset) r1514 <= 1'd0; else if (_12300) r1514 <= _17107;
  wire [1:0] _17108 = {_0, _990} + {_0, _3104};
  wire [1:0] _17109 = {_0, _4192} + {_0, _6781};
  wire [2:0] _17110 = {_0, _17108} + {_0, _17109};
  wire [1:0] _17111 = {_0, _9917} + {_0, _12282};
  wire [3:0] _17112 = {_0, _17110} + {_0, _0, _17111};
  wire _17113 = _12301 < _17112;
  wire _17114 = r1513 ^ _17113;
  wire _17115 = _12298 ? coded_block[1513] : r1513;
  wire _17116 = _12296 ? _17114 : _17115;
  always @ (posedge reset or posedge clock) if (reset) r1513 <= 1'd0; else if (_12300) r1513 <= _17116;
  wire [1:0] _17117 = {_0, _1088} + {_0, _2557};
  wire [1:0] _17118 = {_0, _5116} + {_0, _8028};
  wire [2:0] _17119 = {_0, _17117} + {_0, _17118};
  wire [1:0] _17120 = {_0, _9342} + {_0, _10430};
  wire [3:0] _17121 = {_0, _17119} + {_0, _0, _17120};
  wire _17122 = _12301 < _17121;
  wire _17123 = r1512 ^ _17122;
  wire _17124 = _12298 ? coded_block[1512] : r1512;
  wire _17125 = _12296 ? _17123 : _17124;
  always @ (posedge reset or posedge clock) if (reset) r1512 <= 1'd0; else if (_12300) r1512 <= _17125;
  wire [1:0] _17126 = {_0, _1120} + {_0, _2686};
  wire [1:0] _17127 = {_0, _4640} + {_0, _7199};
  wire [2:0] _17128 = {_0, _17126} + {_0, _17127};
  wire [1:0] _17129 = {_0, _10108} + {_0, _11422};
  wire [3:0] _17130 = {_0, _17128} + {_0, _0, _17129};
  wire _17131 = _12301 < _17130;
  wire _17132 = r1511 ^ _17131;
  wire _17133 = _12298 ? coded_block[1511] : r1511;
  wire _17134 = _12296 ? _17132 : _17133;
  always @ (posedge reset or posedge clock) if (reset) r1511 <= 1'd0; else if (_12300) r1511 <= _17134;
  wire [1:0] _17135 = {_0, _1151} + {_0, _4028};
  wire [1:0] _17136 = {_0, _4767} + {_0, _6718};
  wire [2:0] _17137 = {_0, _17135} + {_0, _17136};
  wire [1:0] _17138 = {_0, _9279} + {_0, _12188};
  wire [3:0] _17139 = {_0, _17137} + {_0, _0, _17138};
  wire _17140 = _12301 < _17139;
  wire _17141 = r1510 ^ _17140;
  wire _17142 = _12298 ? coded_block[1510] : r1510;
  wire _17143 = _12296 ? _17141 : _17142;
  always @ (posedge reset or posedge clock) if (reset) r1510 <= 1'd0; else if (_12300) r1510 <= _17143;
  wire [1:0] _17144 = {_0, _34} + {_0, _2208};
  wire [1:0] _17145 = {_0, _4287} + {_0, _6366};
  wire [2:0] _17146 = {_0, _17144} + {_0, _17145};
  wire [1:0] _17147 = {_0, _8446} + {_0, _10527};
  wire [3:0] _17148 = {_0, _17146} + {_0, _0, _17147};
  wire _17149 = _12301 < _17148;
  wire _17150 = r1509 ^ _17149;
  wire _17151 = _12298 ? coded_block[1509] : r1509;
  wire _17152 = _12296 ? _17150 : _17151;
  always @ (posedge reset or posedge clock) if (reset) r1509 <= 1'd0; else if (_12300) r1509 <= _17152;
  wire [1:0] _17153 = {_0, _672} + {_0, _3262};
  wire [1:0] _17154 = {_0, _5022} + {_0, _8028};
  wire [2:0] _17155 = {_0, _17153} + {_0, _17154};
  wire [1:0] _17156 = {_0, _9566} + {_0, _10590};
  wire [3:0] _17157 = {_0, _17155} + {_0, _0, _17156};
  wire _17158 = _12301 < _17157;
  wire _17159 = r1508 ^ _17158;
  wire _17160 = _12298 ? coded_block[1508] : r1508;
  wire _17161 = _12296 ? _17159 : _17160;
  always @ (posedge reset or posedge clock) if (reset) r1508 <= 1'd0; else if (_12300) r1508 <= _17161;
  wire [1:0] _17162 = {_0, _735} + {_0, _3068};
  wire [1:0] _17163 = {_0, _5790} + {_0, _7420};
  wire [2:0] _17164 = {_0, _17162} + {_0, _17163};
  wire [1:0] _17165 = {_0, _9181} + {_0, _12188};
  wire [3:0] _17166 = {_0, _17164} + {_0, _0, _17165};
  wire _17167 = _12301 < _17166;
  wire _17168 = r1507 ^ _17167;
  wire _17169 = _12298 ? coded_block[1507] : r1507;
  wire _17170 = _12296 ? _17168 : _17169;
  always @ (posedge reset or posedge clock) if (reset) r1507 <= 1'd0; else if (_12300) r1507 <= _17170;
  wire [1:0] _17171 = {_0, _800} + {_0, _4091};
  wire [1:0] _17172 = {_0, _6076} + {_0, _7230};
  wire [2:0] _17173 = {_0, _17171} + {_0, _17172};
  wire [1:0] _17174 = {_0, _9949} + {_0, _11581};
  wire [3:0] _17175 = {_0, _17173} + {_0, _0, _17174};
  wire _17176 = _12301 < _17175;
  wire _17177 = r1506 ^ _17176;
  wire _17178 = _12298 ? coded_block[1506] : r1506;
  wire _17179 = _12296 ? _17177 : _17178;
  always @ (posedge reset or posedge clock) if (reset) r1506 <= 1'd0; else if (_12300) r1506 <= _17179;
  wire [1:0] _17180 = {_0, _34} + {_0, _3549};
  wire [1:0] _17181 = {_0, _5628} + {_0, _7710};
  wire [2:0] _17182 = {_0, _17180} + {_0, _17181};
  wire [1:0] _17183 = {_0, _9790} + {_0, _11869};
  wire [3:0] _17184 = {_0, _17182} + {_0, _0, _17183};
  wire _17185 = _12301 < _17184;
  wire _17186 = r1505 ^ _17185;
  wire _17187 = _12298 ? coded_block[1505] : r1505;
  wire _17188 = _12296 ? _17186 : _17187;
  always @ (posedge reset or posedge clock) if (reset) r1505 <= 1'd0; else if (_12300) r1505 <= _17188;
  wire [1:0] _17189 = {_0, _831} + {_0, _2208};
  wire [1:0] _17190 = {_0, _4511} + {_0, _7454};
  wire [2:0] _17191 = {_0, _17189} + {_0, _17190};
  wire [1:0] _17192 = {_0, _9149} + {_0, _11422};
  wire [3:0] _17193 = {_0, _17191} + {_0, _0, _17192};
  wire _17194 = _12301 < _17193;
  wire _17195 = r1504 ^ _17194;
  wire _17196 = _12298 ? coded_block[1504] : r1504;
  wire _17197 = _12296 ? _17195 : _17196;
  always @ (posedge reset or posedge clock) if (reset) r1504 <= 1'd0; else if (_12300) r1504 <= _17197;
  wire [1:0] _17198 = {_0, _34} + {_0, _3646};
  wire [1:0] _17199 = {_0, _5726} + {_0, _7804};
  wire [2:0] _17200 = {_0, _17198} + {_0, _17199};
  wire [1:0] _17201 = {_0, _9886} + {_0, _11964};
  wire [3:0] _17202 = {_0, _17200} + {_0, _0, _17201};
  wire _17203 = _12301 < _17202;
  wire _17204 = r1503 ^ _17203;
  wire _17205 = _12298 ? coded_block[1503] : r1503;
  wire _17206 = _12296 ? _17204 : _17205;
  always @ (posedge reset or posedge clock) if (reset) r1503 <= 1'd0; else if (_12300) r1503 <= _17206;
  wire [1:0] _17207 = {_0, _34} + {_0, _3294};
  wire [1:0] _17208 = {_0, _5373} + {_0, _7454};
  wire [2:0] _17209 = {_0, _17207} + {_0, _17208};
  wire [1:0] _17210 = {_0, _9534} + {_0, _11613};
  wire [3:0] _17211 = {_0, _17209} + {_0, _0, _17210};
  wire _17212 = _12301 < _17211;
  wire _17213 = r1502 ^ _17212;
  wire _17214 = _12298 ? coded_block[1502] : r1502;
  wire _17215 = _12296 ? _17213 : _17214;
  always @ (posedge reset or posedge clock) if (reset) r1502 <= 1'd0; else if (_12300) r1502 <= _17215;
  wire [1:0] _17216 = {_0, _34} + {_0, _3901};
  wire [1:0] _17217 = {_0, _5981} + {_0, _8059};
  wire [2:0] _17218 = {_0, _17216} + {_0, _17217};
  wire [1:0] _17219 = {_0, _10141} + {_0, _12219};
  wire [3:0] _17220 = {_0, _17218} + {_0, _0, _17219};
  wire _17221 = _12301 < _17220;
  wire _17222 = r1501 ^ _17221;
  wire _17223 = _12298 ? coded_block[1501] : r1501;
  wire _17224 = _12296 ? _17222 : _17223;
  always @ (posedge reset or posedge clock) if (reset) r1501 <= 1'd0; else if (_12300) r1501 <= _17224;
  wire [1:0] _17225 = {_0, _34} + {_0, _2175};
  wire [1:0] _17226 = {_0, _4256} + {_0, _6334};
  wire [2:0] _17227 = {_0, _17225} + {_0, _17226};
  wire [1:0] _17228 = {_0, _8415} + {_0, _10493};
  wire [3:0] _17229 = {_0, _17227} + {_0, _0, _17228};
  wire _17230 = _12301 < _17229;
  wire _17231 = r1500 ^ _17230;
  wire _17232 = _12298 ? coded_block[1500] : r1500;
  wire _17233 = _12296 ? _17231 : _17232;
  always @ (posedge reset or posedge clock) if (reset) r1500 <= 1'd0; else if (_12300) r1500 <= _17233;
  wire [1:0] _17234 = {_0, _34} + {_0, _4091};
  wire [1:0] _17235 = {_0, _4160} + {_0, _6239};
  wire [2:0] _17236 = {_0, _17234} + {_0, _17235};
  wire [1:0] _17237 = {_0, _8319} + {_0, _10399};
  wire [3:0] _17238 = {_0, _17236} + {_0, _0, _17237};
  wire _17239 = _12301 < _17238;
  wire _17240 = r1499 ^ _17239;
  wire _17241 = _12298 ? coded_block[1499] : r1499;
  wire _17242 = _12296 ? _17240 : _17241;
  always @ (posedge reset or posedge clock) if (reset) r1499 <= 1'd0; else if (_12300) r1499 <= _17242;
  wire [1:0] _17243 = {_0, _34} + {_0, _3359};
  wire [1:0] _17244 = {_0, _5438} + {_0, _7517};
  wire [2:0] _17245 = {_0, _17243} + {_0, _17244};
  wire [1:0] _17246 = {_0, _9597} + {_0, _11677};
  wire [3:0] _17247 = {_0, _17245} + {_0, _0, _17246};
  wire _17248 = _12301 < _17247;
  wire _17249 = r1498 ^ _17248;
  wire _17250 = _12298 ? coded_block[1498] : r1498;
  wire _17251 = _12296 ? _17249 : _17250;
  always @ (posedge reset or posedge clock) if (reset) r1498 <= 1'd0; else if (_12300) r1498 <= _17251;
  wire [1:0] _17252 = {_0, _34} + {_0, _3390};
  wire [1:0] _17253 = {_0, _5470} + {_0, _7548};
  wire [2:0] _17254 = {_0, _17252} + {_0, _17253};
  wire [1:0] _17255 = {_0, _9630} + {_0, _11708};
  wire [3:0] _17256 = {_0, _17254} + {_0, _0, _17255};
  wire _17257 = _12301 < _17256;
  wire _17258 = r1497 ^ _17257;
  wire _17259 = _12298 ? coded_block[1497] : r1497;
  wire _17260 = _12296 ? _17258 : _17259;
  always @ (posedge reset or posedge clock) if (reset) r1497 <= 1'd0; else if (_12300) r1497 <= _17260;
  wire [1:0] _17261 = {_0, _34} + {_0, _2623};
  wire [1:0] _17262 = {_0, _4703} + {_0, _6781};
  wire [2:0] _17263 = {_0, _17261} + {_0, _17262};
  wire [1:0] _17264 = {_0, _8863} + {_0, _10941};
  wire [3:0] _17265 = {_0, _17263} + {_0, _0, _17264};
  wire _17266 = _12301 < _17265;
  wire _17267 = r1496 ^ _17266;
  wire _17268 = _12298 ? coded_block[1496] : r1496;
  wire _17269 = _12296 ? _17267 : _17268;
  always @ (posedge reset or posedge clock) if (reset) r1496 <= 1'd0; else if (_12300) r1496 <= _17269;
  wire [1:0] _17270 = {_0, _1823} + {_0, _2271};
  wire [1:0] _17271 = {_0, _5628} + {_0, _7357};
  wire [2:0] _17272 = {_0, _17270} + {_0, _17271};
  wire [1:0] _17273 = {_0, _9566} + {_0, _11422};
  wire [3:0] _17274 = {_0, _17272} + {_0, _0, _17273};
  wire _17275 = _12301 < _17274;
  wire _17276 = r1495 ^ _17275;
  wire _17277 = _12298 ? coded_block[1495] : r1495;
  wire _17278 = _12296 ? _17276 : _17277;
  always @ (posedge reset or posedge clock) if (reset) r1495 <= 1'd0; else if (_12300) r1495 <= _17278;
  wire [1:0] _17279 = {_0, _1789} + {_0, _3549};
  wire [1:0] _17280 = {_0, _5279} + {_0, _7485};
  wire [2:0] _17281 = {_0, _17279} + {_0, _17280};
  wire [1:0] _17282 = {_0, _9342} + {_0, _11771};
  wire [3:0] _17283 = {_0, _17281} + {_0, _0, _17282};
  wire _17284 = _12301 < _17283;
  wire _17285 = r1494 ^ _17284;
  wire _17286 = _12298 ? coded_block[1494] : r1494;
  wire _17287 = _12296 ? _17285 : _17286;
  always @ (posedge reset or posedge clock) if (reset) r1494 <= 1'd0; else if (_12300) r1494 <= _17287;
  wire [1:0] _17288 = {_0, _1823} + {_0, _4028};
  wire [1:0] _17289 = {_0, _4129} + {_0, _8155};
  wire [2:0] _17290 = {_0, _17288} + {_0, _17289};
  wire [1:0] _17291 = {_0, _8383} + {_0, _11069};
  wire [3:0] _17292 = {_0, _17290} + {_0, _0, _17291};
  wire _17293 = _12301 < _17292;
  wire _17294 = r1493 ^ _17293;
  wire _17295 = _12298 ? coded_block[1493] : r1493;
  wire _17296 = _12296 ? _17294 : _17295;
  always @ (posedge reset or posedge clock) if (reset) r1493 <= 1'd0; else if (_12300) r1493 <= _17296;
  wire [1:0] _17297 = {_0, _1950} + {_0, _3805};
  wire [1:0] _17298 = {_0, _4671} + {_0, _7005};
  wire [2:0] _17299 = {_0, _17297} + {_0, _17298};
  wire [1:0] _17300 = {_0, _8446} + {_0, _10335};
  wire [3:0] _17301 = {_0, _17299} + {_0, _0, _17300};
  wire _17302 = _12301 < _17301;
  wire _17303 = r1492 ^ _17302;
  wire _17304 = _12298 ? coded_block[1492] : r1492;
  wire _17305 = _12296 ? _17303 : _17304;
  always @ (posedge reset or posedge clock) if (reset) r1492 <= 1'd0; else if (_12300) r1492 <= _17305;
  wire [1:0] _17306 = {_0, _1981} + {_0, _3870};
  wire [1:0] _17307 = {_0, _5884} + {_0, _6750};
  wire [2:0] _17308 = {_0, _17306} + {_0, _17307};
  wire [1:0] _17309 = {_0, _9085} + {_0, _10527};
  wire [3:0] _17310 = {_0, _17308} + {_0, _0, _17309};
  wire _17311 = _12301 < _17310;
  wire _17312 = r1491 ^ _17311;
  wire _17313 = _12298 ? coded_block[1491] : r1491;
  wire _17314 = _12296 ? _17312 : _17313;
  always @ (posedge reset or posedge clock) if (reset) r1491 <= 1'd0; else if (_12300) r1491 <= _17314;
  wire [1:0] _17315 = {_0, _2013} + {_0, _2655};
  wire [1:0] _17316 = {_0, _5949} + {_0, _7965};
  wire [2:0] _17317 = {_0, _17315} + {_0, _17316};
  wire [1:0] _17318 = {_0, _8830} + {_0, _11165};
  wire [3:0] _17319 = {_0, _17317} + {_0, _0, _17318};
  wire _17320 = _12301 < _17319;
  wire _17321 = r1490 ^ _17320;
  wire _17322 = _12298 ? coded_block[1490] : r1490;
  wire _17323 = _12296 ? _17321 : _17322;
  always @ (posedge reset or posedge clock) if (reset) r1490 <= 1'd0; else if (_12300) r1490 <= _17323;
  wire [1:0] _17324 = {_0, _2044} + {_0, _3359};
  wire [1:0] _17325 = {_0, _4734} + {_0, _8028};
  wire [2:0] _17326 = {_0, _17324} + {_0, _17325};
  wire [1:0] _17327 = {_0, _10045} + {_0, _10910};
  wire [3:0] _17328 = {_0, _17326} + {_0, _0, _17327};
  wire _17329 = _12301 < _17328;
  wire _17330 = r1489 ^ _17329;
  wire _17331 = _12298 ? coded_block[1489] : r1489;
  wire _17332 = _12296 ? _17330 : _17331;
  always @ (posedge reset or posedge clock) if (reset) r1489 <= 1'd0; else if (_12300) r1489 <= _17332;
  wire [1:0] _17333 = {_0, _65} + {_0, _3262};
  wire [1:0] _17334 = {_0, _5438} + {_0, _6814};
  wire [2:0] _17335 = {_0, _17333} + {_0, _17334};
  wire [1:0] _17336 = {_0, _10108} + {_0, _12124};
  wire [3:0] _17337 = {_0, _17335} + {_0, _0, _17336};
  wire _17338 = _12301 < _17337;
  wire _17339 = r1488 ^ _17338;
  wire _17340 = _12298 ? coded_block[1488] : r1488;
  wire _17341 = _12296 ? _17339 : _17340;
  always @ (posedge reset or posedge clock) if (reset) r1488 <= 1'd0; else if (_12300) r1488 <= _17341;
  wire [1:0] _17342 = {_0, _416} + {_0, _3068};
  wire [1:0] _17343 = {_0, _4350} + {_0, _6366};
  wire [2:0] _17344 = {_0, _17342} + {_0, _17343};
  wire [1:0] _17345 = {_0, _9248} + {_0, _11581};
  wire [3:0] _17346 = {_0, _17344} + {_0, _0, _17345};
  wire _17347 = _12301 < _17346;
  wire _17348 = r1487 ^ _17347;
  wire _17349 = _12298 ? coded_block[1487] : r1487;
  wire _17350 = _12296 ? _17348 : _17349;
  always @ (posedge reset or posedge clock) if (reset) r1487 <= 1'd0; else if (_12300) r1487 <= _17350;
  wire [1:0] _17351 = {_0, _479} + {_0, _3678};
  wire [1:0] _17352 = {_0, _5853} + {_0, _7230};
  wire [2:0] _17353 = {_0, _17351} + {_0, _17352};
  wire [1:0] _17354 = {_0, _8511} + {_0, _10527};
  wire [3:0] _17355 = {_0, _17353} + {_0, _0, _17354};
  wire _17356 = _12301 < _17355;
  wire _17357 = r1486 ^ _17356;
  wire _17358 = _12298 ? coded_block[1486] : r1486;
  wire _17359 = _12296 ? _17357 : _17358;
  always @ (posedge reset or posedge clock) if (reset) r1486 <= 1'd0; else if (_12300) r1486 <= _17359;
  wire [1:0] _17360 = {_0, _1854} + {_0, _2208};
  wire [1:0] _17361 = {_0, _6108} + {_0, _6176};
  wire [2:0] _17362 = {_0, _17360} + {_0, _17361};
  wire [1:0] _17363 = {_0, _10235} + {_0, _10462};
  wire [3:0] _17364 = {_0, _17362} + {_0, _0, _17363};
  wire _17365 = _12301 < _17364;
  wire _17366 = r1485 ^ _17365;
  wire _17367 = _12298 ? coded_block[1485] : r1485;
  wire _17368 = _12296 ? _17366 : _17367;
  always @ (posedge reset or posedge clock) if (reset) r1485 <= 1'd0; else if (_12300) r1485 <= _17368;
  wire [1:0] _17369 = {_0, _1917} + {_0, _2592};
  wire [1:0] _17370 = {_0, _4926} + {_0, _6366};
  wire [2:0] _17371 = {_0, _17369} + {_0, _17370};
  wire [1:0] _17372 = {_0, _8256} + {_0, _10272};
  wire [3:0] _17373 = {_0, _17371} + {_0, _0, _17372};
  wire _17374 = _12301 < _17373;
  wire _17375 = r1484 ^ _17374;
  wire _17376 = _12298 ? coded_block[1484] : r1484;
  wire _17377 = _12296 ? _17375 : _17376;
  always @ (posedge reset or posedge clock) if (reset) r1484 <= 1'd0; else if (_12300) r1484 <= _17377;
  wire [1:0] _17378 = {_0, _510} + {_0, _2175};
  wire [1:0] _17379 = {_0, _5757} + {_0, _7931};
  wire [2:0] _17380 = {_0, _17378} + {_0, _17379};
  wire [1:0] _17381 = {_0, _9311} + {_0, _10590};
  wire [3:0] _17382 = {_0, _17380} + {_0, _0, _17381};
  wire _17383 = _12301 < _17382;
  wire _17384 = r1483 ^ _17383;
  wire _17385 = _12298 ? coded_block[1483] : r1483;
  wire _17386 = _12296 ? _17384 : _17385;
  always @ (posedge reset or posedge clock) if (reset) r1483 <= 1'd0; else if (_12300) r1483 <= _17386;
  wire [1:0] _17387 = {_0, _545} + {_0, _3037};
  wire [1:0] _17388 = {_0, _4256} + {_0, _7837};
  wire [2:0] _17389 = {_0, _17387} + {_0, _17388};
  wire [1:0] _17390 = {_0, _10014} + {_0, _11389};
  wire [3:0] _17391 = {_0, _17389} + {_0, _0, _17390};
  wire _17392 = _12301 < _17391;
  wire _17393 = r1482 ^ _17392;
  wire _17394 = _12298 ? coded_block[1482] : r1482;
  wire _17395 = _12296 ? _17393 : _17394;
  always @ (posedge reset or posedge clock) if (reset) r1482 <= 1'd0; else if (_12300) r1482 <= _17395;
  wire [1:0] _17396 = {_0, _576} + {_0, _2302};
  wire [1:0] _17397 = {_0, _5116} + {_0, _6334};
  wire [2:0] _17398 = {_0, _17396} + {_0, _17397};
  wire [1:0] _17399 = {_0, _9917} + {_0, _12092};
  wire [3:0] _17400 = {_0, _17398} + {_0, _0, _17399};
  wire _17401 = _12301 < _17400;
  wire _17402 = r1481 ^ _17401;
  wire _17403 = _12298 ? coded_block[1481] : r1481;
  wire _17404 = _12296 ? _17402 : _17403;
  always @ (posedge reset or posedge clock) if (reset) r1481 <= 1'd0; else if (_12300) r1481 <= _17404;
  wire [1:0] _17405 = {_0, _608} + {_0, _3359};
  wire [1:0] _17406 = {_0, _4384} + {_0, _7199};
  wire [2:0] _17407 = {_0, _17405} + {_0, _17406};
  wire [1:0] _17408 = {_0, _8415} + {_0, _11996};
  wire [3:0] _17409 = {_0, _17407} + {_0, _0, _17408};
  wire _17410 = _12301 < _17409;
  wire _17411 = r1480 ^ _17410;
  wire _17412 = _12298 ? coded_block[1480] : r1480;
  wire _17413 = _12296 ? _17411 : _17412;
  always @ (posedge reset or posedge clock) if (reset) r1480 <= 1'd0; else if (_12300) r1480 <= _17413;
  wire [1:0] _17414 = {_0, _639} + {_0, _3901};
  wire [1:0] _17415 = {_0, _5438} + {_0, _6462};
  wire [2:0] _17416 = {_0, _17414} + {_0, _17415};
  wire [1:0] _17417 = {_0, _9279} + {_0, _10493};
  wire [3:0] _17418 = {_0, _17416} + {_0, _0, _17417};
  wire _17419 = _12301 < _17418;
  wire _17420 = r1479 ^ _17419;
  wire _17421 = _12298 ? coded_block[1479] : r1479;
  wire _17422 = _12296 ? _17420 : _17421;
  always @ (posedge reset or posedge clock) if (reset) r1479 <= 1'd0; else if (_12300) r1479 <= _17422;
  wire [1:0] _17423 = {_0, _672} + {_0, _2974};
  wire [1:0] _17424 = {_0, _5981} + {_0, _7517};
  wire [2:0] _17425 = {_0, _17423} + {_0, _17424};
  wire [1:0] _17426 = {_0, _8543} + {_0, _11358};
  wire [3:0] _17427 = {_0, _17425} + {_0, _0, _17426};
  wire _17428 = _12301 < _17427;
  wire _17429 = r1478 ^ _17428;
  wire _17430 = _12298 ? coded_block[1478] : r1478;
  wire _17431 = _12296 ? _17429 : _17430;
  always @ (posedge reset or posedge clock) if (reset) r1478 <= 1'd0; else if (_12300) r1478 <= _17431;
  wire [1:0] _17432 = {_0, _703} + {_0, _3294};
  wire [1:0] _17433 = {_0, _5053} + {_0, _8059};
  wire [2:0] _17434 = {_0, _17432} + {_0, _17433};
  wire [1:0] _17435 = {_0, _9597} + {_0, _10621};
  wire [3:0] _17436 = {_0, _17434} + {_0, _0, _17435};
  wire _17437 = _12301 < _17436;
  wire _17438 = r1477 ^ _17437;
  wire _17439 = _12298 ? coded_block[1477] : r1477;
  wire _17440 = _12296 ? _17438 : _17439;
  always @ (posedge reset or posedge clock) if (reset) r1477 <= 1'd0; else if (_12300) r1477 <= _17440;
  wire [1:0] _17441 = {_0, _766} + {_0, _3104};
  wire [1:0] _17442 = {_0, _5821} + {_0, _7454};
  wire [2:0] _17443 = {_0, _17441} + {_0, _17442};
  wire [1:0] _17444 = {_0, _9212} + {_0, _12219};
  wire [3:0] _17445 = {_0, _17443} + {_0, _0, _17444};
  wire _17446 = _12301 < _17445;
  wire _17447 = r1476 ^ _17446;
  wire _17448 = _12298 ? coded_block[1476] : r1476;
  wire _17449 = _12296 ? _17447 : _17448;
  always @ (posedge reset or posedge clock) if (reset) r1476 <= 1'd0; else if (_12300) r1476 <= _17449;
  wire [1:0] _17450 = {_0, _1758} + {_0, _2463};
  wire [1:0] _17451 = {_0, _5085} + {_0, _7069};
  wire [2:0] _17452 = {_0, _17450} + {_0, _17451};
  wire [1:0] _17453 = {_0, _10235} + {_0, _10941};
  wire [3:0] _17454 = {_0, _17452} + {_0, _0, _17453};
  wire _17455 = _12301 < _17454;
  wire _17456 = r1475 ^ _17455;
  wire _17457 = _12298 ? coded_block[1475] : r1475;
  wire _17458 = _12296 ? _17456 : _17457;
  always @ (posedge reset or posedge clock) if (reset) r1475 <= 1'd0; else if (_12300) r1475 <= _17458;
  wire [1:0] _17459 = {_0, _1789} + {_0, _2719};
  wire [1:0] _17460 = {_0, _4542} + {_0, _7163};
  wire [2:0] _17461 = {_0, _17459} + {_0, _17460};
  wire [1:0] _17462 = {_0, _9149} + {_0, _10303};
  wire [3:0] _17463 = {_0, _17461} + {_0, _0, _17462};
  wire _17464 = _12301 < _17463;
  wire _17465 = r1474 ^ _17464;
  wire _17466 = _12298 ? coded_block[1474] : r1474;
  wire _17467 = _12296 ? _17465 : _17466;
  always @ (posedge reset or posedge clock) if (reset) r1474 <= 1'd0; else if (_12300) r1474 <= _17467;
  wire [1:0] _17468 = {_0, _1823} + {_0, _3615};
  wire [1:0] _17469 = {_0, _4798} + {_0, _6621};
  wire [2:0] _17470 = {_0, _17468} + {_0, _17469};
  wire [1:0] _17471 = {_0, _9248} + {_0, _11228};
  wire [3:0] _17472 = {_0, _17470} + {_0, _0, _17471};
  wire _17473 = _12301 < _17472;
  wire _17474 = r1473 ^ _17473;
  wire _17475 = _12298 ? coded_block[1473] : r1473;
  wire _17476 = _12296 ? _17474 : _17475;
  always @ (posedge reset or posedge clock) if (reset) r1473 <= 1'd0; else if (_12300) r1473 <= _17476;
  wire [1:0] _17477 = {_0, _1854} + {_0, _3262};
  wire [1:0] _17478 = {_0, _5694} + {_0, _6877};
  wire [2:0] _17479 = {_0, _17477} + {_0, _17478};
  wire [1:0] _17480 = {_0, _8701} + {_0, _11326};
  wire [3:0] _17481 = {_0, _17479} + {_0, _0, _17480};
  wire _17482 = _12301 < _17481;
  wire _17483 = r1472 ^ _17482;
  wire _17484 = _12298 ? coded_block[1472] : r1472;
  wire _17485 = _12296 ? _17483 : _17484;
  always @ (posedge reset or posedge clock) if (reset) r1472 <= 1'd0; else if (_12300) r1472 <= _17485;
  wire [1:0] _17486 = {_0, _1886} + {_0, _3486};
  wire [1:0] _17487 = {_0, _5342} + {_0, _7773};
  wire [2:0] _17488 = {_0, _17486} + {_0, _17487};
  wire [1:0] _17489 = {_0, _8957} + {_0, _10783};
  wire [3:0] _17490 = {_0, _17488} + {_0, _0, _17489};
  wire _17491 = _12301 < _17490;
  wire _17492 = r1471 ^ _17491;
  wire _17493 = _12298 ? coded_block[1471] : r1471;
  wire _17494 = _12296 ? _17492 : _17493;
  always @ (posedge reset or posedge clock) if (reset) r1471 <= 1'd0; else if (_12300) r1471 <= _17494;
  wire [1:0] _17495 = {_0, _1917} + {_0, _3359};
  wire [1:0] _17496 = {_0, _5565} + {_0, _7420};
  wire [2:0] _17497 = {_0, _17495} + {_0, _17496};
  wire [1:0] _17498 = {_0, _9853} + {_0, _11038};
  wire [3:0] _17499 = {_0, _17497} + {_0, _0, _17498};
  wire _17500 = _12301 < _17499;
  wire _17501 = r1470 ^ _17500;
  wire _17502 = _12298 ? coded_block[1470] : r1470;
  wire _17503 = _12296 ? _17501 : _17502;
  always @ (posedge reset or posedge clock) if (reset) r1470 <= 1'd0; else if (_12300) r1470 <= _17503;
  wire [1:0] _17504 = {_0, _1950} + {_0, _3709};
  wire [1:0] _17505 = {_0, _5438} + {_0, _7644};
  wire [2:0] _17506 = {_0, _17504} + {_0, _17505};
  wire [1:0] _17507 = {_0, _9503} + {_0, _11933};
  wire [3:0] _17508 = {_0, _17506} + {_0, _0, _17507};
  wire _17509 = _12301 < _17508;
  wire _17510 = r1469 ^ _17509;
  wire _17511 = _12298 ? coded_block[1469] : r1469;
  wire _17512 = _12296 ? _17510 : _17511;
  always @ (posedge reset or posedge clock) if (reset) r1469 <= 1'd0; else if (_12300) r1469 <= _17512;
  wire [1:0] _17513 = {_0, _1981} + {_0, _2430};
  wire [1:0] _17514 = {_0, _5790} + {_0, _7517};
  wire [2:0] _17515 = {_0, _17513} + {_0, _17514};
  wire [1:0] _17516 = {_0, _9724} + {_0, _11581};
  wire [3:0] _17517 = {_0, _17515} + {_0, _0, _17516};
  wire _17518 = _12301 < _17517;
  wire _17519 = r1468 ^ _17518;
  wire _17520 = _12298 ? coded_block[1468] : r1468;
  wire _17521 = _12296 ? _17519 : _17520;
  always @ (posedge reset or posedge clock) if (reset) r1468 <= 1'd0; else if (_12300) r1468 <= _17521;
  wire [1:0] _17522 = {_0, _2013} + {_0, _3037};
  wire [1:0] _17523 = {_0, _4511} + {_0, _7868};
  wire [2:0] _17524 = {_0, _17522} + {_0, _17523};
  wire [1:0] _17525 = {_0, _9597} + {_0, _11806};
  wire [3:0] _17526 = {_0, _17524} + {_0, _0, _17525};
  wire _17527 = _12301 < _17526;
  wire _17528 = r1467 ^ _17527;
  wire _17529 = _12298 ? coded_block[1467] : r1467;
  wire _17530 = _12296 ? _17528 : _17529;
  always @ (posedge reset or posedge clock) if (reset) r1467 <= 1'd0; else if (_12300) r1467 <= _17530;
  wire [1:0] _17531 = {_0, _831} + {_0, _2112};
  wire [1:0] _17532 = {_0, _6108} + {_0, _7262};
  wire [2:0] _17533 = {_0, _17531} + {_0, _17532};
  wire [1:0] _17534 = {_0, _9980} + {_0, _11613};
  wire [3:0] _17535 = {_0, _17533} + {_0, _0, _17534};
  wire _17536 = _12301 < _17535;
  wire _17537 = r1466 ^ _17536;
  wire _17538 = _12298 ? coded_block[1466] : r1466;
  wire _17539 = _12296 ? _17537 : _17538;
  always @ (posedge reset or posedge clock) if (reset) r1466 <= 1'd0; else if (_12300) r1466 <= _17539;
  wire [1:0] _17540 = {_0, _863} + {_0, _3580};
  wire [1:0] _17541 = {_0, _4192} + {_0, _8186};
  wire [2:0] _17542 = {_0, _17540} + {_0, _17541};
  wire [1:0] _17543 = {_0, _9342} + {_0, _12061};
  wire [3:0] _17544 = {_0, _17542} + {_0, _0, _17543};
  wire _17545 = _12301 < _17544;
  wire _17546 = r1465 ^ _17545;
  wire _17547 = _12298 ? coded_block[1465] : r1465;
  wire _17548 = _12296 ? _17546 : _17547;
  always @ (posedge reset or posedge clock) if (reset) r1465 <= 1'd0; else if (_12300) r1465 <= _17548;
  wire [1:0] _17549 = {_0, _894} + {_0, _3836};
  wire [1:0] _17550 = {_0, _5663} + {_0, _6270};
  wire [2:0] _17551 = {_0, _17549} + {_0, _17550};
  wire [1:0] _17552 = {_0, _8256} + {_0, _11422};
  wire [3:0] _17553 = {_0, _17551} + {_0, _0, _17552};
  wire _17554 = _12301 < _17553;
  wire _17555 = r1464 ^ _17554;
  wire _17556 = _12298 ? coded_block[1464] : r1464;
  wire _17557 = _12296 ? _17555 : _17556;
  always @ (posedge reset or posedge clock) if (reset) r1464 <= 1'd0; else if (_12300) r1464 <= _17557;
  wire [1:0] _17558 = {_0, _927} + {_0, _2719};
  wire [1:0] _17559 = {_0, _5918} + {_0, _7741};
  wire [2:0] _17560 = {_0, _17558} + {_0, _17559};
  wire [1:0] _17561 = {_0, _8352} + {_0, _10335};
  wire [3:0] _17562 = {_0, _17560} + {_0, _0, _17561};
  wire _17563 = _12301 < _17562;
  wire _17564 = r1463 ^ _17563;
  wire _17565 = _12298 ? coded_block[1463] : r1463;
  wire _17566 = _12296 ? _17564 : _17565;
  always @ (posedge reset or posedge clock) if (reset) r1463 <= 1'd0; else if (_12300) r1463 <= _17566;
  wire [1:0] _17567 = {_0, _958} + {_0, _2367};
  wire [1:0] _17568 = {_0, _4798} + {_0, _7996};
  wire [2:0] _17569 = {_0, _17567} + {_0, _17568};
  wire [1:0] _17570 = {_0, _9822} + {_0, _10430};
  wire [3:0] _17571 = {_0, _17569} + {_0, _0, _17570};
  wire _17572 = _12301 < _17571;
  wire _17573 = r1462 ^ _17572;
  wire _17574 = _12298 ? coded_block[1462] : r1462;
  wire _17575 = _12296 ? _17573 : _17574;
  always @ (posedge reset or posedge clock) if (reset) r1462 <= 1'd0; else if (_12300) r1462 <= _17575;
  wire [1:0] _17576 = {_0, _990} + {_0, _2592};
  wire [1:0] _17577 = {_0, _4447} + {_0, _6877};
  wire [2:0] _17578 = {_0, _17576} + {_0, _17577};
  wire [1:0] _17579 = {_0, _10077} + {_0, _11900};
  wire [3:0] _17580 = {_0, _17578} + {_0, _0, _17579};
  wire _17581 = _12301 < _17580;
  wire _17582 = r1461 ^ _17581;
  wire _17583 = _12298 ? coded_block[1461] : r1461;
  wire _17584 = _12296 ? _17582 : _17583;
  always @ (posedge reset or posedge clock) if (reset) r1461 <= 1'd0; else if (_12300) r1461 <= _17584;
  wire [1:0] _17585 = {_0, _1021} + {_0, _2463};
  wire [1:0] _17586 = {_0, _4671} + {_0, _6525};
  wire [2:0] _17587 = {_0, _17585} + {_0, _17586};
  wire [1:0] _17588 = {_0, _8957} + {_0, _12155};
  wire [3:0] _17589 = {_0, _17587} + {_0, _0, _17588};
  wire _17590 = _12301 < _17589;
  wire _17591 = r1460 ^ _17590;
  wire _17592 = _12298 ? coded_block[1460] : r1460;
  wire _17593 = _12296 ? _17591 : _17592;
  always @ (posedge reset or posedge clock) if (reset) r1460 <= 1'd0; else if (_12300) r1460 <= _17593;
  wire [1:0] _17594 = {_0, _1057} + {_0, _2813};
  wire [1:0] _17595 = {_0, _4542} + {_0, _6750};
  wire [2:0] _17596 = {_0, _17594} + {_0, _17595};
  wire [1:0] _17597 = {_0, _8607} + {_0, _11038};
  wire [3:0] _17598 = {_0, _17596} + {_0, _0, _17597};
  wire _17599 = _12301 < _17598;
  wire _17600 = r1459 ^ _17599;
  wire _17601 = _12298 ? coded_block[1459] : r1459;
  wire _17602 = _12296 ? _17600 : _17601;
  always @ (posedge reset or posedge clock) if (reset) r1459 <= 1'd0; else if (_12300) r1459 <= _17602;
  wire [1:0] _17603 = {_0, _1088} + {_0, _3549};
  wire [1:0] _17604 = {_0, _4895} + {_0, _6621};
  wire [2:0] _17605 = {_0, _17603} + {_0, _17604};
  wire [1:0] _17606 = {_0, _8830} + {_0, _10685};
  wire [3:0] _17607 = {_0, _17605} + {_0, _0, _17606};
  wire _17608 = _12301 < _17607;
  wire _17609 = r1458 ^ _17608;
  wire _17610 = _12298 ? coded_block[1458] : r1458;
  wire _17611 = _12296 ? _17609 : _17610;
  always @ (posedge reset or posedge clock) if (reset) r1458 <= 1'd0; else if (_12300) r1458 <= _17611;
  wire [1:0] _17612 = {_0, _1662} + {_0, _3997};
  wire [1:0] _17613 = {_0, _4703} + {_0, _6334};
  wire [2:0] _17614 = {_0, _17612} + {_0, _17613};
  wire [1:0] _17615 = {_0, _10108} + {_0, _11101};
  wire [3:0] _17616 = {_0, _17614} + {_0, _0, _17615};
  wire _17617 = _12301 < _17616;
  wire _17618 = r1457 ^ _17617;
  wire _17619 = _12298 ? coded_block[1457] : r1457;
  wire _17620 = _12296 ? _17618 : _17619;
  always @ (posedge reset or posedge clock) if (reset) r1457 <= 1'd0; else if (_12300) r1457 <= _17620;
  wire [1:0] _17621 = {_0, _1726} + {_0, _3005};
  wire [1:0] _17622 = {_0, _4989} + {_0, _8155};
  wire [2:0] _17623 = {_0, _17621} + {_0, _17622};
  wire [1:0] _17624 = {_0, _8863} + {_0, _10493};
  wire [3:0] _17625 = {_0, _17623} + {_0, _0, _17624};
  wire _17626 = _12301 < _17625;
  wire _17627 = r1456 ^ _17626;
  wire _17628 = _12298 ? coded_block[1456] : r1456;
  wire _17629 = _12296 ? _17627 : _17628;
  always @ (posedge reset or posedge clock) if (reset) r1456 <= 1'd0; else if (_12300) r1456 <= _17629;
  wire [1:0] _17630 = {_0, _352} + {_0, _2719};
  wire [1:0] _17631 = {_0, _4605} + {_0, _6176};
  wire [2:0] _17632 = {_0, _17630} + {_0, _17631};
  wire [1:0] _17633 = {_0, _8736} + {_0, _10973};
  wire [3:0] _17634 = {_0, _17632} + {_0, _0, _17633};
  wire _17635 = _12301 < _17634;
  wire _17636 = r1455 ^ _17635;
  wire _17637 = _12298 ? coded_block[1455] : r1455;
  wire _17638 = _12296 ? _17636 : _17637;
  always @ (posedge reset or posedge clock) if (reset) r1455 <= 1'd0; else if (_12300) r1455 <= _17638;
  wire [1:0] _17639 = {_0, _383} + {_0, _3359};
  wire [1:0] _17640 = {_0, _4798} + {_0, _6687};
  wire [2:0] _17641 = {_0, _17639} + {_0, _17640};
  wire [1:0] _17642 = {_0, _8225} + {_0, _10814};
  wire [3:0] _17643 = {_0, _17641} + {_0, _0, _17642};
  wire _17644 = _12301 < _17643;
  wire _17645 = r1454 ^ _17644;
  wire _17646 = _12298 ? coded_block[1454] : r1454;
  wire _17647 = _12296 ? _17645 : _17646;
  always @ (posedge reset or posedge clock) if (reset) r1454 <= 1'd0; else if (_12300) r1454 <= _17647;
  wire [1:0] _17648 = {_0, _416} + {_0, _3104};
  wire [1:0] _17649 = {_0, _5438} + {_0, _6877};
  wire [2:0] _17650 = {_0, _17648} + {_0, _17649};
  wire [1:0] _17651 = {_0, _8767} + {_0, _10272};
  wire [3:0] _17652 = {_0, _17650} + {_0, _0, _17651};
  wire _17653 = _12301 < _17652;
  wire _17654 = r1453 ^ _17653;
  wire _17655 = _12298 ? coded_block[1453] : r1453;
  wire _17656 = _12296 ? _17654 : _17655;
  always @ (posedge reset or posedge clock) if (reset) r1453 <= 1'd0; else if (_12300) r1453 <= _17656;
  wire [1:0] _17657 = {_0, _447} + {_0, _2302};
  wire [1:0] _17658 = {_0, _5183} + {_0, _7517};
  wire [2:0] _17659 = {_0, _17657} + {_0, _17658};
  wire [1:0] _17660 = {_0, _8957} + {_0, _10846};
  wire [3:0] _17661 = {_0, _17659} + {_0, _0, _17660};
  wire _17662 = _12301 < _17661;
  wire _17663 = r1452 ^ _17662;
  wire _17664 = _12298 ? coded_block[1452] : r1452;
  wire _17665 = _12296 ? _17663 : _17664;
  always @ (posedge reset or posedge clock) if (reset) r1452 <= 1'd0; else if (_12300) r1452 <= _17665;
  wire [1:0] _17666 = {_0, _479} + {_0, _2367};
  wire [1:0] _17667 = {_0, _4384} + {_0, _7262};
  wire [2:0] _17668 = {_0, _17666} + {_0, _17667};
  wire [1:0] _17669 = {_0, _9597} + {_0, _11038};
  wire [3:0] _17670 = {_0, _17668} + {_0, _0, _17669};
  wire _17671 = _12301 < _17670;
  wire _17672 = r1451 ^ _17671;
  wire _17673 = _12298 ? coded_block[1451] : r1451;
  wire _17674 = _12296 ? _17672 : _17673;
  always @ (posedge reset or posedge clock) if (reset) r1451 <= 1'd0; else if (_12300) r1451 <= _17674;
  wire [1:0] _17675 = {_0, _510} + {_0, _3167};
  wire [1:0] _17676 = {_0, _4447} + {_0, _6462};
  wire [2:0] _17677 = {_0, _17675} + {_0, _17676};
  wire [1:0] _17678 = {_0, _9342} + {_0, _11677};
  wire [3:0] _17679 = {_0, _17677} + {_0, _0, _17678};
  wire _17680 = _12301 < _17679;
  wire _17681 = r1450 ^ _17680;
  wire _17682 = _12298 ? coded_block[1450] : r1450;
  wire _17683 = _12296 ? _17681 : _17682;
  always @ (posedge reset or posedge clock) if (reset) r1450 <= 1'd0; else if (_12300) r1450 <= _17683;
  wire [1:0] _17684 = {_0, _576} + {_0, _3773};
  wire [1:0] _17685 = {_0, _5949} + {_0, _7326};
  wire [2:0] _17686 = {_0, _17684} + {_0, _17685};
  wire [1:0] _17687 = {_0, _8607} + {_0, _10621};
  wire [3:0] _17688 = {_0, _17686} + {_0, _0, _17687};
  wire _17689 = _12301 < _17688;
  wire _17690 = r1449 ^ _17689;
  wire _17691 = _12298 ? coded_block[1449] : r1449;
  wire _17692 = _12296 ? _17690 : _17691;
  always @ (posedge reset or posedge clock) if (reset) r1449 <= 1'd0; else if (_12300) r1449 <= _17692;
  wire [1:0] _17693 = {_0, _608} + {_0, _2271};
  wire [1:0] _17694 = {_0, _5853} + {_0, _8028};
  wire [2:0] _17695 = {_0, _17693} + {_0, _17694};
  wire [1:0] _17696 = {_0, _9406} + {_0, _10685};
  wire [3:0] _17697 = {_0, _17695} + {_0, _0, _17696};
  wire _17698 = _12301 < _17697;
  wire _17699 = r1448 ^ _17698;
  wire _17700 = _12298 ? coded_block[1448] : r1448;
  wire _17701 = _12296 ? _17699 : _17700;
  always @ (posedge reset or posedge clock) if (reset) r1448 <= 1'd0; else if (_12300) r1448 <= _17701;
  wire [1:0] _17702 = {_0, _639} + {_0, _3135};
  wire [1:0] _17703 = {_0, _4350} + {_0, _7931};
  wire [2:0] _17704 = {_0, _17702} + {_0, _17703};
  wire [1:0] _17705 = {_0, _10108} + {_0, _11485};
  wire [3:0] _17706 = {_0, _17704} + {_0, _0, _17705};
  wire _17707 = _12301 < _17706;
  wire _17708 = r1447 ^ _17707;
  wire _17709 = _12298 ? coded_block[1447] : r1447;
  wire _17710 = _12296 ? _17708 : _17709;
  always @ (posedge reset or posedge clock) if (reset) r1447 <= 1'd0; else if (_12300) r1447 <= _17710;
  wire [1:0] _17711 = {_0, _672} + {_0, _2399};
  wire [1:0] _17712 = {_0, _5215} + {_0, _6431};
  wire [2:0] _17713 = {_0, _17711} + {_0, _17712};
  wire [1:0] _17714 = {_0, _10014} + {_0, _12188};
  wire [3:0] _17715 = {_0, _17713} + {_0, _0, _17714};
  wire _17716 = _12301 < _17715;
  wire _17717 = r1446 ^ _17716;
  wire _17718 = _12298 ? coded_block[1446] : r1446;
  wire _17719 = _12296 ? _17717 : _17718;
  always @ (posedge reset or posedge clock) if (reset) r1446 <= 1'd0; else if (_12300) r1446 <= _17719;
  wire [1:0] _17720 = {_0, _703} + {_0, _3453};
  wire [1:0] _17721 = {_0, _4478} + {_0, _7293};
  wire [2:0] _17722 = {_0, _17720} + {_0, _17721};
  wire [1:0] _17723 = {_0, _8511} + {_0, _12092};
  wire [3:0] _17724 = {_0, _17722} + {_0, _0, _17723};
  wire _17725 = _12301 < _17724;
  wire _17726 = r1445 ^ _17725;
  wire _17727 = _12298 ? coded_block[1445] : r1445;
  wire _17728 = _12296 ? _17726 : _17727;
  always @ (posedge reset or posedge clock) if (reset) r1445 <= 1'd0; else if (_12300) r1445 <= _17728;
  wire [1:0] _17729 = {_0, _766} + {_0, _3068};
  wire [1:0] _17730 = {_0, _6076} + {_0, _7612};
  wire [2:0] _17731 = {_0, _17729} + {_0, _17730};
  wire [1:0] _17732 = {_0, _8638} + {_0, _11453};
  wire [3:0] _17733 = {_0, _17731} + {_0, _0, _17732};
  wire _17734 = _12301 < _17733;
  wire _17735 = r1444 ^ _17734;
  wire _17736 = _12298 ? coded_block[1444] : r1444;
  wire _17737 = _12296 ? _17735 : _17736;
  always @ (posedge reset or posedge clock) if (reset) r1444 <= 1'd0; else if (_12300) r1444 <= _17737;
  wire [1:0] _17738 = {_0, _800} + {_0, _3390};
  wire [1:0] _17739 = {_0, _5152} + {_0, _8155};
  wire [2:0] _17740 = {_0, _17738} + {_0, _17739};
  wire [1:0] _17741 = {_0, _9693} + {_0, _10717};
  wire [3:0] _17742 = {_0, _17740} + {_0, _0, _17741};
  wire _17743 = _12301 < _17742;
  wire _17744 = r1443 ^ _17743;
  wire _17745 = _12298 ? coded_block[1443] : r1443;
  wire _17746 = _12296 ? _17744 : _17745;
  always @ (posedge reset or posedge clock) if (reset) r1443 <= 1'd0; else if (_12300) r1443 <= _17746;
  wire [1:0] _17747 = {_0, _65} + {_0, _2208};
  wire [1:0] _17748 = {_0, _4671} + {_0, _7199};
  wire [2:0] _17749 = {_0, _17747} + {_0, _17748};
  wire [1:0] _17750 = {_0, _8670} + {_0, _12027};
  wire [3:0] _17751 = {_0, _17749} + {_0, _0, _17750};
  wire _17752 = _12301 < _17751;
  wire _17753 = r1442 ^ _17752;
  wire _17754 = _12298 ? coded_block[1442] : r1442;
  wire _17755 = _12296 ? _17753 : _17754;
  always @ (posedge reset or posedge clock) if (reset) r1442 <= 1'd0; else if (_12300) r1442 <= _17755;
  wire [1:0] _17756 = {_0, _97} + {_0, _3231};
  wire [1:0] _17757 = {_0, _4287} + {_0, _6750};
  wire [2:0] _17758 = {_0, _17756} + {_0, _17757};
  wire [1:0] _17759 = {_0, _9279} + {_0, _10748};
  wire [3:0] _17760 = {_0, _17758} + {_0, _0, _17759};
  wire _17761 = _12301 < _17760;
  wire _17762 = r1441 ^ _17761;
  wire _17763 = _12298 ? coded_block[1441] : r1441;
  wire _17764 = _12296 ? _17762 : _17763;
  always @ (posedge reset or posedge clock) if (reset) r1441 <= 1'd0; else if (_12300) r1441 <= _17764;
  wire [1:0] _17765 = {_0, _128} + {_0, _3646};
  wire [1:0] _17766 = {_0, _5310} + {_0, _6366};
  wire [2:0] _17767 = {_0, _17765} + {_0, _17766};
  wire [1:0] _17768 = {_0, _8830} + {_0, _11358};
  wire [3:0] _17769 = {_0, _17767} + {_0, _0, _17768};
  wire _17770 = _12301 < _17769;
  wire _17771 = r1440 ^ _17770;
  wire _17772 = _12298 ? coded_block[1440] : r1440;
  wire _17773 = _12296 ? _17771 : _17772;
  always @ (posedge reset or posedge clock) if (reset) r1440 <= 1'd0; else if (_12300) r1440 <= _17773;
  wire [1:0] _17774 = {_0, _192} + {_0, _3549};
  wire [1:0] _17775 = {_0, _4192} + {_0, _7804};
  wire [2:0] _17776 = {_0, _17774} + {_0, _17775};
  wire [1:0] _17777 = {_0, _9469} + {_0, _10527};
  wire [3:0] _17778 = {_0, _17776} + {_0, _0, _17777};
  wire _17779 = _12301 < _17778;
  wire _17780 = r1439 ^ _17779;
  wire _17781 = _12298 ? coded_block[1439] : r1439;
  wire _17782 = _12296 ? _17780 : _17781;
  always @ (posedge reset or posedge clock) if (reset) r1439 <= 1'd0; else if (_12300) r1439 <= _17782;
  wire [1:0] _17783 = {_0, _224} + {_0, _2847};
  wire [1:0] _17784 = {_0, _5628} + {_0, _6270};
  wire [2:0] _17785 = {_0, _17783} + {_0, _17784};
  wire [1:0] _17786 = {_0, _9886} + {_0, _11550};
  wire [3:0] _17787 = {_0, _17785} + {_0, _0, _17786};
  wire _17788 = _12301 < _17787;
  wire _17789 = r1438 ^ _17788;
  wire _17790 = _12298 ? coded_block[1438] : r1438;
  wire _17791 = _12296 ? _17789 : _17790;
  always @ (posedge reset or posedge clock) if (reset) r1438 <= 1'd0; else if (_12300) r1438 <= _17791;
  wire [1:0] _17792 = {_0, _255} + {_0, _2526};
  wire [1:0] _17793 = {_0, _4926} + {_0, _7710};
  wire [2:0] _17794 = {_0, _17792} + {_0, _17793};
  wire [1:0] _17795 = {_0, _8352} + {_0, _11964};
  wire [3:0] _17796 = {_0, _17794} + {_0, _0, _17795};
  wire _17797 = _12301 < _17796;
  wire _17798 = r1437 ^ _17797;
  wire _17799 = _12298 ? coded_block[1437] : r1437;
  wire _17800 = _12296 ? _17798 : _17799;
  always @ (posedge reset or posedge clock) if (reset) r1437 <= 1'd0; else if (_12300) r1437 <= _17800;
  wire [1:0] _17801 = {_0, _289} + {_0, _2686};
  wire [1:0] _17802 = {_0, _4605} + {_0, _7005};
  wire [2:0] _17803 = {_0, _17801} + {_0, _17802};
  wire [1:0] _17804 = {_0, _9790} + {_0, _10430};
  wire [3:0] _17805 = {_0, _17803} + {_0, _0, _17804};
  wire _17806 = _12301 < _17805;
  wire _17807 = r1436 ^ _17806;
  wire _17808 = _12298 ? coded_block[1436] : r1436;
  wire _17809 = _12296 ? _17807 : _17808;
  always @ (posedge reset or posedge clock) if (reset) r1436 <= 1'd0; else if (_12300) r1436 <= _17809;
  wire [1:0] _17810 = {_0, _320} + {_0, _2494};
  wire [1:0] _17811 = {_0, _4767} + {_0, _6687};
  wire [2:0] _17812 = {_0, _17810} + {_0, _17811};
  wire [1:0] _17813 = {_0, _9085} + {_0, _11869};
  wire [3:0] _17814 = {_0, _17812} + {_0, _0, _17813};
  wire _17815 = _12301 < _17814;
  wire _17816 = r1435 ^ _17815;
  wire _17817 = _12298 ? coded_block[1435] : r1435;
  wire _17818 = _12296 ? _17816 : _17817;
  always @ (posedge reset or posedge clock) if (reset) r1435 <= 1'd0; else if (_12300) r1435 <= _17818;
  wire [1:0] _17819 = {_0, _383} + {_0, _4028};
  wire [1:0] _17820 = {_0, _4958} + {_0, _6652};
  wire [2:0] _17821 = {_0, _17819} + {_0, _17820};
  wire [1:0] _17822 = {_0, _8926} + {_0, _10846};
  wire [3:0] _17823 = {_0, _17821} + {_0, _0, _17822};
  wire _17824 = _12301 < _17823;
  wire _17825 = r1434 ^ _17824;
  wire _17826 = _12298 ? coded_block[1434] : r1434;
  wire _17827 = _12296 ? _17825 : _17826;
  always @ (posedge reset or posedge clock) if (reset) r1434 <= 1'd0; else if (_12300) r1434 <= _17827;
  wire [1:0] _17828 = {_0, _416} + {_0, _3805};
  wire [1:0] _17829 = {_0, _6108} + {_0, _7036};
  wire [2:0] _17830 = {_0, _17828} + {_0, _17829};
  wire [1:0] _17831 = {_0, _8736} + {_0, _11004};
  wire [3:0] _17832 = {_0, _17830} + {_0, _0, _17831};
  wire _17833 = _12301 < _17832;
  wire _17834 = r1433 ^ _17833;
  wire _17835 = _12298 ? coded_block[1433] : r1433;
  wire _17836 = _12296 ? _17834 : _17835;
  always @ (posedge reset or posedge clock) if (reset) r1433 <= 1'd0; else if (_12300) r1433 <= _17836;
  wire [1:0] _17837 = {_0, _447} + {_0, _2367};
  wire [1:0] _17838 = {_0, _5884} + {_0, _8186};
  wire [2:0] _17839 = {_0, _17837} + {_0, _17838};
  wire [1:0] _17840 = {_0, _9118} + {_0, _10814};
  wire [3:0] _17841 = {_0, _17839} + {_0, _0, _17840};
  wire _17842 = _12301 < _17841;
  wire _17843 = r1432 ^ _17842;
  wire _17844 = _12298 ? coded_block[1432] : r1432;
  wire _17845 = _12296 ? _17843 : _17844;
  always @ (posedge reset or posedge clock) if (reset) r1432 <= 1'd0; else if (_12300) r1432 <= _17845;
  wire [1:0] _17846 = {_0, _479} + {_0, _2302};
  wire [1:0] _17847 = {_0, _4447} + {_0, _7965};
  wire [2:0] _17848 = {_0, _17846} + {_0, _17847};
  wire [1:0] _17849 = {_0, _8256} + {_0, _11196};
  wire [3:0] _17850 = {_0, _17848} + {_0, _0, _17849};
  wire _17851 = _12301 < _17850;
  wire _17852 = r1431 ^ _17851;
  wire _17853 = _12298 ? coded_block[1431] : r1431;
  wire _17854 = _12296 ? _17852 : _17853;
  always @ (posedge reset or posedge clock) if (reset) r1431 <= 1'd0; else if (_12300) r1431 <= _17854;
  wire [1:0] _17855 = {_0, _545} + {_0, _4091};
  wire [1:0] _17856 = {_0, _5501} + {_0, _6462};
  wire [2:0] _17857 = {_0, _17855} + {_0, _17856};
  wire [1:0] _17858 = {_0, _8607} + {_0, _12124};
  wire [3:0] _17859 = {_0, _17857} + {_0, _0, _17858};
  wire _17860 = _12301 < _17859;
  wire _17861 = r1430 ^ _17860;
  wire _17862 = _12298 ? coded_block[1430] : r1430;
  wire _17863 = _12296 ? _17861 : _17862;
  always @ (posedge reset or posedge clock) if (reset) r1430 <= 1'd0; else if (_12300) r1430 <= _17863;
  wire [1:0] _17864 = {_0, _576} + {_0, _3678};
  wire [1:0] _17865 = {_0, _4160} + {_0, _7581};
  wire [2:0] _17866 = {_0, _17864} + {_0, _17865};
  wire [1:0] _17867 = {_0, _8543} + {_0, _10685};
  wire [3:0] _17868 = {_0, _17866} + {_0, _0, _17867};
  wire _17869 = _12301 < _17868;
  wire _17870 = r1429 ^ _17869;
  wire _17871 = _12298 ? coded_block[1429] : r1429;
  wire _17872 = _12296 ? _17870 : _17871;
  always @ (posedge reset or posedge clock) if (reset) r1429 <= 1'd0; else if (_12300) r1429 <= _17872;
  wire [1:0] _17873 = {_0, _608} + {_0, _3390};
  wire [1:0] _17874 = {_0, _5757} + {_0, _6239};
  wire [2:0] _17875 = {_0, _17873} + {_0, _17874};
  wire [1:0] _17876 = {_0, _9661} + {_0, _10621};
  wire [3:0] _17877 = {_0, _17875} + {_0, _0, _17876};
  wire _17878 = _12301 < _17877;
  wire _17879 = r1428 ^ _17878;
  wire _17880 = _12298 ? coded_block[1428] : r1428;
  wire _17881 = _12296 ? _17879 : _17880;
  always @ (posedge reset or posedge clock) if (reset) r1428 <= 1'd0; else if (_12300) r1428 <= _17881;
  wire [1:0] _17882 = {_0, _672} + {_0, _3836};
  wire [1:0] _17883 = {_0, _4415} + {_0, _7548};
  wire [2:0] _17884 = {_0, _17882} + {_0, _17883};
  wire [1:0] _17885 = {_0, _9917} + {_0, _10399};
  wire [3:0] _17886 = {_0, _17884} + {_0, _0, _17885};
  wire _17887 = _12301 < _17886;
  wire _17888 = r1427 ^ _17887;
  wire _17889 = _12298 ? coded_block[1427] : r1427;
  wire _17890 = _12296 ? _17888 : _17889;
  always @ (posedge reset or posedge clock) if (reset) r1427 <= 1'd0; else if (_12300) r1427 <= _17890;
  wire [1:0] _17891 = {_0, _703} + {_0, _2813};
  wire [1:0] _17892 = {_0, _5918} + {_0, _6494};
  wire [2:0] _17893 = {_0, _17891} + {_0, _17892};
  wire [1:0] _17894 = {_0, _9630} + {_0, _11996};
  wire [3:0] _17895 = {_0, _17893} + {_0, _0, _17894};
  wire _17896 = _12301 < _17895;
  wire _17897 = r1426 ^ _17896;
  wire _17898 = _12298 ? coded_block[1426] : r1426;
  wire _17899 = _12296 ? _17897 : _17898;
  always @ (posedge reset or posedge clock) if (reset) r1426 <= 1'd0; else if (_12300) r1426 <= _17899;
  wire [1:0] _17900 = {_0, _703} + {_0, _2686};
  wire [1:0] _17901 = {_0, _5597} + {_0, _6908};
  wire [2:0] _17902 = {_0, _17900} + {_0, _17901};
  wire [1:0] _17903 = {_0, _10014} + {_0, _10590};
  wire [3:0] _17904 = {_0, _17902} + {_0, _0, _17903};
  wire _17905 = _12301 < _17904;
  wire _17906 = r1425 ^ _17905;
  wire _17907 = _12298 ? coded_block[1425] : r1425;
  wire _17908 = _12296 ? _17906 : _17907;
  always @ (posedge reset or posedge clock) if (reset) r1425 <= 1'd0; else if (_12300) r1425 <= _17908;
  wire [1:0] _17909 = {_0, _735} + {_0, _2208};
  wire [1:0] _17910 = {_0, _4767} + {_0, _7675};
  wire [2:0] _17911 = {_0, _17909} + {_0, _17910};
  wire [1:0] _17912 = {_0, _8991} + {_0, _12092};
  wire [3:0] _17913 = {_0, _17911} + {_0, _0, _17912};
  wire _17914 = _12301 < _17913;
  wire _17915 = r1424 ^ _17914;
  wire _17916 = _12298 ? coded_block[1424] : r1424;
  wire _17917 = _12296 ? _17915 : _17916;
  always @ (posedge reset or posedge clock) if (reset) r1424 <= 1'd0; else if (_12300) r1424 <= _17917;
  wire [1:0] _17918 = {_0, _766} + {_0, _2336};
  wire [1:0] _17919 = {_0, _4287} + {_0, _6845};
  wire [2:0] _17920 = {_0, _17918} + {_0, _17919};
  wire [1:0] _17921 = {_0, _9759} + {_0, _11069};
  wire [3:0] _17922 = {_0, _17920} + {_0, _0, _17921};
  wire _17923 = _12301 < _17922;
  wire _17924 = r1423 ^ _17923;
  wire _17925 = _12298 ? coded_block[1423] : r1423;
  wire _17926 = _12296 ? _17924 : _17925;
  always @ (posedge reset or posedge clock) if (reset) r1423 <= 1'd0; else if (_12300) r1423 <= _17926;
  wire [1:0] _17927 = {_0, _800} + {_0, _3678};
  wire [1:0] _17928 = {_0, _4415} + {_0, _6366};
  wire [2:0] _17929 = {_0, _17927} + {_0, _17928};
  wire [1:0] _17930 = {_0, _8926} + {_0, _11837};
  wire [3:0] _17931 = {_0, _17929} + {_0, _0, _17930};
  wire _17932 = _12301 < _17931;
  wire _17933 = r1422 ^ _17932;
  wire _17934 = _12298 ? coded_block[1422] : r1422;
  wire _17935 = _12296 ? _17933 : _17934;
  always @ (posedge reset or posedge clock) if (reset) r1422 <= 1'd0; else if (_12300) r1422 <= _17935;
  wire [1:0] _17936 = {_0, _863} + {_0, _2878};
  wire [1:0] _17937 = {_0, _4989} + {_0, _7837};
  wire [2:0] _17938 = {_0, _17936} + {_0, _17937};
  wire [1:0] _17939 = {_0, _8574} + {_0, _10527};
  wire [3:0] _17940 = {_0, _17938} + {_0, _0, _17939};
  wire _17941 = _12301 < _17940;
  wire _17942 = r1421 ^ _17941;
  wire _17943 = _12298 ? coded_block[1421] : r1421;
  wire _17944 = _12296 ? _17942 : _17943;
  always @ (posedge reset or posedge clock) if (reset) r1421 <= 1'd0; else if (_12300) r1421 <= _17944;
  wire [1:0] _17945 = {_0, _894} + {_0, _3709};
  wire [1:0] _17946 = {_0, _4958} + {_0, _7069};
  wire [2:0] _17947 = {_0, _17945} + {_0, _17946};
  wire [1:0] _17948 = {_0, _9917} + {_0, _10654};
  wire [3:0] _17949 = {_0, _17947} + {_0, _0, _17948};
  wire _17950 = _12301 < _17949;
  wire _17951 = r1420 ^ _17950;
  wire _17952 = _12298 ? coded_block[1420] : r1420;
  wire _17953 = _12296 ? _17951 : _17952;
  always @ (posedge reset or posedge clock) if (reset) r1420 <= 1'd0; else if (_12300) r1420 <= _17953;
  wire [1:0] _17954 = {_0, _927} + {_0, _3997};
  wire [1:0] _17955 = {_0, _5790} + {_0, _7036};
  wire [2:0] _17956 = {_0, _17954} + {_0, _17955};
  wire [1:0] _17957 = {_0, _9149} + {_0, _11996};
  wire [3:0] _17958 = {_0, _17956} + {_0, _0, _17957};
  wire _17959 = _12301 < _17958;
  wire _17960 = r1419 ^ _17959;
  wire _17961 = _12298 ? coded_block[1419] : r1419;
  wire _17962 = _12296 ? _17960 : _17961;
  always @ (posedge reset or posedge clock) if (reset) r1419 <= 1'd0; else if (_12300) r1419 <= _17962;
  wire [1:0] _17963 = {_0, _958} + {_0, _3390};
  wire [1:0] _17964 = {_0, _6076} + {_0, _7868};
  wire [2:0] _17965 = {_0, _17963} + {_0, _17964};
  wire [1:0] _17966 = {_0, _9118} + {_0, _11228};
  wire [3:0] _17967 = {_0, _17965} + {_0, _0, _17966};
  wire _17968 = _12301 < _17967;
  wire _17969 = r1418 ^ _17968;
  wire _17970 = _12298 ? coded_block[1418] : r1418;
  wire _17971 = _12296 ? _17969 : _17970;
  always @ (posedge reset or posedge clock) if (reset) r1418 <= 1'd0; else if (_12300) r1418 <= _17971;
  wire [1:0] _17972 = {_0, _990} + {_0, _3231};
  wire [1:0] _17973 = {_0, _5470} + {_0, _8155};
  wire [2:0] _17974 = {_0, _17972} + {_0, _17973};
  wire [1:0] _17975 = {_0, _9949} + {_0, _11196};
  wire [3:0] _17976 = {_0, _17974} + {_0, _0, _17975};
  wire _17977 = _12301 < _17976;
  wire _17978 = r1417 ^ _17977;
  wire _17979 = _12298 ? coded_block[1417] : r1417;
  wire _17980 = _12296 ? _17978 : _17979;
  always @ (posedge reset or posedge clock) if (reset) r1417 <= 1'd0; else if (_12300) r1417 <= _17980;
  wire [1:0] _17981 = {_0, _1021} + {_0, _2081};
  wire [1:0] _17982 = {_0, _5310} + {_0, _7548};
  wire [2:0] _17983 = {_0, _17981} + {_0, _17982};
  wire [1:0] _17984 = {_0, _10235} + {_0, _12027};
  wire [3:0] _17985 = {_0, _17983} + {_0, _0, _17984};
  wire _17986 = _12301 < _17985;
  wire _17987 = r1416 ^ _17986;
  wire _17988 = _12298 ? coded_block[1416] : r1416;
  wire _17989 = _12296 ? _17987 : _17988;
  always @ (posedge reset or posedge clock) if (reset) r1416 <= 1'd0; else if (_12300) r1416 <= _17989;
  wire [1:0] _17990 = {_0, _1088} + {_0, _3453};
  wire [1:0] _17991 = {_0, _5342} + {_0, _6176};
  wire [2:0] _17992 = {_0, _17990} + {_0, _17991};
  wire [1:0] _17993 = {_0, _9469} + {_0, _11708};
  wire [3:0] _17994 = {_0, _17992} + {_0, _0, _17993};
  wire _17995 = _12301 < _17994;
  wire _17996 = r1415 ^ _17995;
  wire _17997 = _12298 ? coded_block[1415] : r1415;
  wire _17998 = _12296 ? _17996 : _17997;
  always @ (posedge reset or posedge clock) if (reset) r1415 <= 1'd0; else if (_12300) r1415 <= _17998;
  wire [1:0] _17999 = {_0, _1120} + {_0, _4091};
  wire [1:0] _18000 = {_0, _5534} + {_0, _7420};
  wire [2:0] _18001 = {_0, _17999} + {_0, _18000};
  wire [1:0] _18002 = {_0, _8225} + {_0, _11550};
  wire [3:0] _18003 = {_0, _18001} + {_0, _0, _18002};
  wire _18004 = _12301 < _18003;
  wire _18005 = r1414 ^ _18004;
  wire _18006 = _12298 ? coded_block[1414] : r1414;
  wire _18007 = _12296 ? _18005 : _18006;
  always @ (posedge reset or posedge clock) if (reset) r1414 <= 1'd0; else if (_12300) r1414 <= _18007;
  wire [1:0] _18008 = {_0, _1151} + {_0, _3836};
  wire [1:0] _18009 = {_0, _4160} + {_0, _7612};
  wire [2:0] _18010 = {_0, _18008} + {_0, _18009};
  wire [1:0] _18011 = {_0, _9503} + {_0, _10272};
  wire [3:0] _18012 = {_0, _18010} + {_0, _0, _18011};
  wire _18013 = _12301 < _18012;
  wire _18014 = r1413 ^ _18013;
  wire _18015 = _12298 ? coded_block[1413] : r1413;
  wire _18016 = _12296 ? _18014 : _18015;
  always @ (posedge reset or posedge clock) if (reset) r1413 <= 1'd0; else if (_12300) r1413 <= _18016;
  wire [1:0] _18017 = {_0, _1184} + {_0, _3037};
  wire [1:0] _18018 = {_0, _5918} + {_0, _6239};
  wire [2:0] _18019 = {_0, _18017} + {_0, _18018};
  wire [1:0] _18020 = {_0, _9693} + {_0, _11581};
  wire [3:0] _18021 = {_0, _18019} + {_0, _0, _18020};
  wire _18022 = _12301 < _18021;
  wire _18023 = r1412 ^ _18022;
  wire _18024 = _12298 ? coded_block[1412] : r1412;
  wire _18025 = _12296 ? _18023 : _18024;
  always @ (posedge reset or posedge clock) if (reset) r1412 <= 1'd0; else if (_12300) r1412 <= _18025;
  wire [1:0] _18026 = {_0, _1247} + {_0, _3901};
  wire [1:0] _18027 = {_0, _5183} + {_0, _7199};
  wire [2:0] _18028 = {_0, _18026} + {_0, _18027};
  wire [1:0] _18029 = {_0, _10077} + {_0, _10399};
  wire [3:0] _18030 = {_0, _18028} + {_0, _0, _18029};
  wire _18031 = _12301 < _18030;
  wire _18032 = r1411 ^ _18031;
  wire _18033 = _12298 ? coded_block[1411] : r1411;
  wire _18034 = _12296 ? _18032 : _18033;
  always @ (posedge reset or posedge clock) if (reset) r1411 <= 1'd0; else if (_12300) r1411 <= _18034;
  wire [1:0] _18035 = {_0, _1278} + {_0, _2592};
  wire [1:0] _18036 = {_0, _5981} + {_0, _7262};
  wire [2:0] _18037 = {_0, _18035} + {_0, _18036};
  wire [1:0] _18038 = {_0, _9279} + {_0, _12155};
  wire [3:0] _18039 = {_0, _18037} + {_0, _0, _18038};
  wire _18040 = _12301 < _18039;
  wire _18041 = r1410 ^ _18040;
  wire _18042 = _12298 ? coded_block[1410] : r1410;
  wire _18043 = _12296 ? _18041 : _18042;
  always @ (posedge reset or posedge clock) if (reset) r1410 <= 1'd0; else if (_12300) r1410 <= _18043;
  wire [1:0] _18044 = {_0, _1312} + {_0, _2494};
  wire [1:0] _18045 = {_0, _4671} + {_0, _8059};
  wire [2:0] _18046 = {_0, _18044} + {_0, _18045};
  wire [1:0] _18047 = {_0, _9342} + {_0, _11358};
  wire [3:0] _18048 = {_0, _18046} + {_0, _0, _18047};
  wire _18049 = _12301 < _18048;
  wire _18050 = r1409 ^ _18049;
  wire _18051 = _12298 ? coded_block[1409] : r1409;
  wire _18052 = _12296 ? _18050 : _18051;
  always @ (posedge reset or posedge clock) if (reset) r1409 <= 1'd0; else if (_12300) r1409 <= _18052;
  wire [1:0] _18053 = {_0, _1343} + {_0, _3005};
  wire [1:0] _18054 = {_0, _4574} + {_0, _6750};
  wire [2:0] _18055 = {_0, _18053} + {_0, _18054};
  wire [1:0] _18056 = {_0, _10141} + {_0, _11422};
  wire [3:0] _18057 = {_0, _18055} + {_0, _0, _18056};
  wire _18058 = _12301 < _18057;
  wire _18059 = r1408 ^ _18058;
  wire _18060 = _12298 ? coded_block[1408] : r1408;
  wire _18061 = _12296 ? _18059 : _18060;
  always @ (posedge reset or posedge clock) if (reset) r1408 <= 1'd0; else if (_12300) r1408 <= _18061;
  wire [1:0] _18062 = {_0, _1375} + {_0, _3870};
  wire [1:0] _18063 = {_0, _5085} + {_0, _6652};
  wire [2:0] _18064 = {_0, _18062} + {_0, _18063};
  wire [1:0] _18065 = {_0, _8830} + {_0, _12219};
  wire [3:0] _18066 = {_0, _18064} + {_0, _0, _18065};
  wire _18067 = _12301 < _18066;
  wire _18068 = r1407 ^ _18067;
  wire _18069 = _12298 ? coded_block[1407] : r1407;
  wire _18070 = _12296 ? _18068 : _18069;
  always @ (posedge reset or posedge clock) if (reset) r1407 <= 1'd0; else if (_12300) r1407 <= _18070;
  wire [1:0] _18071 = {_0, _1406} + {_0, _3135};
  wire [1:0] _18072 = {_0, _5949} + {_0, _7163};
  wire [2:0] _18073 = {_0, _18071} + {_0, _18072};
  wire [1:0] _18074 = {_0, _8736} + {_0, _10910};
  wire [3:0] _18075 = {_0, _18073} + {_0, _0, _18074};
  wire _18076 = _12301 < _18075;
  wire _18077 = r1406 ^ _18076;
  wire _18078 = _12298 ? coded_block[1406] : r1406;
  wire _18079 = _12296 ? _18077 : _18078;
  always @ (posedge reset or posedge clock) if (reset) r1406 <= 1'd0; else if (_12300) r1406 <= _18079;
  wire [1:0] _18080 = {_0, _1439} + {_0, _2175};
  wire [1:0] _18081 = {_0, _5215} + {_0, _8028};
  wire [2:0] _18082 = {_0, _18080} + {_0, _18081};
  wire [1:0] _18083 = {_0, _9248} + {_0, _10814};
  wire [3:0] _18084 = {_0, _18082} + {_0, _0, _18083};
  wire _18085 = _12301 < _18084;
  wire _18086 = r1405 ^ _18085;
  wire _18087 = _12298 ? coded_block[1405] : r1405;
  wire _18088 = _12296 ? _18086 : _18087;
  always @ (posedge reset or posedge clock) if (reset) r1405 <= 1'd0; else if (_12300) r1405 <= _18088;
  wire [1:0] _18089 = {_0, _1470} + {_0, _2719};
  wire [1:0] _18090 = {_0, _4256} + {_0, _7293};
  wire [2:0] _18091 = {_0, _18089} + {_0, _18090};
  wire [1:0] _18092 = {_0, _10108} + {_0, _11326};
  wire [3:0] _18093 = {_0, _18091} + {_0, _0, _18092};
  wire _18094 = _12301 < _18093;
  wire _18095 = r1404 ^ _18094;
  wire _18096 = _12298 ? coded_block[1404] : r1404;
  wire _18097 = _12296 ? _18095 : _18096;
  always @ (posedge reset or posedge clock) if (reset) r1404 <= 1'd0; else if (_12300) r1404 <= _18097;
  wire [1:0] _18098 = {_0, _1502} + {_0, _3805};
  wire [1:0] _18099 = {_0, _4798} + {_0, _6334};
  wire [2:0] _18100 = {_0, _18098} + {_0, _18099};
  wire [1:0] _18101 = {_0, _9375} + {_0, _12188};
  wire [3:0] _18102 = {_0, _18100} + {_0, _0, _18101};
  wire _18103 = _12301 < _18102;
  wire _18104 = r1403 ^ _18103;
  wire _18105 = _12298 ? coded_block[1403] : r1403;
  wire _18106 = _12296 ? _18104 : _18105;
  always @ (posedge reset or posedge clock) if (reset) r1403 <= 1'd0; else if (_12300) r1403 <= _18106;
  wire [1:0] _18107 = {_0, _1533} + {_0, _2112};
  wire [1:0] _18108 = {_0, _5884} + {_0, _6877};
  wire [2:0] _18109 = {_0, _18107} + {_0, _18108};
  wire [1:0] _18110 = {_0, _8415} + {_0, _11453};
  wire [3:0] _18111 = {_0, _18109} + {_0, _0, _18110};
  wire _18112 = _12301 < _18111;
  wire _18113 = r1402 ^ _18112;
  wire _18114 = _12298 ? coded_block[1402] : r1402;
  wire _18115 = _12296 ? _18113 : _18114;
  always @ (posedge reset or posedge clock) if (reset) r1402 <= 1'd0; else if (_12300) r1402 <= _18115;
  wire [1:0] _18116 = {_0, _1568} + {_0, _2557};
  wire [1:0] _18117 = {_0, _4192} + {_0, _7965};
  wire [2:0] _18118 = {_0, _18116} + {_0, _18117};
  wire [1:0] _18119 = {_0, _8957} + {_0, _10493};
  wire [3:0] _18120 = {_0, _18118} + {_0, _0, _18119};
  wire _18121 = _12301 < _18120;
  wire _18122 = r1401 ^ _18121;
  wire _18123 = _12298 ? coded_block[1401] : r1401;
  wire _18124 = _12296 ? _18122 : _18123;
  always @ (posedge reset or posedge clock) if (reset) r1401 <= 1'd0; else if (_12300) r1401 <= _18124;
  wire [1:0] _18125 = {_0, _1599} + {_0, _3933};
  wire [1:0] _18126 = {_0, _4640} + {_0, _6270};
  wire [2:0] _18127 = {_0, _18125} + {_0, _18126};
  wire [1:0] _18128 = {_0, _10045} + {_0, _11038};
  wire [3:0] _18129 = {_0, _18127} + {_0, _0, _18128};
  wire _18130 = _12301 < _18129;
  wire _18131 = r1400 ^ _18130;
  wire _18132 = _12298 ? coded_block[1400] : r1400;
  wire _18133 = _12296 ? _18131 : _18132;
  always @ (posedge reset or posedge clock) if (reset) r1400 <= 1'd0; else if (_12300) r1400 <= _18133;
  wire [1:0] _18134 = {_0, _1631} + {_0, _2847};
  wire [1:0] _18135 = {_0, _6012} + {_0, _6718};
  wire [2:0] _18136 = {_0, _18134} + {_0, _18135};
  wire [1:0] _18137 = {_0, _8352} + {_0, _12124};
  wire [3:0] _18138 = {_0, _18136} + {_0, _0, _18137};
  wire _18139 = _12301 < _18138;
  wire _18140 = r1399 ^ _18139;
  wire _18141 = _12298 ? coded_block[1399] : r1399;
  wire _18142 = _12296 ? _18140 : _18141;
  always @ (posedge reset or posedge clock) if (reset) r1399 <= 1'd0; else if (_12300) r1399 <= _18142;
  wire [1:0] _18143 = {_0, _1662} + {_0, _2941};
  wire [1:0] _18144 = {_0, _4926} + {_0, _8092};
  wire [2:0] _18145 = {_0, _18143} + {_0, _18144};
  wire [1:0] _18146 = {_0, _8799} + {_0, _10430};
  wire [3:0] _18147 = {_0, _18145} + {_0, _0, _18146};
  wire _18148 = _12301 < _18147;
  wire _18149 = r1398 ^ _18148;
  wire _18150 = _12298 ? coded_block[1398] : r1398;
  wire _18151 = _12296 ? _18149 : _18150;
  always @ (posedge reset or posedge clock) if (reset) r1398 <= 1'd0; else if (_12300) r1398 <= _18151;
  wire [1:0] _18152 = {_0, _1695} + {_0, _2399};
  wire [1:0] _18153 = {_0, _5022} + {_0, _7005};
  wire [2:0] _18154 = {_0, _18152} + {_0, _18153};
  wire [1:0] _18155 = {_0, _10172} + {_0, _10877};
  wire [3:0] _18156 = {_0, _18154} + {_0, _0, _18155};
  wire _18157 = _12301 < _18156;
  wire _18158 = r1397 ^ _18157;
  wire _18159 = _12298 ? coded_block[1397] : r1397;
  wire _18160 = _12296 ? _18158 : _18159;
  always @ (posedge reset or posedge clock) if (reset) r1397 <= 1'd0; else if (_12300) r1397 <= _18160;
  wire [1:0] _18161 = {_0, _1726} + {_0, _2655};
  wire [1:0] _18162 = {_0, _4478} + {_0, _7100};
  wire [2:0] _18163 = {_0, _18161} + {_0, _18162};
  wire [1:0] _18164 = {_0, _9085} + {_0, _12251};
  wire [3:0] _18165 = {_0, _18163} + {_0, _0, _18164};
  wire _18166 = _12301 < _18165;
  wire _18167 = r1396 ^ _18166;
  wire _18168 = _12298 ? coded_block[1396] : r1396;
  wire _18169 = _12296 ? _18167 : _18168;
  always @ (posedge reset or posedge clock) if (reset) r1396 <= 1'd0; else if (_12300) r1396 <= _18169;
  wire [1:0] _18170 = {_0, _1789} + {_0, _3198};
  wire [1:0] _18171 = {_0, _5628} + {_0, _6814};
  wire [2:0] _18172 = {_0, _18170} + {_0, _18171};
  wire [1:0] _18173 = {_0, _8638} + {_0, _11259};
  wire [3:0] _18174 = {_0, _18172} + {_0, _0, _18173};
  wire _18175 = _12301 < _18174;
  wire _18176 = r1395 ^ _18175;
  wire _18177 = _12298 ? coded_block[1395] : r1395;
  wire _18178 = _12296 ? _18176 : _18177;
  always @ (posedge reset or posedge clock) if (reset) r1395 <= 1'd0; else if (_12300) r1395 <= _18178;
  wire [1:0] _18179 = {_0, _1823} + {_0, _3422};
  wire [1:0] _18180 = {_0, _5279} + {_0, _7710};
  wire [2:0] _18181 = {_0, _18179} + {_0, _18180};
  wire [1:0] _18182 = {_0, _8894} + {_0, _10717};
  wire [3:0] _18183 = {_0, _18181} + {_0, _0, _18182};
  wire _18184 = _12301 < _18183;
  wire _18185 = r1394 ^ _18184;
  wire _18186 = _12298 ? coded_block[1394] : r1394;
  wire _18187 = _12296 ? _18185 : _18186;
  always @ (posedge reset or posedge clock) if (reset) r1394 <= 1'd0; else if (_12300) r1394 <= _18187;
  wire [1:0] _18188 = {_0, _1886} + {_0, _3646};
  wire [1:0] _18189 = {_0, _5373} + {_0, _7581};
  wire [2:0] _18190 = {_0, _18188} + {_0, _18189};
  wire [1:0] _18191 = {_0, _9438} + {_0, _11869};
  wire [3:0] _18192 = {_0, _18190} + {_0, _0, _18191};
  wire _18193 = _12301 < _18192;
  wire _18194 = r1393 ^ _18193;
  wire _18195 = _12298 ? coded_block[1393] : r1393;
  wire _18196 = _12296 ? _18194 : _18195;
  always @ (posedge reset or posedge clock) if (reset) r1393 <= 1'd0; else if (_12300) r1393 <= _18196;
  wire [1:0] _18197 = {_0, _1981} + {_0, _2526};
  wire [1:0] _18198 = {_0, _5053} + {_0, _6525};
  wire [2:0] _18199 = {_0, _18197} + {_0, _18198};
  wire [1:0] _18200 = {_0, _9886} + {_0, _11613};
  wire [3:0] _18201 = {_0, _18199} + {_0, _0, _18200};
  wire _18202 = _12301 < _18201;
  wire _18203 = r1392 ^ _18202;
  wire _18204 = _12298 ? coded_block[1392] : r1392;
  wire _18205 = _12296 ? _18203 : _18204;
  always @ (posedge reset or posedge clock) if (reset) r1392 <= 1'd0; else if (_12300) r1392 <= _18205;
  wire [1:0] _18206 = {_0, _2013} + {_0, _2144};
  wire [1:0] _18207 = {_0, _4605} + {_0, _7132};
  wire [2:0] _18208 = {_0, _18206} + {_0, _18207};
  wire [1:0] _18209 = {_0, _8607} + {_0, _11964};
  wire [3:0] _18210 = {_0, _18208} + {_0, _0, _18209};
  wire _18211 = _12301 < _18210;
  wire _18212 = r1391 ^ _18211;
  wire _18213 = _12298 ? coded_block[1391] : r1391;
  wire _18214 = _12296 ? _18212 : _18213;
  always @ (posedge reset or posedge clock) if (reset) r1391 <= 1'd0; else if (_12300) r1391 <= _18214;
  wire [1:0] _18215 = {_0, _735} + {_0, _3580};
  wire [1:0] _18216 = {_0, _4895} + {_0, _7996};
  wire [2:0] _18217 = {_0, _18215} + {_0, _18216};
  wire [1:0] _18218 = {_0, _8574} + {_0, _11708};
  wire [3:0] _18219 = {_0, _18217} + {_0, _0, _18218};
  wire _18220 = _12301 < _18219;
  wire _18221 = r1390 ^ _18220;
  wire _18222 = _12298 ? coded_block[1390] : r1390;
  wire _18223 = _12296 ? _18221 : _18222;
  always @ (posedge reset or posedge clock) if (reset) r1390 <= 1'd0; else if (_12300) r1390 <= _18223;
  wire [1:0] _18224 = {_0, _766} + {_0, _2750};
  wire [1:0] _18225 = {_0, _5663} + {_0, _6973};
  wire [2:0] _18226 = {_0, _18224} + {_0, _18225};
  wire [1:0] _18227 = {_0, _10077} + {_0, _10654};
  wire [3:0] _18228 = {_0, _18226} + {_0, _0, _18227};
  wire _18229 = _12301 < _18228;
  wire _18230 = r1389 ^ _18229;
  wire _18231 = _12298 ? coded_block[1389] : r1389;
  wire _18232 = _12296 ? _18230 : _18231;
  always @ (posedge reset or posedge clock) if (reset) r1389 <= 1'd0; else if (_12300) r1389 <= _18232;
  wire [1:0] _18233 = {_0, _800} + {_0, _2271};
  wire [1:0] _18234 = {_0, _4830} + {_0, _7741};
  wire [2:0] _18235 = {_0, _18233} + {_0, _18234};
  wire [1:0] _18236 = {_0, _9054} + {_0, _12155};
  wire [3:0] _18237 = {_0, _18235} + {_0, _0, _18236};
  wire _18238 = _12301 < _18237;
  wire _18239 = r1388 ^ _18238;
  wire _18240 = _12298 ? coded_block[1388] : r1388;
  wire _18241 = _12296 ? _18239 : _18240;
  always @ (posedge reset or posedge clock) if (reset) r1388 <= 1'd0; else if (_12300) r1388 <= _18241;
  wire [1:0] _18242 = {_0, _831} + {_0, _2399};
  wire [1:0] _18243 = {_0, _4350} + {_0, _6908};
  wire [2:0] _18244 = {_0, _18242} + {_0, _18243};
  wire [1:0] _18245 = {_0, _9822} + {_0, _11132};
  wire [3:0] _18246 = {_0, _18244} + {_0, _0, _18245};
  wire _18247 = _12301 < _18246;
  wire _18248 = r1387 ^ _18247;
  wire _18249 = _12298 ? coded_block[1387] : r1387;
  wire _18250 = _12296 ? _18248 : _18249;
  always @ (posedge reset or posedge clock) if (reset) r1387 <= 1'd0; else if (_12300) r1387 <= _18250;
  wire [1:0] _18251 = {_0, _863} + {_0, _3742};
  wire [1:0] _18252 = {_0, _4478} + {_0, _6431};
  wire [2:0] _18253 = {_0, _18251} + {_0, _18252};
  wire [1:0] _18254 = {_0, _8991} + {_0, _11900};
  wire [3:0] _18255 = {_0, _18253} + {_0, _0, _18254};
  wire _18256 = _12301 < _18255;
  wire _18257 = r1386 ^ _18256;
  wire _18258 = _12298 ? coded_block[1386] : r1386;
  wire _18259 = _12296 ? _18257 : _18258;
  always @ (posedge reset or posedge clock) if (reset) r1386 <= 1'd0; else if (_12300) r1386 <= _18259;
  wire [1:0] _18260 = {_0, _894} + {_0, _2974};
  wire [1:0] _18261 = {_0, _5821} + {_0, _6558};
  wire [2:0] _18262 = {_0, _18260} + {_0, _18261};
  wire [1:0] _18263 = {_0, _8511} + {_0, _11069};
  wire [3:0] _18264 = {_0, _18262} + {_0, _0, _18263};
  wire _18265 = _12301 < _18264;
  wire _18266 = r1385 ^ _18265;
  wire _18267 = _12298 ? coded_block[1385] : r1385;
  wire _18268 = _12296 ? _18266 : _18267;
  always @ (posedge reset or posedge clock) if (reset) r1385 <= 1'd0; else if (_12300) r1385 <= _18268;
  wire [1:0] _18269 = {_0, _927} + {_0, _2941};
  wire [1:0] _18270 = {_0, _5053} + {_0, _7900};
  wire [2:0] _18271 = {_0, _18269} + {_0, _18270};
  wire [1:0] _18272 = {_0, _8638} + {_0, _10590};
  wire [3:0] _18273 = {_0, _18271} + {_0, _0, _18272};
  wire _18274 = _12301 < _18273;
  wire _18275 = r1384 ^ _18274;
  wire _18276 = _12298 ? coded_block[1384] : r1384;
  wire _18277 = _12296 ? _18275 : _18276;
  always @ (posedge reset or posedge clock) if (reset) r1384 <= 1'd0; else if (_12300) r1384 <= _18277;
  wire [1:0] _18278 = {_0, _192} + {_0, _2910};
  wire [1:0] _18279 = {_0, _5534} + {_0, _7517};
  wire [2:0] _18280 = {_0, _18278} + {_0, _18279};
  wire [1:0] _18281 = {_0, _8670} + {_0, _11389};
  wire [3:0] _18282 = {_0, _18280} + {_0, _0, _18281};
  wire _18283 = _12301 < _18282;
  wire _18284 = r1383 ^ _18283;
  wire _18285 = _12298 ? coded_block[1383] : r1383;
  wire _18286 = _12296 ? _18284 : _18285;
  always @ (posedge reset or posedge clock) if (reset) r1383 <= 1'd0; else if (_12300) r1383 <= _18286;
  wire [1:0] _18287 = {_0, _224} + {_0, _3167};
  wire [1:0] _18288 = {_0, _4989} + {_0, _7612};
  wire [2:0] _18289 = {_0, _18287} + {_0, _18288};
  wire [1:0] _18290 = {_0, _9597} + {_0, _10748};
  wire [3:0] _18291 = {_0, _18289} + {_0, _0, _18290};
  wire _18292 = _12301 < _18291;
  wire _18293 = r1382 ^ _18292;
  wire _18294 = _12298 ? coded_block[1382] : r1382;
  wire _18295 = _12296 ? _18293 : _18294;
  always @ (posedge reset or posedge clock) if (reset) r1382 <= 1'd0; else if (_12300) r1382 <= _18295;
  wire [1:0] _18296 = {_0, _255} + {_0, _4060};
  wire [1:0] _18297 = {_0, _5246} + {_0, _7069};
  wire [2:0] _18298 = {_0, _18296} + {_0, _18297};
  wire [1:0] _18299 = {_0, _9693} + {_0, _11677};
  wire [3:0] _18300 = {_0, _18298} + {_0, _0, _18299};
  wire _18301 = _12301 < _18300;
  wire _18302 = r1381 ^ _18301;
  wire _18303 = _12298 ? coded_block[1381] : r1381;
  wire _18304 = _12296 ? _18302 : _18303;
  always @ (posedge reset or posedge clock) if (reset) r1381 <= 1'd0; else if (_12300) r1381 <= _18304;
  wire [1:0] _18305 = {_0, _289} + {_0, _3709};
  wire [1:0] _18306 = {_0, _6139} + {_0, _7326};
  wire [2:0] _18307 = {_0, _18305} + {_0, _18306};
  wire [1:0] _18308 = {_0, _9149} + {_0, _11771};
  wire [3:0] _18309 = {_0, _18307} + {_0, _0, _18308};
  wire _18310 = _12301 < _18309;
  wire _18311 = r1380 ^ _18310;
  wire _18312 = _12298 ? coded_block[1380] : r1380;
  wire _18313 = _12296 ? _18311 : _18312;
  always @ (posedge reset or posedge clock) if (reset) r1380 <= 1'd0; else if (_12300) r1380 <= _18313;
  wire [1:0] _18314 = {_0, _320} + {_0, _3933};
  wire [1:0] _18315 = {_0, _5790} + {_0, _6207};
  wire [2:0] _18316 = {_0, _18314} + {_0, _18315};
  wire [1:0] _18317 = {_0, _9406} + {_0, _11228};
  wire [3:0] _18318 = {_0, _18316} + {_0, _0, _18317};
  wire _18319 = _12301 < _18318;
  wire _18320 = r1379 ^ _18319;
  wire _18321 = _12298 ? coded_block[1379] : r1379;
  wire _18322 = _12296 ? _18320 : _18321;
  always @ (posedge reset or posedge clock) if (reset) r1379 <= 1'd0; else if (_12300) r1379 <= _18322;
  wire [1:0] _18323 = {_0, _352} + {_0, _3805};
  wire [1:0] _18324 = {_0, _6012} + {_0, _7868};
  wire [2:0] _18325 = {_0, _18323} + {_0, _18324};
  wire [1:0] _18326 = {_0, _8288} + {_0, _11485};
  wire [3:0] _18327 = {_0, _18325} + {_0, _0, _18326};
  wire _18328 = _12301 < _18327;
  wire _18329 = r1378 ^ _18328;
  wire _18330 = _12298 ? coded_block[1378] : r1378;
  wire _18331 = _12296 ? _18329 : _18330;
  always @ (posedge reset or posedge clock) if (reset) r1378 <= 1'd0; else if (_12300) r1378 <= _18331;
  wire [1:0] _18332 = {_0, _416} + {_0, _2878};
  wire [1:0] _18333 = {_0, _4223} + {_0, _7965};
  wire [2:0] _18334 = {_0, _18332} + {_0, _18333};
  wire [1:0] _18335 = {_0, _10172} + {_0, _12027};
  wire [3:0] _18336 = {_0, _18334} + {_0, _0, _18335};
  wire _18337 = _12301 < _18336;
  wire _18338 = r1377 ^ _18337;
  wire _18339 = _12298 ? coded_block[1377] : r1377;
  wire _18340 = _12296 ? _18338 : _18339;
  always @ (posedge reset or posedge clock) if (reset) r1377 <= 1'd0; else if (_12300) r1377 <= _18340;
  wire [1:0] _18341 = {_0, _447} + {_0, _3486};
  wire [1:0] _18342 = {_0, _4958} + {_0, _6303};
  wire [2:0] _18343 = {_0, _18341} + {_0, _18342};
  wire [1:0] _18344 = {_0, _10045} + {_0, _12251};
  wire [3:0] _18345 = {_0, _18343} + {_0, _0, _18344};
  wire _18346 = _12301 < _18345;
  wire _18347 = r1376 ^ _18346;
  wire _18348 = _12298 ? coded_block[1376] : r1376;
  wire _18349 = _12296 ? _18347 : _18348;
  always @ (posedge reset or posedge clock) if (reset) r1376 <= 1'd0; else if (_12300) r1376 <= _18349;
  wire [1:0] _18350 = {_0, _479} + {_0, _3037};
  wire [1:0] _18351 = {_0, _5565} + {_0, _7036};
  wire [2:0] _18352 = {_0, _18350} + {_0, _18351};
  wire [1:0] _18353 = {_0, _8383} + {_0, _12124};
  wire [3:0] _18354 = {_0, _18352} + {_0, _0, _18353};
  wire _18355 = _12301 < _18354;
  wire _18356 = r1375 ^ _18355;
  wire _18357 = _12298 ? coded_block[1375] : r1375;
  wire _18358 = _12296 ? _18356 : _18357;
  always @ (posedge reset or posedge clock) if (reset) r1375 <= 1'd0; else if (_12300) r1375 <= _18358;
  wire [1:0] _18359 = {_0, _510} + {_0, _2655};
  wire [1:0] _18360 = {_0, _5116} + {_0, _7644};
  wire [2:0] _18361 = {_0, _18359} + {_0, _18360};
  wire [1:0] _18362 = {_0, _9118} + {_0, _10462};
  wire [3:0] _18363 = {_0, _18361} + {_0, _0, _18362};
  wire _18364 = _12301 < _18363;
  wire _18365 = r1374 ^ _18364;
  wire _18366 = _12298 ? coded_block[1374] : r1374;
  wire _18367 = _12296 ? _18365 : _18366;
  always @ (posedge reset or posedge clock) if (reset) r1374 <= 1'd0; else if (_12300) r1374 <= _18367;
  wire [1:0] _18368 = {_0, _545} + {_0, _3678};
  wire [1:0] _18369 = {_0, _4734} + {_0, _7199};
  wire [2:0] _18370 = {_0, _18368} + {_0, _18369};
  wire [1:0] _18371 = {_0, _9724} + {_0, _11196};
  wire [3:0] _18372 = {_0, _18370} + {_0, _0, _18371};
  wire _18373 = _12301 < _18372;
  wire _18374 = r1373 ^ _18373;
  wire _18375 = _12298 ? coded_block[1373] : r1373;
  wire _18376 = _12296 ? _18374 : _18375;
  always @ (posedge reset or posedge clock) if (reset) r1373 <= 1'd0; else if (_12300) r1373 <= _18376;
  wire [1:0] _18377 = {_0, _576} + {_0, _4091};
  wire [1:0] _18378 = {_0, _5757} + {_0, _6814};
  wire [2:0] _18379 = {_0, _18377} + {_0, _18378};
  wire [1:0] _18380 = {_0, _9279} + {_0, _11806};
  wire [3:0] _18381 = {_0, _18379} + {_0, _0, _18380};
  wire _18382 = _12301 < _18381;
  wire _18383 = r1372 ^ _18382;
  wire _18384 = _12298 ? coded_block[1372] : r1372;
  wire _18385 = _12296 ? _18383 : _18384;
  always @ (posedge reset or posedge clock) if (reset) r1372 <= 1'd0; else if (_12300) r1372 <= _18385;
  wire [1:0] _18386 = {_0, _608} + {_0, _2557};
  wire [1:0] _18387 = {_0, _4160} + {_0, _7837};
  wire [2:0] _18388 = {_0, _18386} + {_0, _18387};
  wire [1:0] _18389 = {_0, _8894} + {_0, _11358};
  wire [3:0] _18390 = {_0, _18388} + {_0, _0, _18389};
  wire _18391 = _12301 < _18390;
  wire _18392 = r1371 ^ _18391;
  wire _18393 = _12298 ? coded_block[1371] : r1371;
  wire _18394 = _12296 ? _18392 : _18393;
  always @ (posedge reset or posedge clock) if (reset) r1371 <= 1'd0; else if (_12300) r1371 <= _18394;
  wire [1:0] _18395 = {_0, _639} + {_0, _3997};
  wire [1:0] _18396 = {_0, _4640} + {_0, _6239};
  wire [2:0] _18397 = {_0, _18395} + {_0, _18396};
  wire [1:0] _18398 = {_0, _9917} + {_0, _10973};
  wire [3:0] _18399 = {_0, _18397} + {_0, _0, _18398};
  wire _18400 = _12301 < _18399;
  wire _18401 = r1370 ^ _18400;
  wire _18402 = _12298 ? coded_block[1370] : r1370;
  wire _18403 = _12296 ? _18401 : _18402;
  always @ (posedge reset or posedge clock) if (reset) r1370 <= 1'd0; else if (_12300) r1370 <= _18403;
  wire [1:0] _18404 = {_0, _703} + {_0, _2974};
  wire [1:0] _18405 = {_0, _5373} + {_0, _8155};
  wire [2:0] _18406 = {_0, _18404} + {_0, _18405};
  wire [1:0] _18407 = {_0, _8799} + {_0, _10399};
  wire [3:0] _18408 = {_0, _18406} + {_0, _0, _18407};
  wire _18409 = _12301 < _18408;
  wire _18410 = r1369 ^ _18409;
  wire _18411 = _12298 ? coded_block[1369] : r1369;
  wire _18412 = _12296 ? _18410 : _18411;
  always @ (posedge reset or posedge clock) if (reset) r1369 <= 1'd0; else if (_12300) r1369 <= _18412;
  wire [1:0] _18413 = {_0, _735} + {_0, _3135};
  wire [1:0] _18414 = {_0, _5053} + {_0, _7454};
  wire [2:0] _18415 = {_0, _18413} + {_0, _18414};
  wire [1:0] _18416 = {_0, _10235} + {_0, _10877};
  wire [3:0] _18417 = {_0, _18415} + {_0, _0, _18416};
  wire _18418 = _12301 < _18417;
  wire _18419 = r1368 ^ _18418;
  wire _18420 = _12298 ? coded_block[1368] : r1368;
  wire _18421 = _12296 ? _18419 : _18420;
  always @ (posedge reset or posedge clock) if (reset) r1368 <= 1'd0; else if (_12300) r1368 <= _18421;
  wire [1:0] _18422 = {_0, _766} + {_0, _2941};
  wire [1:0] _18423 = {_0, _5215} + {_0, _7132};
  wire [2:0] _18424 = {_0, _18422} + {_0, _18423};
  wire [1:0] _18425 = {_0, _9534} + {_0, _10303};
  wire [3:0] _18426 = {_0, _18424} + {_0, _0, _18425};
  wire _18427 = _12301 < _18426;
  wire _18428 = r1367 ^ _18427;
  wire _18429 = _12298 ? coded_block[1367] : r1367;
  wire _18430 = _12296 ? _18428 : _18429;
  always @ (posedge reset or posedge clock) if (reset) r1367 <= 1'd0; else if (_12300) r1367 <= _18430;
  wire [1:0] _18431 = {_0, _800} + {_0, _3325};
  wire [1:0] _18432 = {_0, _5022} + {_0, _7293};
  wire [2:0] _18433 = {_0, _18431} + {_0, _18432};
  wire [1:0] _18434 = {_0, _9212} + {_0, _11613};
  wire [3:0] _18435 = {_0, _18433} + {_0, _0, _18434};
  wire _18436 = _12301 < _18435;
  wire _18437 = r1366 ^ _18436;
  wire _18438 = _12298 ? coded_block[1366] : r1366;
  wire _18439 = _12296 ? _18437 : _18438;
  always @ (posedge reset or posedge clock) if (reset) r1366 <= 1'd0; else if (_12300) r1366 <= _18439;
  wire [1:0] _18440 = {_0, _831} + {_0, _2463};
  wire [1:0] _18441 = {_0, _5407} + {_0, _7100};
  wire [2:0] _18442 = {_0, _18440} + {_0, _18441};
  wire [1:0] _18443 = {_0, _9375} + {_0, _11295};
  wire [3:0] _18444 = {_0, _18442} + {_0, _0, _18443};
  wire _18445 = _12301 < _18444;
  wire _18446 = r1365 ^ _18445;
  wire _18447 = _12298 ? coded_block[1365] : r1365;
  wire _18448 = _12296 ? _18446 : _18447;
  always @ (posedge reset or posedge clock) if (reset) r1365 <= 1'd0; else if (_12300) r1365 <= _18448;
  wire [1:0] _18449 = {_0, _863} + {_0, _2239};
  wire [1:0] _18450 = {_0, _4542} + {_0, _7485};
  wire [2:0] _18451 = {_0, _18449} + {_0, _18450};
  wire [1:0] _18452 = {_0, _9181} + {_0, _11453};
  wire [3:0] _18453 = {_0, _18451} + {_0, _0, _18452};
  wire _18454 = _12301 < _18453;
  wire _18455 = r1364 ^ _18454;
  wire _18456 = _12298 ? coded_block[1364] : r1364;
  wire _18457 = _12296 ? _18455 : _18456;
  always @ (posedge reset or posedge clock) if (reset) r1364 <= 1'd0; else if (_12300) r1364 <= _18457;
  wire [1:0] _18458 = {_0, _927} + {_0, _2750};
  wire [1:0] _18459 = {_0, _4895} + {_0, _6397};
  wire [2:0] _18460 = {_0, _18458} + {_0, _18459};
  wire [1:0] _18461 = {_0, _8701} + {_0, _11644};
  wire [3:0] _18462 = {_0, _18460} + {_0, _0, _18461};
  wire _18463 = _12301 < _18462;
  wire _18464 = r1363 ^ _18463;
  wire _18465 = _12298 ? coded_block[1363] : r1363;
  wire _18466 = _12296 ? _18464 : _18465;
  always @ (posedge reset or posedge clock) if (reset) r1363 <= 1'd0; else if (_12300) r1363 <= _18466;
  wire [1:0] _18467 = {_0, _958} + {_0, _3870};
  wire [1:0] _18468 = {_0, _4830} + {_0, _6973};
  wire [2:0] _18469 = {_0, _18467} + {_0, _18468};
  wire [1:0] _18470 = {_0, _8480} + {_0, _10783};
  wire [3:0] _18471 = {_0, _18469} + {_0, _0, _18470};
  wire _18472 = _12301 < _18471;
  wire _18473 = r1362 ^ _18472;
  wire _18474 = _12298 ? coded_block[1362] : r1362;
  wire _18475 = _12296 ? _18473 : _18474;
  always @ (posedge reset or posedge clock) if (reset) r1362 <= 1'd0; else if (_12300) r1362 <= _18475;
  wire [1:0] _18476 = {_0, _990} + {_0, _2526};
  wire [1:0] _18477 = {_0, _5949} + {_0, _6908};
  wire [2:0] _18478 = {_0, _18476} + {_0, _18477};
  wire [1:0] _18479 = {_0, _9054} + {_0, _10558};
  wire [3:0] _18480 = {_0, _18478} + {_0, _0, _18479};
  wire _18481 = _12301 < _18480;
  wire _18482 = r1361 ^ _18481;
  wire _18483 = _12298 ? coded_block[1361] : r1361;
  wire _18484 = _12296 ? _18482 : _18483;
  always @ (posedge reset or posedge clock) if (reset) r1361 <= 1'd0; else if (_12300) r1361 <= _18484;
  wire [1:0] _18485 = {_0, _1021} + {_0, _2112};
  wire [1:0] _18486 = {_0, _4605} + {_0, _8028};
  wire [2:0] _18487 = {_0, _18485} + {_0, _18486};
  wire [1:0] _18488 = {_0, _8991} + {_0, _11132};
  wire [3:0] _18489 = {_0, _18487} + {_0, _0, _18488};
  wire _18490 = _12301 < _18489;
  wire _18491 = r1360 ^ _18490;
  wire _18492 = _12298 ? coded_block[1360] : r1360;
  wire _18493 = _12296 ? _18491 : _18492;
  always @ (posedge reset or posedge clock) if (reset) r1360 <= 1'd0; else if (_12300) r1360 <= _18493;
  wire [1:0] _18494 = {_0, _1057} + {_0, _3836};
  wire [1:0] _18495 = {_0, _4192} + {_0, _6687};
  wire [2:0] _18496 = {_0, _18494} + {_0, _18495};
  wire [1:0] _18497 = {_0, _10108} + {_0, _11069};
  wire [3:0] _18498 = {_0, _18496} + {_0, _0, _18497};
  wire _18499 = _12301 < _18498;
  wire _18500 = r1359 ^ _18499;
  wire _18501 = _12298 ? coded_block[1359] : r1359;
  wire _18502 = _12296 ? _18500 : _18501;
  always @ (posedge reset or posedge clock) if (reset) r1359 <= 1'd0; else if (_12300) r1359 <= _18502;
  wire [1:0] _18503 = {_0, _1088} + {_0, _2782};
  wire [1:0] _18504 = {_0, _5918} + {_0, _6270};
  wire [2:0] _18505 = {_0, _18503} + {_0, _18504};
  wire [1:0] _18506 = {_0, _8767} + {_0, _12188};
  wire [3:0] _18507 = {_0, _18505} + {_0, _0, _18506};
  wire _18508 = _12301 < _18507;
  wire _18509 = r1358 ^ _18508;
  wire _18510 = _12298 ? coded_block[1358] : r1358;
  wire _18511 = _12296 ? _18509 : _18510;
  always @ (posedge reset or posedge clock) if (reset) r1358 <= 1'd0; else if (_12300) r1358 <= _18511;
  wire [1:0] _18512 = {_0, _1151} + {_0, _3262};
  wire [1:0] _18513 = {_0, _4350} + {_0, _6942};
  wire [2:0] _18514 = {_0, _18512} + {_0, _18513};
  wire [1:0] _18515 = {_0, _10077} + {_0, _10430};
  wire [3:0] _18516 = {_0, _18514} + {_0, _0, _18515};
  wire _18517 = _12301 < _18516;
  wire _18518 = r1357 ^ _18517;
  wire _18519 = _12298 ? coded_block[1357] : r1357;
  wire _18520 = _12296 ? _18518 : _18519;
  always @ (posedge reset or posedge clock) if (reset) r1357 <= 1'd0; else if (_12300) r1357 <= _18520;
  wire [1:0] _18521 = {_0, _1184} + {_0, _4028};
  wire [1:0] _18522 = {_0, _5342} + {_0, _6431};
  wire [2:0] _18523 = {_0, _18521} + {_0, _18522};
  wire [1:0] _18524 = {_0, _9022} + {_0, _12155};
  wire [3:0] _18525 = {_0, _18523} + {_0, _0, _18524};
  wire _18526 = _12301 < _18525;
  wire _18527 = r1356 ^ _18526;
  wire _18528 = _12298 ? coded_block[1356] : r1356;
  wire _18529 = _12296 ? _18527 : _18528;
  always @ (posedge reset or posedge clock) if (reset) r1356 <= 1'd0; else if (_12300) r1356 <= _18529;
  wire [1:0] _18530 = {_0, _1215} + {_0, _3198};
  wire [1:0] _18531 = {_0, _6108} + {_0, _7420};
  wire [2:0] _18532 = {_0, _18530} + {_0, _18531};
  wire [1:0] _18533 = {_0, _8511} + {_0, _11101};
  wire [3:0] _18534 = {_0, _18532} + {_0, _0, _18533};
  wire _18535 = _12301 < _18534;
  wire _18536 = r1355 ^ _18535;
  wire _18537 = _12298 ? coded_block[1355] : r1355;
  wire _18538 = _12296 ? _18536 : _18537;
  always @ (posedge reset or posedge clock) if (reset) r1355 <= 1'd0; else if (_12300) r1355 <= _18538;
  wire [1:0] _18539 = {_0, _1278} + {_0, _2847};
  wire [1:0] _18540 = {_0, _4798} + {_0, _7357};
  wire [2:0] _18541 = {_0, _18539} + {_0, _18540};
  wire [1:0] _18542 = {_0, _8256} + {_0, _11581};
  wire [3:0] _18543 = {_0, _18541} + {_0, _0, _18542};
  wire _18544 = _12301 < _18543;
  wire _18545 = r1354 ^ _18544;
  wire _18546 = _12298 ? coded_block[1354] : r1354;
  wire _18547 = _12296 ? _18545 : _18546;
  always @ (posedge reset or posedge clock) if (reset) r1354 <= 1'd0; else if (_12300) r1354 <= _18547;
  wire [1:0] _18548 = {_0, _1312} + {_0, _2175};
  wire [1:0] _18549 = {_0, _4926} + {_0, _6877};
  wire [2:0] _18550 = {_0, _18548} + {_0, _18549};
  wire [1:0] _18551 = {_0, _9438} + {_0, _10335};
  wire [3:0] _18552 = {_0, _18550} + {_0, _0, _18551};
  wire _18553 = _12301 < _18552;
  wire _18554 = r1353 ^ _18553;
  wire _18555 = _12298 ? coded_block[1353] : r1353;
  wire _18556 = _12296 ? _18554 : _18555;
  always @ (posedge reset or posedge clock) if (reset) r1353 <= 1'd0; else if (_12300) r1353 <= _18556;
  wire [1:0] _18557 = {_0, _1343} + {_0, _3422};
  wire [1:0] _18558 = {_0, _4256} + {_0, _7005};
  wire [2:0] _18559 = {_0, _18557} + {_0, _18558};
  wire [1:0] _18560 = {_0, _8957} + {_0, _11516};
  wire [3:0] _18561 = {_0, _18559} + {_0, _0, _18560};
  wire _18562 = _12301 < _18561;
  wire _18563 = r1352 ^ _18562;
  wire _18564 = _12298 ? coded_block[1352] : r1352;
  wire _18565 = _12296 ? _18563 : _18564;
  always @ (posedge reset or posedge clock) if (reset) r1352 <= 1'd0; else if (_12300) r1352 <= _18565;
  wire [1:0] _18566 = {_0, _1375} + {_0, _3390};
  wire [1:0] _18567 = {_0, _5501} + {_0, _6334};
  wire [2:0] _18568 = {_0, _18566} + {_0, _18567};
  wire [1:0] _18569 = {_0, _9085} + {_0, _11038};
  wire [3:0] _18570 = {_0, _18568} + {_0, _0, _18569};
  wire _18571 = _12301 < _18570;
  wire _18572 = r1351 ^ _18571;
  wire _18573 = _12298 ? coded_block[1351] : r1351;
  wire _18574 = _12296 ? _18572 : _18573;
  always @ (posedge reset or posedge clock) if (reset) r1351 <= 1'd0; else if (_12300) r1351 <= _18574;
  wire [1:0] _18575 = {_0, _1406} + {_0, _2208};
  wire [1:0] _18576 = {_0, _5470} + {_0, _7581};
  wire [2:0] _18577 = {_0, _18575} + {_0, _18576};
  wire [1:0] _18578 = {_0, _8415} + {_0, _11165};
  wire [3:0] _18579 = {_0, _18577} + {_0, _0, _18578};
  wire _18580 = _12301 < _18579;
  wire _18581 = r1350 ^ _18580;
  wire _18582 = _12298 ? coded_block[1350] : r1350;
  wire _18583 = _12296 ? _18581 : _18582;
  always @ (posedge reset or posedge clock) if (reset) r1350 <= 1'd0; else if (_12300) r1350 <= _18583;
  wire [1:0] _18584 = {_0, _1439} + {_0, _2494};
  wire [1:0] _18585 = {_0, _4287} + {_0, _7548};
  wire [2:0] _18586 = {_0, _18584} + {_0, _18585};
  wire [1:0] _18587 = {_0, _9661} + {_0, _10493};
  wire [3:0] _18588 = {_0, _18586} + {_0, _0, _18587};
  wire _18589 = _12301 < _18588;
  wire _18590 = r1349 ^ _18589;
  wire _18591 = _12298 ? coded_block[1349] : r1349;
  wire _18592 = _12296 ? _18590 : _18591;
  always @ (posedge reset or posedge clock) if (reset) r1349 <= 1'd0; else if (_12300) r1349 <= _18592;
  wire [1:0] _18593 = {_0, _1470} + {_0, _3901};
  wire [1:0] _18594 = {_0, _4574} + {_0, _6366};
  wire [2:0] _18595 = {_0, _18593} + {_0, _18594};
  wire [1:0] _18596 = {_0, _9630} + {_0, _11740};
  wire [3:0] _18597 = {_0, _18595} + {_0, _0, _18596};
  wire _18598 = _12301 < _18597;
  wire _18599 = r1348 ^ _18598;
  wire _18600 = _12298 ? coded_block[1348] : r1348;
  wire _18601 = _12296 ? _18599 : _18600;
  always @ (posedge reset or posedge clock) if (reset) r1348 <= 1'd0; else if (_12300) r1348 <= _18601;
  wire [1:0] _18602 = {_0, _1502} + {_0, _3742};
  wire [1:0] _18603 = {_0, _5981} + {_0, _6652};
  wire [2:0] _18604 = {_0, _18602} + {_0, _18603};
  wire [1:0] _18605 = {_0, _8446} + {_0, _11708};
  wire [3:0] _18606 = {_0, _18604} + {_0, _0, _18605};
  wire _18607 = _12301 < _18606;
  wire _18608 = r1347 ^ _18607;
  wire _18609 = _12298 ? coded_block[1347] : r1347;
  wire _18610 = _12296 ? _18608 : _18609;
  always @ (posedge reset or posedge clock) if (reset) r1347 <= 1'd0; else if (_12300) r1347 <= _18610;
  wire [1:0] _18611 = {_0, _1533} + {_0, _2081};
  wire [1:0] _18612 = {_0, _5821} + {_0, _8059};
  wire [2:0] _18613 = {_0, _18611} + {_0, _18612};
  wire [1:0] _18614 = {_0, _8736} + {_0, _10527};
  wire [3:0] _18615 = {_0, _18613} + {_0, _0, _18614};
  wire _18616 = _12301 < _18615;
  wire _18617 = r1346 ^ _18616;
  wire _18618 = _12298 ? coded_block[1346] : r1346;
  wire _18619 = _12296 ? _18617 : _18618;
  always @ (posedge reset or posedge clock) if (reset) r1346 <= 1'd0; else if (_12300) r1346 <= _18619;
  wire [1:0] _18620 = {_0, _1568} + {_0, _3773};
  wire [1:0] _18621 = {_0, _4129} + {_0, _7900};
  wire [2:0] _18622 = {_0, _18620} + {_0, _18621};
  wire [1:0] _18623 = {_0, _10141} + {_0, _10814};
  wire [3:0] _18624 = {_0, _18622} + {_0, _0, _18623};
  wire _18625 = _12301 < _18624;
  wire _18626 = r1345 ^ _18625;
  wire _18627 = _12298 ? coded_block[1345] : r1345;
  wire _18628 = _12296 ? _18626 : _18627;
  always @ (posedge reset or posedge clock) if (reset) r1345 <= 1'd0; else if (_12300) r1345 <= _18628;
  wire [1:0] _18629 = {_0, _1599} + {_0, _3964};
  wire [1:0] _18630 = {_0, _5853} + {_0, _6176};
  wire [2:0] _18631 = {_0, _18629} + {_0, _18630};
  wire [1:0] _18632 = {_0, _9980} + {_0, _12219};
  wire [3:0] _18633 = {_0, _18631} + {_0, _0, _18632};
  wire _18634 = _12301 < _18633;
  wire _18635 = r1344 ^ _18634;
  wire _18636 = _12298 ? coded_block[1344] : r1344;
  wire _18637 = _12296 ? _18635 : _18636;
  always @ (posedge reset or posedge clock) if (reset) r1344 <= 1'd0; else if (_12300) r1344 <= _18637;
  wire [1:0] _18638 = {_0, _1631} + {_0, _2592};
  wire [1:0] _18639 = {_0, _6045} + {_0, _7931};
  wire [2:0] _18640 = {_0, _18638} + {_0, _18639};
  wire [1:0] _18641 = {_0, _8225} + {_0, _12061};
  wire [3:0] _18642 = {_0, _18640} + {_0, _0, _18641};
  wire _18643 = _12301 < _18642;
  wire _18644 = r1343 ^ _18643;
  wire _18645 = _12298 ? coded_block[1343] : r1343;
  wire _18646 = _12296 ? _18644 : _18645;
  always @ (posedge reset or posedge clock) if (reset) r1343 <= 1'd0; else if (_12300) r1343 <= _18646;
  wire [1:0] _18647 = {_0, _1662} + {_0, _2336};
  wire [1:0] _18648 = {_0, _4671} + {_0, _8123};
  wire [2:0] _18649 = {_0, _18647} + {_0, _18648};
  wire [1:0] _18650 = {_0, _10014} + {_0, _10272};
  wire [3:0] _18651 = {_0, _18649} + {_0, _0, _18650};
  wire _18652 = _12301 < _18651;
  wire _18653 = r1342 ^ _18652;
  wire _18654 = _12298 ? coded_block[1342] : r1342;
  wire _18655 = _12296 ? _18653 : _18654;
  always @ (posedge reset or posedge clock) if (reset) r1342 <= 1'd0; else if (_12300) r1342 <= _18655;
  wire [1:0] _18656 = {_0, _1695} + {_0, _3549};
  wire [1:0] _18657 = {_0, _4415} + {_0, _6750};
  wire [2:0] _18658 = {_0, _18656} + {_0, _18657};
  wire [1:0] _18659 = {_0, _10204} + {_0, _12092};
  wire [3:0] _18660 = {_0, _18658} + {_0, _0, _18659};
  wire _18661 = _12301 < _18660;
  wire _18662 = r1341 ^ _18661;
  wire _18663 = _12298 ? coded_block[1341] : r1341;
  wire _18664 = _12296 ? _18662 : _18663;
  always @ (posedge reset or posedge clock) if (reset) r1341 <= 1'd0; else if (_12300) r1341 <= _18664;
  wire [1:0] _18665 = {_0, _1726} + {_0, _3615};
  wire [1:0] _18666 = {_0, _5628} + {_0, _6494};
  wire [2:0] _18667 = {_0, _18665} + {_0, _18666};
  wire [1:0] _18668 = {_0, _8830} + {_0, _12282};
  wire [3:0] _18669 = {_0, _18667} + {_0, _0, _18668};
  wire _18670 = _12301 < _18669;
  wire _18671 = r1340 ^ _18670;
  wire _18672 = _12298 ? coded_block[1340] : r1340;
  wire _18673 = _12296 ? _18671 : _18672;
  always @ (posedge reset or posedge clock) if (reset) r1340 <= 1'd0; else if (_12300) r1340 <= _18673;
  wire [1:0] _18674 = {_0, _1758} + {_0, _2399};
  wire [1:0] _18675 = {_0, _5694} + {_0, _7710};
  wire [2:0] _18676 = {_0, _18674} + {_0, _18675};
  wire [1:0] _18677 = {_0, _8574} + {_0, _10910};
  wire [3:0] _18678 = {_0, _18676} + {_0, _0, _18677};
  wire _18679 = _12301 < _18678;
  wire _18680 = r1339 ^ _18679;
  wire _18681 = _12298 ? coded_block[1339] : r1339;
  wire _18682 = _12296 ? _18680 : _18681;
  always @ (posedge reset or posedge clock) if (reset) r1339 <= 1'd0; else if (_12300) r1339 <= _18682;
  wire [1:0] _18683 = {_0, _1789} + {_0, _3104};
  wire [1:0] _18684 = {_0, _4478} + {_0, _7773};
  wire [2:0] _18685 = {_0, _18683} + {_0, _18684};
  wire [1:0] _18686 = {_0, _9790} + {_0, _10654};
  wire [3:0] _18687 = {_0, _18685} + {_0, _0, _18686};
  wire _18688 = _12301 < _18687;
  wire _18689 = r1338 ^ _18688;
  wire _18690 = _12298 ? coded_block[1338] : r1338;
  wire _18691 = _12296 ? _18689 : _18690;
  always @ (posedge reset or posedge clock) if (reset) r1338 <= 1'd0; else if (_12300) r1338 <= _18691;
  wire [1:0] _18692 = {_0, _1854} + {_0, _3517};
  wire [1:0] _18693 = {_0, _5085} + {_0, _7262};
  wire [2:0] _18694 = {_0, _18692} + {_0, _18693};
  wire [1:0] _18695 = {_0, _8638} + {_0, _11933};
  wire [3:0] _18696 = {_0, _18694} + {_0, _0, _18695};
  wire _18697 = _12301 < _18696;
  wire _18698 = r1337 ^ _18697;
  wire _18699 = _12298 ? coded_block[1337] : r1337;
  wire _18700 = _12296 ? _18698 : _18699;
  always @ (posedge reset or posedge clock) if (reset) r1337 <= 1'd0; else if (_12300) r1337 <= _18700;
  wire [1:0] _18701 = {_0, _1886} + {_0, _2367};
  wire [1:0] _18702 = {_0, _5597} + {_0, _7163};
  wire [2:0] _18703 = {_0, _18701} + {_0, _18702};
  wire [1:0] _18704 = {_0, _9342} + {_0, _10717};
  wire [3:0] _18705 = {_0, _18703} + {_0, _0, _18704};
  wire _18706 = _12301 < _18705;
  wire _18707 = r1336 ^ _18706;
  wire _18708 = _12298 ? coded_block[1336] : r1336;
  wire _18709 = _12296 ? _18707 : _18708;
  always @ (posedge reset or posedge clock) if (reset) r1336 <= 1'd0; else if (_12300) r1336 <= _18709;
  wire [1:0] _18710 = {_0, _1981} + {_0, _3231};
  wire [1:0] _18711 = {_0, _4767} + {_0, _7804};
  wire [2:0] _18712 = {_0, _18710} + {_0, _18711};
  wire [1:0] _18713 = {_0, _8607} + {_0, _11837};
  wire [3:0] _18714 = {_0, _18712} + {_0, _0, _18713};
  wire _18715 = _12301 < _18714;
  wire _18716 = r1335 ^ _18715;
  wire _18717 = _12298 ? coded_block[1335] : r1335;
  wire _18718 = _12296 ? _18716 : _18717;
  always @ (posedge reset or posedge clock) if (reset) r1335 <= 1'd0; else if (_12300) r1335 <= _18718;
  wire [1:0] _18719 = {_0, _990} + {_0, _4060};
  wire [1:0] _18720 = {_0, _5853} + {_0, _7100};
  wire [2:0] _18721 = {_0, _18719} + {_0, _18720};
  wire [1:0] _18722 = {_0, _9212} + {_0, _12061};
  wire [3:0] _18723 = {_0, _18721} + {_0, _0, _18722};
  wire _18724 = _12301 < _18723;
  wire _18725 = r1334 ^ _18724;
  wire _18726 = _12298 ? coded_block[1334] : r1334;
  wire _18727 = _12296 ? _18725 : _18726;
  always @ (posedge reset or posedge clock) if (reset) r1334 <= 1'd0; else if (_12300) r1334 <= _18727;
  wire [1:0] _18728 = {_0, _1021} + {_0, _3453};
  wire [1:0] _18729 = {_0, _6139} + {_0, _7931};
  wire [2:0] _18730 = {_0, _18728} + {_0, _18729};
  wire [1:0] _18731 = {_0, _9181} + {_0, _11295};
  wire [3:0] _18732 = {_0, _18730} + {_0, _0, _18731};
  wire _18733 = _12301 < _18732;
  wire _18734 = r1333 ^ _18733;
  wire _18735 = _12298 ? coded_block[1333] : r1333;
  wire _18736 = _12296 ? _18734 : _18735;
  always @ (posedge reset or posedge clock) if (reset) r1333 <= 1'd0; else if (_12300) r1333 <= _18736;
  wire [1:0] _18737 = {_0, _1088} + {_0, _2686};
  wire [1:0] _18738 = {_0, _4542} + {_0, _6973};
  wire [2:0] _18739 = {_0, _18737} + {_0, _18738};
  wire [1:0] _18740 = {_0, _10172} + {_0, _11996};
  wire [3:0] _18741 = {_0, _18739} + {_0, _0, _18740};
  wire _18742 = _12301 < _18741;
  wire _18743 = r1332 ^ _18742;
  wire _18744 = _12298 ? coded_block[1332] : r1332;
  wire _18745 = _12296 ? _18743 : _18744;
  always @ (posedge reset or posedge clock) if (reset) r1332 <= 1'd0; else if (_12300) r1332 <= _18745;
  wire [1:0] _18746 = {_0, _1120} + {_0, _2557};
  wire [1:0] _18747 = {_0, _4767} + {_0, _6621};
  wire [2:0] _18748 = {_0, _18746} + {_0, _18747};
  wire [1:0] _18749 = {_0, _9054} + {_0, _12251};
  wire [3:0] _18750 = {_0, _18748} + {_0, _0, _18749};
  wire _18751 = _12301 < _18750;
  wire _18752 = r1331 ^ _18751;
  wire _18753 = _12298 ? coded_block[1331] : r1331;
  wire _18754 = _12296 ? _18752 : _18753;
  always @ (posedge reset or posedge clock) if (reset) r1331 <= 1'd0; else if (_12300) r1331 <= _18754;
  wire [1:0] _18755 = {_0, _1151} + {_0, _2910};
  wire [1:0] _18756 = {_0, _4640} + {_0, _6845};
  wire [2:0] _18757 = {_0, _18755} + {_0, _18756};
  wire [1:0] _18758 = {_0, _8701} + {_0, _11132};
  wire [3:0] _18759 = {_0, _18757} + {_0, _0, _18758};
  wire _18760 = _12301 < _18759;
  wire _18761 = r1330 ^ _18760;
  wire _18762 = _12298 ? coded_block[1330] : r1330;
  wire _18763 = _12296 ? _18761 : _18762;
  always @ (posedge reset or posedge clock) if (reset) r1330 <= 1'd0; else if (_12300) r1330 <= _18763;
  wire [1:0] _18764 = {_0, _1184} + {_0, _3646};
  wire [1:0] _18765 = {_0, _4989} + {_0, _6718};
  wire [2:0] _18766 = {_0, _18764} + {_0, _18765};
  wire [1:0] _18767 = {_0, _8926} + {_0, _10783};
  wire [3:0] _18768 = {_0, _18766} + {_0, _0, _18767};
  wire _18769 = _12301 < _18768;
  wire _18770 = r1329 ^ _18769;
  wire _18771 = _12298 ? coded_block[1329] : r1329;
  wire _18772 = _12296 ? _18770 : _18771;
  always @ (posedge reset or posedge clock) if (reset) r1329 <= 1'd0; else if (_12300) r1329 <= _18772;
  wire [1:0] _18773 = {_0, _672} + {_0, _3933};
  wire [1:0] _18774 = {_0, _5470} + {_0, _6494};
  wire [2:0] _18775 = {_0, _18773} + {_0, _18774};
  wire [1:0] _18776 = {_0, _9311} + {_0, _10527};
  wire [3:0] _18777 = {_0, _18775} + {_0, _0, _18776};
  wire _18778 = _12301 < _18777;
  wire _18779 = r1328 ^ _18778;
  wire _18780 = _12298 ? coded_block[1328] : r1328;
  wire _18781 = _12296 ? _18779 : _18780;
  always @ (posedge reset or posedge clock) if (reset) r1328 <= 1'd0; else if (_12300) r1328 <= _18781;
  wire [1:0] _18782 = {_0, _703} + {_0, _3005};
  wire [1:0] _18783 = {_0, _6012} + {_0, _7548};
  wire [2:0] _18784 = {_0, _18782} + {_0, _18783};
  wire [1:0] _18785 = {_0, _8574} + {_0, _11389};
  wire [3:0] _18786 = {_0, _18784} + {_0, _0, _18785};
  wire _18787 = _12301 < _18786;
  wire _18788 = r1327 ^ _18787;
  wire _18789 = _12298 ? coded_block[1327] : r1327;
  wire _18790 = _12296 ? _18788 : _18789;
  always @ (posedge reset or posedge clock) if (reset) r1327 <= 1'd0; else if (_12300) r1327 <= _18790;
  wire [1:0] _18791 = {_0, _735} + {_0, _3325};
  wire [1:0] _18792 = {_0, _5085} + {_0, _8092};
  wire [2:0] _18793 = {_0, _18791} + {_0, _18792};
  wire [1:0] _18794 = {_0, _9630} + {_0, _10654};
  wire [3:0] _18795 = {_0, _18793} + {_0, _0, _18794};
  wire _18796 = _12301 < _18795;
  wire _18797 = r1326 ^ _18796;
  wire _18798 = _12298 ? coded_block[1326] : r1326;
  wire _18799 = _12296 ? _18797 : _18798;
  always @ (posedge reset or posedge clock) if (reset) r1326 <= 1'd0; else if (_12300) r1326 <= _18799;
  wire [1:0] _18800 = {_0, _766} + {_0, _3773};
  wire [1:0] _18801 = {_0, _5407} + {_0, _7163};
  wire [2:0] _18802 = {_0, _18800} + {_0, _18801};
  wire [1:0] _18803 = {_0, _10172} + {_0, _11708};
  wire [3:0] _18804 = {_0, _18802} + {_0, _0, _18803};
  wire _18805 = _12301 < _18804;
  wire _18806 = r1325 ^ _18805;
  wire _18807 = _12298 ? coded_block[1325] : r1325;
  wire _18808 = _12296 ? _18806 : _18807;
  always @ (posedge reset or posedge clock) if (reset) r1325 <= 1'd0; else if (_12300) r1325 <= _18808;
  wire [1:0] _18809 = {_0, _800} + {_0, _3135};
  wire [1:0] _18810 = {_0, _5853} + {_0, _7485};
  wire [2:0] _18811 = {_0, _18809} + {_0, _18810};
  wire [1:0] _18812 = {_0, _9248} + {_0, _12251};
  wire [3:0] _18813 = {_0, _18811} + {_0, _0, _18812};
  wire _18814 = _12301 < _18813;
  wire _18815 = r1324 ^ _18814;
  wire _18816 = _12298 ? coded_block[1324] : r1324;
  wire _18817 = _12296 ? _18815 : _18816;
  always @ (posedge reset or posedge clock) if (reset) r1324 <= 1'd0; else if (_12300) r1324 <= _18817;
  wire [1:0] _18818 = {_0, _831} + {_0, _4060};
  wire [1:0] _18819 = {_0, _5215} + {_0, _7931};
  wire [2:0] _18820 = {_0, _18818} + {_0, _18819};
  wire [1:0] _18821 = {_0, _9566} + {_0, _11326};
  wire [3:0] _18822 = {_0, _18820} + {_0, _0, _18821};
  wire _18823 = _12301 < _18822;
  wire _18824 = r1323 ^ _18823;
  wire _18825 = _12298 ? coded_block[1323] : r1323;
  wire _18826 = _12296 ? _18824 : _18825;
  always @ (posedge reset or posedge clock) if (reset) r1323 <= 1'd0; else if (_12300) r1323 <= _18826;
  wire [1:0] _18827 = {_0, _863} + {_0, _2144};
  wire [1:0] _18828 = {_0, _6139} + {_0, _7293};
  wire [2:0] _18829 = {_0, _18827} + {_0, _18828};
  wire [1:0] _18830 = {_0, _10014} + {_0, _11644};
  wire [3:0] _18831 = {_0, _18829} + {_0, _0, _18830};
  wire _18832 = _12301 < _18831;
  wire _18833 = r1322 ^ _18832;
  wire _18834 = _12298 ? coded_block[1322] : r1322;
  wire _18835 = _12296 ? _18833 : _18834;
  always @ (posedge reset or posedge clock) if (reset) r1322 <= 1'd0; else if (_12300) r1322 <= _18835;
  wire [1:0] _18836 = {_0, _894} + {_0, _3615};
  wire [1:0] _18837 = {_0, _4223} + {_0, _6207};
  wire [2:0] _18838 = {_0, _18836} + {_0, _18837};
  wire [1:0] _18839 = {_0, _9375} + {_0, _12092};
  wire [3:0] _18840 = {_0, _18838} + {_0, _0, _18839};
  wire _18841 = _12301 < _18840;
  wire _18842 = r1321 ^ _18841;
  wire _18843 = _12298 ? coded_block[1321] : r1321;
  wire _18844 = _12296 ? _18842 : _18843;
  always @ (posedge reset or posedge clock) if (reset) r1321 <= 1'd0; else if (_12300) r1321 <= _18844;
  wire [1:0] _18845 = {_0, _927} + {_0, _3870};
  wire [1:0] _18846 = {_0, _5694} + {_0, _6303};
  wire [2:0] _18847 = {_0, _18845} + {_0, _18846};
  wire [1:0] _18848 = {_0, _8288} + {_0, _11453};
  wire [3:0] _18849 = {_0, _18847} + {_0, _0, _18848};
  wire _18850 = _12301 < _18849;
  wire _18851 = r1320 ^ _18850;
  wire _18852 = _12298 ? coded_block[1320] : r1320;
  wire _18853 = _12296 ? _18851 : _18852;
  always @ (posedge reset or posedge clock) if (reset) r1320 <= 1'd0; else if (_12300) r1320 <= _18853;
  wire [1:0] _18854 = {_0, _958} + {_0, _2750};
  wire [1:0] _18855 = {_0, _5949} + {_0, _7773};
  wire [2:0] _18856 = {_0, _18854} + {_0, _18855};
  wire [1:0] _18857 = {_0, _8383} + {_0, _10366};
  wire [3:0] _18858 = {_0, _18856} + {_0, _0, _18857};
  wire _18859 = _12301 < _18858;
  wire _18860 = r1319 ^ _18859;
  wire _18861 = _12298 ? coded_block[1319] : r1319;
  wire _18862 = _12296 ? _18860 : _18861;
  always @ (posedge reset or posedge clock) if (reset) r1319 <= 1'd0; else if (_12300) r1319 <= _18862;
  wire [1:0] _18863 = {_0, _990} + {_0, _2399};
  wire [1:0] _18864 = {_0, _4830} + {_0, _8028};
  wire [2:0] _18865 = {_0, _18863} + {_0, _18864};
  wire [1:0] _18866 = {_0, _9853} + {_0, _10462};
  wire [3:0] _18867 = {_0, _18865} + {_0, _0, _18866};
  wire _18868 = _12301 < _18867;
  wire _18869 = r1318 ^ _18868;
  wire _18870 = _12298 ? coded_block[1318] : r1318;
  wire _18871 = _12296 ? _18869 : _18870;
  always @ (posedge reset or posedge clock) if (reset) r1318 <= 1'd0; else if (_12300) r1318 <= _18871;
  wire [1:0] _18872 = {_0, _1021} + {_0, _2623};
  wire [1:0] _18873 = {_0, _4478} + {_0, _6908};
  wire [2:0] _18874 = {_0, _18872} + {_0, _18873};
  wire [1:0] _18875 = {_0, _10108} + {_0, _11933};
  wire [3:0] _18876 = {_0, _18874} + {_0, _0, _18875};
  wire _18877 = _12301 < _18876;
  wire _18878 = r1317 ^ _18877;
  wire _18879 = _12298 ? coded_block[1317] : r1317;
  wire _18880 = _12296 ? _18878 : _18879;
  always @ (posedge reset or posedge clock) if (reset) r1317 <= 1'd0; else if (_12300) r1317 <= _18880;
  wire [1:0] _18881 = {_0, _1057} + {_0, _2494};
  wire [1:0] _18882 = {_0, _4703} + {_0, _6558};
  wire [2:0] _18883 = {_0, _18881} + {_0, _18882};
  wire [1:0] _18884 = {_0, _8991} + {_0, _12188};
  wire [3:0] _18885 = {_0, _18883} + {_0, _0, _18884};
  wire _18886 = _12301 < _18885;
  wire _18887 = r1316 ^ _18886;
  wire _18888 = _12298 ? coded_block[1316] : r1316;
  wire _18889 = _12296 ? _18887 : _18888;
  always @ (posedge reset or posedge clock) if (reset) r1316 <= 1'd0; else if (_12300) r1316 <= _18889;
  wire [1:0] _18890 = {_0, _1088} + {_0, _2847};
  wire [1:0] _18891 = {_0, _4574} + {_0, _6781};
  wire [2:0] _18892 = {_0, _18890} + {_0, _18891};
  wire [1:0] _18893 = {_0, _8638} + {_0, _11069};
  wire [3:0] _18894 = {_0, _18892} + {_0, _0, _18893};
  wire _18895 = _12301 < _18894;
  wire _18896 = r1315 ^ _18895;
  wire _18897 = _12298 ? coded_block[1315] : r1315;
  wire _18898 = _12296 ? _18896 : _18897;
  always @ (posedge reset or posedge clock) if (reset) r1315 <= 1'd0; else if (_12300) r1315 <= _18898;
  wire [1:0] _18899 = {_0, _1120} + {_0, _3580};
  wire [1:0] _18900 = {_0, _4926} + {_0, _6652};
  wire [2:0] _18901 = {_0, _18899} + {_0, _18900};
  wire [1:0] _18902 = {_0, _8863} + {_0, _10717};
  wire [3:0] _18903 = {_0, _18901} + {_0, _0, _18902};
  wire _18904 = _12301 < _18903;
  wire _18905 = r1314 ^ _18904;
  wire _18906 = _12298 ? coded_block[1314] : r1314;
  wire _18907 = _12296 ? _18905 : _18906;
  always @ (posedge reset or posedge clock) if (reset) r1314 <= 1'd0; else if (_12300) r1314 <= _18907;
  wire [1:0] _18908 = {_0, _1151} + {_0, _2175};
  wire [1:0] _18909 = {_0, _5663} + {_0, _7005};
  wire [2:0] _18910 = {_0, _18908} + {_0, _18909};
  wire [1:0] _18911 = {_0, _8736} + {_0, _10941};
  wire [3:0] _18912 = {_0, _18910} + {_0, _0, _18911};
  wire _18913 = _12301 < _18912;
  wire _18914 = r1313 ^ _18913;
  wire _18915 = _12298 ? coded_block[1313] : r1313;
  wire _18916 = _12296 ? _18914 : _18915;
  always @ (posedge reset or posedge clock) if (reset) r1313 <= 1'd0; else if (_12300) r1313 <= _18916;
  wire [1:0] _18917 = {_0, _1215} + {_0, _3359};
  wire [1:0] _18918 = {_0, _5821} + {_0, _6334};
  wire [2:0] _18919 = {_0, _18917} + {_0, _18918};
  wire [1:0] _18920 = {_0, _9822} + {_0, _11165};
  wire [3:0] _18921 = {_0, _18919} + {_0, _0, _18920};
  wire _18922 = _12301 < _18921;
  wire _18923 = r1312 ^ _18922;
  wire _18924 = _12298 ? coded_block[1312] : r1312;
  wire _18925 = _12296 ? _18923 : _18924;
  always @ (posedge reset or posedge clock) if (reset) r1312 <= 1'd0; else if (_12300) r1312 <= _18925;
  wire [1:0] _18926 = {_0, _1247} + {_0, _2367};
  wire [1:0] _18927 = {_0, _5438} + {_0, _7900};
  wire [2:0] _18928 = {_0, _18926} + {_0, _18927};
  wire [1:0] _18929 = {_0, _8415} + {_0, _11900};
  wire [3:0] _18930 = {_0, _18928} + {_0, _0, _18929};
  wire _18931 = _12301 < _18930;
  wire _18932 = r1311 ^ _18931;
  wire _18933 = _12298 ? coded_block[1311] : r1311;
  wire _18934 = _12296 ? _18932 : _18933;
  always @ (posedge reset or posedge clock) if (reset) r1311 <= 1'd0; else if (_12300) r1311 <= _18934;
  wire [1:0] _18935 = {_0, _1278} + {_0, _2782};
  wire [1:0] _18936 = {_0, _4447} + {_0, _7517};
  wire [2:0] _18937 = {_0, _18935} + {_0, _18936};
  wire [1:0] _18938 = {_0, _9980} + {_0, _10493};
  wire [3:0] _18939 = {_0, _18937} + {_0, _0, _18938};
  wire _18940 = _12301 < _18939;
  wire _18941 = r1310 ^ _18940;
  wire _18942 = _12298 ? coded_block[1310] : r1310;
  wire _18943 = _12296 ? _18941 : _18942;
  always @ (posedge reset or posedge clock) if (reset) r1310 <= 1'd0; else if (_12300) r1310 <= _18943;
  wire [1:0] _18944 = {_0, _1343} + {_0, _2686};
  wire [1:0] _18945 = {_0, _5342} + {_0, _6942};
  wire [2:0] _18946 = {_0, _18944} + {_0, _18945};
  wire [1:0] _18947 = {_0, _8607} + {_0, _11677};
  wire [3:0] _18948 = {_0, _18946} + {_0, _0, _18947};
  wire _18949 = _12301 < _18948;
  wire _18950 = r1309 ^ _18949;
  wire _18951 = _12298 ? coded_block[1309] : r1309;
  wire _18952 = _12296 ? _18950 : _18951;
  always @ (posedge reset or posedge clock) if (reset) r1309 <= 1'd0; else if (_12300) r1309 <= _18952;
  wire [1:0] _18953 = {_0, _1375} + {_0, _3997};
  wire [1:0] _18954 = {_0, _4767} + {_0, _7420};
  wire [2:0] _18955 = {_0, _18953} + {_0, _18954};
  wire [1:0] _18956 = {_0, _9022} + {_0, _10685};
  wire [3:0] _18957 = {_0, _18955} + {_0, _0, _18956};
  wire _18958 = _12301 < _18957;
  wire _18959 = r1308 ^ _18958;
  wire _18960 = _12298 ? coded_block[1308] : r1308;
  wire _18961 = _12296 ? _18959 : _18960;
  always @ (posedge reset or posedge clock) if (reset) r1308 <= 1'd0; else if (_12300) r1308 <= _18961;
  wire [1:0] _18962 = {_0, _1406} + {_0, _3678};
  wire [1:0] _18963 = {_0, _6076} + {_0, _6845};
  wire [2:0] _18964 = {_0, _18962} + {_0, _18963};
  wire [1:0] _18965 = {_0, _9503} + {_0, _11101};
  wire [3:0] _18966 = {_0, _18964} + {_0, _0, _18965};
  wire _18967 = _12301 < _18966;
  wire _18968 = r1307 ^ _18967;
  wire _18969 = _12298 ? coded_block[1307] : r1307;
  wire _18970 = _12296 ? _18968 : _18969;
  always @ (posedge reset or posedge clock) if (reset) r1307 <= 1'd0; else if (_12300) r1307 <= _18970;
  wire [1:0] _18971 = {_0, _1439} + {_0, _3836};
  wire [1:0] _18972 = {_0, _5757} + {_0, _8155};
  wire [2:0] _18973 = {_0, _18971} + {_0, _18972};
  wire [1:0] _18974 = {_0, _8926} + {_0, _11581};
  wire [3:0] _18975 = {_0, _18973} + {_0, _0, _18974};
  wire _18976 = _12301 < _18975;
  wire _18977 = r1306 ^ _18976;
  wire _18978 = _12298 ? coded_block[1306] : r1306;
  wire _18979 = _12296 ? _18977 : _18978;
  always @ (posedge reset or posedge clock) if (reset) r1306 <= 1'd0; else if (_12300) r1306 <= _18979;
  wire [1:0] _18980 = {_0, _1470} + {_0, _3646};
  wire [1:0] _18981 = {_0, _5918} + {_0, _7837};
  wire [2:0] _18982 = {_0, _18980} + {_0, _18981};
  wire [1:0] _18983 = {_0, _10235} + {_0, _11004};
  wire [3:0] _18984 = {_0, _18982} + {_0, _0, _18983};
  wire _18985 = _12301 < _18984;
  wire _18986 = r1305 ^ _18985;
  wire _18987 = _12298 ? coded_block[1305] : r1305;
  wire _18988 = _12296 ? _18986 : _18987;
  always @ (posedge reset or posedge clock) if (reset) r1305 <= 1'd0; else if (_12300) r1305 <= _18988;
  wire [1:0] _18989 = {_0, _1502} + {_0, _4028};
  wire [1:0] _18990 = {_0, _5726} + {_0, _7996};
  wire [2:0] _18991 = {_0, _18989} + {_0, _18990};
  wire [1:0] _18992 = {_0, _9917} + {_0, _10303};
  wire [3:0] _18993 = {_0, _18991} + {_0, _0, _18992};
  wire _18994 = _12301 < _18993;
  wire _18995 = r1304 ^ _18994;
  wire _18996 = _12298 ? coded_block[1304] : r1304;
  wire _18997 = _12296 ? _18995 : _18996;
  always @ (posedge reset or posedge clock) if (reset) r1304 <= 1'd0; else if (_12300) r1304 <= _18997;
  wire [1:0] _18998 = {_0, _1599} + {_0, _3517};
  wire [1:0] _18999 = {_0, _5022} + {_0, _7326};
  wire [2:0] _19000 = {_0, _18998} + {_0, _18999};
  wire [1:0] _19001 = {_0, _8256} + {_0, _11964};
  wire [3:0] _19002 = {_0, _19000} + {_0, _0, _19001};
  wire _19003 = _12301 < _19002;
  wire _19004 = r1303 ^ _19003;
  wire _19005 = _12298 ? coded_block[1303] : r1303;
  wire _19006 = _12296 ? _19004 : _19005;
  always @ (posedge reset or posedge clock) if (reset) r1303 <= 1'd0; else if (_12300) r1303 <= _19006;
  wire [1:0] _19007 = {_0, _1631} + {_0, _3453};
  wire [1:0] _19008 = {_0, _5597} + {_0, _7100};
  wire [2:0] _19009 = {_0, _19007} + {_0, _19008};
  wire [1:0] _19010 = {_0, _9406} + {_0, _10335};
  wire [3:0] _19011 = {_0, _19009} + {_0, _0, _19010};
  wire _19012 = _12301 < _19011;
  wire _19013 = r1302 ^ _19012;
  wire _19014 = _12298 ? coded_block[1302] : r1302;
  wire _19015 = _12296 ? _19013 : _19014;
  always @ (posedge reset or posedge clock) if (reset) r1302 <= 1'd0; else if (_12300) r1302 <= _19015;
  wire [1:0] _19016 = {_0, _1695} + {_0, _3231};
  wire [1:0] _19017 = {_0, _4640} + {_0, _7612};
  wire [2:0] _19018 = {_0, _19016} + {_0, _19017};
  wire [1:0] _19019 = {_0, _9759} + {_0, _11259};
  wire [3:0] _19020 = {_0, _19018} + {_0, _0, _19019};
  wire _19021 = _12301 < _19020;
  wire _19022 = r1301 ^ _19021;
  wire _19023 = _12298 ? coded_block[1301] : r1301;
  wire _19024 = _12296 ? _19022 : _19023;
  always @ (posedge reset or posedge clock) if (reset) r1301 <= 1'd0; else if (_12300) r1301 <= _19024;
  wire [1:0] _19025 = {_0, _1758} + {_0, _2526};
  wire [1:0] _19026 = {_0, _4895} + {_0, _7389};
  wire [2:0] _19027 = {_0, _19025} + {_0, _19026};
  wire [1:0] _19028 = {_0, _8799} + {_0, _11771};
  wire [3:0] _19029 = {_0, _19027} + {_0, _0, _19028};
  wire _19030 = _12301 < _19029;
  wire _19031 = r1300 ^ _19030;
  wire _19032 = _12298 ? coded_block[1300] : r1300;
  wire _19033 = _12296 ? _19031 : _19032;
  always @ (posedge reset or posedge clock) if (reset) r1300 <= 1'd0; else if (_12300) r1300 <= _19033;
  wire [1:0] _19034 = {_0, _1789} + {_0, _3486};
  wire [1:0] _19035 = {_0, _4605} + {_0, _6973};
  wire [2:0] _19036 = {_0, _19034} + {_0, _19035};
  wire [1:0] _19037 = {_0, _9469} + {_0, _10877};
  wire [3:0] _19038 = {_0, _19036} + {_0, _0, _19037};
  wire _19039 = _12301 < _19038;
  wire _19040 = r1299 ^ _19039;
  wire _19041 = _12298 ? coded_block[1299] : r1299;
  wire _19042 = _12296 ? _19040 : _19041;
  always @ (posedge reset or posedge clock) if (reset) r1299 <= 1'd0; else if (_12300) r1299 <= _19042;
  wire [1:0] _19043 = {_0, _1823} + {_0, _2974};
  wire [1:0] _19044 = {_0, _5565} + {_0, _6687};
  wire [2:0] _19045 = {_0, _19043} + {_0, _19044};
  wire [1:0] _19046 = {_0, _9054} + {_0, _11550};
  wire [3:0] _19047 = {_0, _19045} + {_0, _0, _19046};
  wire _19048 = _12301 < _19047;
  wire _19049 = r1298 ^ _19048;
  wire _19050 = _12298 ? coded_block[1298] : r1298;
  wire _19051 = _12296 ? _19049 : _19050;
  always @ (posedge reset or posedge clock) if (reset) r1298 <= 1'd0; else if (_12300) r1298 <= _19051;
  wire [1:0] _19052 = {_0, _1854} + {_0, _3964};
  wire [1:0] _19053 = {_0, _5053} + {_0, _7644};
  wire [2:0] _19054 = {_0, _19052} + {_0, _19053};
  wire [1:0] _19055 = {_0, _8767} + {_0, _11132};
  wire [3:0] _19056 = {_0, _19054} + {_0, _0, _19055};
  wire _19057 = _12301 < _19056;
  wire _19058 = r1297 ^ _19057;
  wire _19059 = _12298 ? coded_block[1297] : r1297;
  wire _19060 = _12296 ? _19058 : _19059;
  always @ (posedge reset or posedge clock) if (reset) r1297 <= 1'd0; else if (_12300) r1297 <= _19060;
  wire [1:0] _19061 = {_0, _1917} + {_0, _3901};
  wire [1:0] _19062 = {_0, _4798} + {_0, _8123};
  wire [2:0] _19063 = {_0, _19061} + {_0, _19062};
  wire [1:0] _19064 = {_0, _9212} + {_0, _11806};
  wire [3:0] _19065 = {_0, _19063} + {_0, _0, _19064};
  wire _19066 = _12301 < _19065;
  wire _19067 = r1296 ^ _19066;
  wire _19068 = _12298 ? coded_block[1296] : r1296;
  wire _19069 = _12296 ? _19067 : _19068;
  always @ (posedge reset or posedge clock) if (reset) r1296 <= 1'd0; else if (_12300) r1296 <= _19069;
  wire [1:0] _19070 = {_0, _1950} + {_0, _3422};
  wire [1:0] _19071 = {_0, _5981} + {_0, _6877};
  wire [2:0] _19072 = {_0, _19070} + {_0, _19071};
  wire [1:0] _19073 = {_0, _10204} + {_0, _11295};
  wire [3:0] _19074 = {_0, _19072} + {_0, _0, _19073};
  wire _19075 = _12301 < _19074;
  wire _19076 = r1295 ^ _19075;
  wire _19077 = _12298 ? coded_block[1295] : r1295;
  wire _19078 = _12296 ? _19076 : _19077;
  always @ (posedge reset or posedge clock) if (reset) r1295 <= 1'd0; else if (_12300) r1295 <= _19078;
  wire [1:0] _19079 = {_0, _1981} + {_0, _3549};
  wire [1:0] _19080 = {_0, _5501} + {_0, _8059};
  wire [2:0] _19081 = {_0, _19079} + {_0, _19080};
  wire [1:0] _19082 = {_0, _8957} + {_0, _12282};
  wire [3:0] _19083 = {_0, _19081} + {_0, _0, _19082};
  wire _19084 = _12301 < _19083;
  wire _19085 = r1294 ^ _19084;
  wire _19086 = _12298 ? coded_block[1294] : r1294;
  wire _19087 = _12296 ? _19085 : _19086;
  always @ (posedge reset or posedge clock) if (reset) r1294 <= 1'd0; else if (_12300) r1294 <= _19087;
  wire [1:0] _19088 = {_0, _2013} + {_0, _2878};
  wire [1:0] _19089 = {_0, _5628} + {_0, _7581};
  wire [2:0] _19090 = {_0, _19088} + {_0, _19089};
  wire [1:0] _19091 = {_0, _10141} + {_0, _11038};
  wire [3:0] _19092 = {_0, _19090} + {_0, _0, _19091};
  wire _19093 = _12301 < _19092;
  wire _19094 = r1293 ^ _19093;
  wire _19095 = _12298 ? coded_block[1293] : r1293;
  wire _19096 = _12296 ? _19094 : _19095;
  always @ (posedge reset or posedge clock) if (reset) r1293 <= 1'd0; else if (_12300) r1293 <= _19096;
  wire [1:0] _19097 = {_0, _65} + {_0, _4091};
  wire [1:0] _19098 = {_0, _4192} + {_0, _7036};
  wire [2:0] _19099 = {_0, _19097} + {_0, _19098};
  wire [1:0] _19100 = {_0, _9790} + {_0, _11740};
  wire [3:0] _19101 = {_0, _19099} + {_0, _0, _19100};
  wire _19102 = _12301 < _19101;
  wire _19103 = r1292 ^ _19102;
  wire _19104 = _12298 ? coded_block[1292] : r1292;
  wire _19105 = _12296 ? _19103 : _19104;
  always @ (posedge reset or posedge clock) if (reset) r1292 <= 1'd0; else if (_12300) r1292 <= _19105;
  wire [1:0] _19106 = {_0, _97} + {_0, _2910};
  wire [1:0] _19107 = {_0, _4160} + {_0, _6270};
  wire [2:0] _19108 = {_0, _19106} + {_0, _19107};
  wire [1:0] _19109 = {_0, _9118} + {_0, _11869};
  wire [3:0] _19110 = {_0, _19108} + {_0, _0, _19109};
  wire _19111 = _12301 < _19110;
  wire _19112 = r1291 ^ _19111;
  wire _19113 = _12298 ? coded_block[1291] : r1291;
  wire _19114 = _12296 ? _19112 : _19113;
  always @ (posedge reset or posedge clock) if (reset) r1291 <= 1'd0; else if (_12300) r1291 <= _19114;
  wire [1:0] _19115 = {_0, _128} + {_0, _3198};
  wire [1:0] _19116 = {_0, _4989} + {_0, _6239};
  wire [2:0] _19117 = {_0, _19115} + {_0, _19116};
  wire [1:0] _19118 = {_0, _8352} + {_0, _11196};
  wire [3:0] _19119 = {_0, _19117} + {_0, _0, _19118};
  wire _19120 = _12301 < _19119;
  wire _19121 = r1290 ^ _19120;
  wire _19122 = _12298 ? coded_block[1290] : r1290;
  wire _19123 = _12296 ? _19121 : _19122;
  always @ (posedge reset or posedge clock) if (reset) r1290 <= 1'd0; else if (_12300) r1290 <= _19123;
  wire [1:0] _19124 = {_0, _161} + {_0, _2592};
  wire [1:0] _19125 = {_0, _5279} + {_0, _7069};
  wire [2:0] _19126 = {_0, _19124} + {_0, _19125};
  wire [1:0] _19127 = {_0, _8319} + {_0, _10430};
  wire [3:0] _19128 = {_0, _19126} + {_0, _0, _19127};
  wire _19129 = _12301 < _19128;
  wire _19130 = r1289 ^ _19129;
  wire _19131 = _12298 ? coded_block[1289] : r1289;
  wire _19132 = _12296 ? _19130 : _19131;
  always @ (posedge reset or posedge clock) if (reset) r1289 <= 1'd0; else if (_12300) r1289 <= _19132;
  wire [1:0] _19133 = {_0, _192} + {_0, _2430};
  wire [1:0] _19134 = {_0, _4671} + {_0, _7357};
  wire [2:0] _19135 = {_0, _19133} + {_0, _19134};
  wire [1:0] _19136 = {_0, _9149} + {_0, _10399};
  wire [3:0] _19137 = {_0, _19135} + {_0, _0, _19136};
  wire _19138 = _12301 < _19137;
  wire _19139 = r1288 ^ _19138;
  wire _19140 = _12298 ? coded_block[1288] : r1288;
  wire _19141 = _12296 ? _19139 : _19140;
  always @ (posedge reset or posedge clock) if (reset) r1288 <= 1'd0; else if (_12300) r1288 <= _19141;
  wire [1:0] _19142 = {_0, _224} + {_0, _2081};
  wire [1:0] _19143 = {_0, _4511} + {_0, _6750};
  wire [2:0] _19144 = {_0, _19142} + {_0, _19143};
  wire [1:0] _19145 = {_0, _9438} + {_0, _11228};
  wire [3:0] _19146 = {_0, _19144} + {_0, _0, _19145};
  wire _19147 = _12301 < _19146;
  wire _19148 = r1287 ^ _19147;
  wire _19149 = _12298 ? coded_block[1287] : r1287;
  wire _19150 = _12296 ? _19148 : _19149;
  always @ (posedge reset or posedge clock) if (reset) r1287 <= 1'd0; else if (_12300) r1287 <= _19150;
  wire [1:0] _19151 = {_0, _255} + {_0, _2463};
  wire [1:0] _19152 = {_0, _4129} + {_0, _6589};
  wire [2:0] _19153 = {_0, _19151} + {_0, _19152};
  wire [1:0] _19154 = {_0, _8830} + {_0, _11516};
  wire [3:0] _19155 = {_0, _19153} + {_0, _0, _19154};
  wire _19156 = _12301 < _19155;
  wire _19157 = r1286 ^ _19156;
  wire _19158 = _12298 ? coded_block[1286] : r1286;
  wire _19159 = _12296 ? _19157 : _19158;
  always @ (posedge reset or posedge clock) if (reset) r1286 <= 1'd0; else if (_12300) r1286 <= _19159;
  wire [1:0] _19160 = {_0, _320} + {_0, _3294};
  wire [1:0] _19161 = {_0, _4734} + {_0, _6621};
  wire [2:0] _19162 = {_0, _19160} + {_0, _19161};
  wire [1:0] _19163 = {_0, _8225} + {_0, _10748};
  wire [3:0] _19164 = {_0, _19162} + {_0, _0, _19163};
  wire _19165 = _12301 < _19164;
  wire _19166 = r1285 ^ _19165;
  wire _19167 = _12298 ? coded_block[1285] : r1285;
  wire _19168 = _12296 ? _19166 : _19167;
  always @ (posedge reset or posedge clock) if (reset) r1285 <= 1'd0; else if (_12300) r1285 <= _19168;
  wire [1:0] _19169 = {_0, _416} + {_0, _2302};
  wire [1:0] _19170 = {_0, _4319} + {_0, _7199};
  wire [2:0] _19171 = {_0, _19169} + {_0, _19170};
  wire [1:0] _19172 = {_0, _9534} + {_0, _10973};
  wire [3:0] _19173 = {_0, _19171} + {_0, _0, _19172};
  wire _19174 = _12301 < _19173;
  wire _19175 = r1284 ^ _19174;
  wire _19176 = _12298 ? coded_block[1284] : r1284;
  wire _19177 = _12296 ? _19175 : _19176;
  always @ (posedge reset or posedge clock) if (reset) r1284 <= 1'd0; else if (_12300) r1284 <= _19177;
  wire [1:0] _19178 = {_0, _447} + {_0, _3104};
  wire [1:0] _19179 = {_0, _4384} + {_0, _6397};
  wire [2:0] _19180 = {_0, _19178} + {_0, _19179};
  wire [1:0] _19181 = {_0, _9279} + {_0, _11613};
  wire [3:0] _19182 = {_0, _19180} + {_0, _0, _19181};
  wire _19183 = _12301 < _19182;
  wire _19184 = r1283 ^ _19183;
  wire _19185 = _12298 ? coded_block[1283] : r1283;
  wire _19186 = _12296 ? _19184 : _19185;
  always @ (posedge reset or posedge clock) if (reset) r1283 <= 1'd0; else if (_12300) r1283 <= _19186;
  wire [1:0] _19187 = {_0, _1215} + {_0, _2239};
  wire [1:0] _19188 = {_0, _5726} + {_0, _7069};
  wire [2:0] _19189 = {_0, _19187} + {_0, _19188};
  wire [1:0] _19190 = {_0, _8799} + {_0, _11004};
  wire [3:0] _19191 = {_0, _19189} + {_0, _0, _19190};
  wire _19192 = _12301 < _19191;
  wire _19193 = r1282 ^ _19192;
  wire _19194 = _12298 ? coded_block[1282] : r1282;
  wire _19195 = _12296 ? _19193 : _19194;
  always @ (posedge reset or posedge clock) if (reset) r1282 <= 1'd0; else if (_12300) r1282 <= _19195;
  wire [1:0] _19196 = {_0, _1247} + {_0, _3805};
  wire [1:0] _19197 = {_0, _4319} + {_0, _7804};
  wire [2:0] _19198 = {_0, _19196} + {_0, _19197};
  wire [1:0] _19199 = {_0, _9149} + {_0, _10877};
  wire [3:0] _19200 = {_0, _19198} + {_0, _0, _19199};
  wire _19201 = _12301 < _19200;
  wire _19202 = r1281 ^ _19201;
  wire _19203 = _12298 ? coded_block[1281] : r1281;
  wire _19204 = _12296 ? _19202 : _19203;
  always @ (posedge reset or posedge clock) if (reset) r1281 <= 1'd0; else if (_12300) r1281 <= _19204;
  wire [1:0] _19205 = {_0, _1278} + {_0, _3422};
  wire [1:0] _19206 = {_0, _5884} + {_0, _6397};
  wire [2:0] _19207 = {_0, _19205} + {_0, _19206};
  wire [1:0] _19208 = {_0, _9886} + {_0, _11228};
  wire [3:0] _19209 = {_0, _19207} + {_0, _0, _19208};
  wire _19210 = _12301 < _19209;
  wire _19211 = r1280 ^ _19210;
  wire _19212 = _12298 ? coded_block[1280] : r1280;
  wire _19213 = _12296 ? _19211 : _19212;
  always @ (posedge reset or posedge clock) if (reset) r1280 <= 1'd0; else if (_12300) r1280 <= _19213;
  wire [1:0] _19214 = {_0, _1312} + {_0, _2430};
  wire [1:0] _19215 = {_0, _5501} + {_0, _7965};
  wire [2:0] _19216 = {_0, _19214} + {_0, _19215};
  wire [1:0] _19217 = {_0, _8480} + {_0, _11964};
  wire [3:0] _19218 = {_0, _19216} + {_0, _0, _19217};
  wire _19219 = _12301 < _19218;
  wire _19220 = r1279 ^ _19219;
  wire _19221 = _12298 ? coded_block[1279] : r1279;
  wire _19222 = _12296 ? _19220 : _19221;
  always @ (posedge reset or posedge clock) if (reset) r1279 <= 1'd0; else if (_12300) r1279 <= _19222;
  wire [1:0] _19223 = {_0, _1343} + {_0, _2847};
  wire [1:0] _19224 = {_0, _4511} + {_0, _7581};
  wire [2:0] _19225 = {_0, _19223} + {_0, _19224};
  wire [1:0] _19226 = {_0, _10045} + {_0, _10558};
  wire [3:0] _19227 = {_0, _19225} + {_0, _0, _19226};
  wire _19228 = _12301 < _19227;
  wire _19229 = r1278 ^ _19228;
  wire _19230 = _12298 ? coded_block[1278] : r1278;
  wire _19231 = _12296 ? _19229 : _19230;
  always @ (posedge reset or posedge clock) if (reset) r1278 <= 1'd0; else if (_12300) r1278 <= _19231;
  wire [1:0] _19232 = {_0, _1406} + {_0, _2750};
  wire [1:0] _19233 = {_0, _5407} + {_0, _7005};
  wire [2:0] _19234 = {_0, _19232} + {_0, _19233};
  wire [1:0] _19235 = {_0, _8670} + {_0, _11740};
  wire [3:0] _19236 = {_0, _19234} + {_0, _0, _19235};
  wire _19237 = _12301 < _19236;
  wire _19238 = r1277 ^ _19237;
  wire _19239 = _12298 ? coded_block[1277] : r1277;
  wire _19240 = _12296 ? _19238 : _19239;
  always @ (posedge reset or posedge clock) if (reset) r1277 <= 1'd0; else if (_12300) r1277 <= _19240;
  wire [1:0] _19241 = {_0, _1439} + {_0, _4060};
  wire [1:0] _19242 = {_0, _4830} + {_0, _7485};
  wire [2:0] _19243 = {_0, _19241} + {_0, _19242};
  wire [1:0] _19244 = {_0, _9085} + {_0, _10748};
  wire [3:0] _19245 = {_0, _19243} + {_0, _0, _19244};
  wire _19246 = _12301 < _19245;
  wire _19247 = r1276 ^ _19246;
  wire _19248 = _12298 ? coded_block[1276] : r1276;
  wire _19249 = _12296 ? _19247 : _19248;
  always @ (posedge reset or posedge clock) if (reset) r1276 <= 1'd0; else if (_12300) r1276 <= _19249;
  wire [1:0] _19250 = {_0, _192} + {_0, _2336};
  wire [1:0] _19251 = {_0, _4798} + {_0, _7326};
  wire [2:0] _19252 = {_0, _19250} + {_0, _19251};
  wire [1:0] _19253 = {_0, _8799} + {_0, _12155};
  wire [3:0] _19254 = {_0, _19252} + {_0, _0, _19253};
  wire _19255 = _12301 < _19254;
  wire _19256 = r1275 ^ _19255;
  wire _19257 = _12298 ? coded_block[1275] : r1275;
  wire _19258 = _12296 ? _19256 : _19257;
  always @ (posedge reset or posedge clock) if (reset) r1275 <= 1'd0; else if (_12300) r1275 <= _19258;
  wire [1:0] _19259 = {_0, _224} + {_0, _3359};
  wire [1:0] _19260 = {_0, _4415} + {_0, _6877};
  wire [2:0] _19261 = {_0, _19259} + {_0, _19260};
  wire [1:0] _19262 = {_0, _9406} + {_0, _10877};
  wire [3:0] _19263 = {_0, _19261} + {_0, _0, _19262};
  wire _19264 = _12301 < _19263;
  wire _19265 = r1274 ^ _19264;
  wire _19266 = _12298 ? coded_block[1274] : r1274;
  wire _19267 = _12296 ? _19265 : _19266;
  always @ (posedge reset or posedge clock) if (reset) r1274 <= 1'd0; else if (_12300) r1274 <= _19267;
  wire [1:0] _19268 = {_0, _255} + {_0, _3773};
  wire [1:0] _19269 = {_0, _5438} + {_0, _6494};
  wire [2:0] _19270 = {_0, _19268} + {_0, _19269};
  wire [1:0] _19271 = {_0, _8957} + {_0, _11485};
  wire [3:0] _19272 = {_0, _19270} + {_0, _0, _19271};
  wire _19273 = _12301 < _19272;
  wire _19274 = r1273 ^ _19273;
  wire _19275 = _12298 ? coded_block[1273] : r1273;
  wire _19276 = _12296 ? _19274 : _19275;
  always @ (posedge reset or posedge clock) if (reset) r1273 <= 1'd0; else if (_12300) r1273 <= _19276;
  wire [1:0] _19277 = {_0, _289} + {_0, _2239};
  wire [1:0] _19278 = {_0, _5853} + {_0, _7517};
  wire [2:0] _19279 = {_0, _19277} + {_0, _19278};
  wire [1:0] _19280 = {_0, _8574} + {_0, _11038};
  wire [3:0] _19281 = {_0, _19279} + {_0, _0, _19280};
  wire _19282 = _12301 < _19281;
  wire _19283 = r1272 ^ _19282;
  wire _19284 = _12298 ? coded_block[1272] : r1272;
  wire _19285 = _12296 ? _19283 : _19284;
  always @ (posedge reset or posedge clock) if (reset) r1272 <= 1'd0; else if (_12300) r1272 <= _19285;
  wire [1:0] _19286 = {_0, _320} + {_0, _3678};
  wire [1:0] _19287 = {_0, _4319} + {_0, _7931};
  wire [2:0] _19288 = {_0, _19286} + {_0, _19287};
  wire [1:0] _19289 = {_0, _9597} + {_0, _10654};
  wire [3:0] _19290 = {_0, _19288} + {_0, _0, _19289};
  wire _19291 = _12301 < _19290;
  wire _19292 = r1271 ^ _19291;
  wire _19293 = _12298 ? coded_block[1271] : r1271;
  wire _19294 = _12296 ? _19292 : _19293;
  always @ (posedge reset or posedge clock) if (reset) r1271 <= 1'd0; else if (_12300) r1271 <= _19294;
  wire [1:0] _19295 = {_0, _352} + {_0, _2974};
  wire [1:0] _19296 = {_0, _5757} + {_0, _6397};
  wire [2:0] _19297 = {_0, _19295} + {_0, _19296};
  wire [1:0] _19298 = {_0, _10014} + {_0, _11677};
  wire [3:0] _19299 = {_0, _19297} + {_0, _0, _19298};
  wire _19300 = _12301 < _19299;
  wire _19301 = r1270 ^ _19300;
  wire _19302 = _12298 ? coded_block[1270] : r1270;
  wire _19303 = _12296 ? _19301 : _19302;
  always @ (posedge reset or posedge clock) if (reset) r1270 <= 1'd0; else if (_12300) r1270 <= _19303;
  wire [1:0] _19304 = {_0, _383} + {_0, _2655};
  wire [1:0] _19305 = {_0, _5053} + {_0, _7837};
  wire [2:0] _19306 = {_0, _19304} + {_0, _19305};
  wire [1:0] _19307 = {_0, _8480} + {_0, _12092};
  wire [3:0] _19308 = {_0, _19306} + {_0, _0, _19307};
  wire _19309 = _12301 < _19308;
  wire _19310 = r1269 ^ _19309;
  wire _19311 = _12298 ? coded_block[1269] : r1269;
  wire _19312 = _12296 ? _19310 : _19311;
  always @ (posedge reset or posedge clock) if (reset) r1269 <= 1'd0; else if (_12300) r1269 <= _19312;
  wire [1:0] _19313 = {_0, _416} + {_0, _2813};
  wire [1:0] _19314 = {_0, _4734} + {_0, _7132};
  wire [2:0] _19315 = {_0, _19313} + {_0, _19314};
  wire [1:0] _19316 = {_0, _9917} + {_0, _10558};
  wire [3:0] _19317 = {_0, _19315} + {_0, _0, _19316};
  wire _19318 = _12301 < _19317;
  wire _19319 = r1268 ^ _19318;
  wire _19320 = _12298 ? coded_block[1268] : r1268;
  wire _19321 = _12296 ? _19319 : _19320;
  always @ (posedge reset or posedge clock) if (reset) r1268 <= 1'd0; else if (_12300) r1268 <= _19321;
  wire [1:0] _19322 = {_0, _447} + {_0, _2623};
  wire [1:0] _19323 = {_0, _4895} + {_0, _6814};
  wire [2:0] _19324 = {_0, _19322} + {_0, _19323};
  wire [1:0] _19325 = {_0, _9212} + {_0, _11996};
  wire [3:0] _19326 = {_0, _19324} + {_0, _0, _19325};
  wire _19327 = _12301 < _19326;
  wire _19328 = r1267 ^ _19327;
  wire _19329 = _12298 ? coded_block[1267] : r1267;
  wire _19330 = _12296 ? _19328 : _19329;
  always @ (posedge reset or posedge clock) if (reset) r1267 <= 1'd0; else if (_12300) r1267 <= _19330;
  wire [1:0] _19331 = {_0, _479} + {_0, _3005};
  wire [1:0] _19332 = {_0, _4703} + {_0, _6973};
  wire [2:0] _19333 = {_0, _19331} + {_0, _19332};
  wire [1:0] _19334 = {_0, _8894} + {_0, _11295};
  wire [3:0] _19335 = {_0, _19333} + {_0, _0, _19334};
  wire _19336 = _12301 < _19335;
  wire _19337 = r1266 ^ _19336;
  wire _19338 = _12298 ? coded_block[1266] : r1266;
  wire _19339 = _12296 ? _19337 : _19338;
  always @ (posedge reset or posedge clock) if (reset) r1266 <= 1'd0; else if (_12300) r1266 <= _19339;
  wire [1:0] _19340 = {_0, _510} + {_0, _2144};
  wire [1:0] _19341 = {_0, _5085} + {_0, _6781};
  wire [2:0] _19342 = {_0, _19340} + {_0, _19341};
  wire [1:0] _19343 = {_0, _9054} + {_0, _10973};
  wire [3:0] _19344 = {_0, _19342} + {_0, _0, _19343};
  wire _19345 = _12301 < _19344;
  wire _19346 = r1265 ^ _19345;
  wire _19347 = _12298 ? coded_block[1265] : r1265;
  wire _19348 = _12296 ? _19346 : _19347;
  always @ (posedge reset or posedge clock) if (reset) r1265 <= 1'd0; else if (_12300) r1265 <= _19348;
  wire [1:0] _19349 = {_0, _545} + {_0, _3933};
  wire [1:0] _19350 = {_0, _4223} + {_0, _7163};
  wire [2:0] _19351 = {_0, _19349} + {_0, _19350};
  wire [1:0] _19352 = {_0, _8863} + {_0, _11132};
  wire [3:0] _19353 = {_0, _19351} + {_0, _0, _19352};
  wire _19354 = _12301 < _19353;
  wire _19355 = r1264 ^ _19354;
  wire _19356 = _12298 ? coded_block[1264] : r1264;
  wire _19357 = _12296 ? _19355 : _19356;
  always @ (posedge reset or posedge clock) if (reset) r1264 <= 1'd0; else if (_12300) r1264 <= _19357;
  wire [1:0] _19358 = {_0, _576} + {_0, _2494};
  wire [1:0] _19359 = {_0, _6012} + {_0, _6303};
  wire [2:0] _19360 = {_0, _19358} + {_0, _19359};
  wire [1:0] _19361 = {_0, _9248} + {_0, _10941};
  wire [3:0] _19362 = {_0, _19360} + {_0, _0, _19361};
  wire _19363 = _12301 < _19362;
  wire _19364 = r1263 ^ _19363;
  wire _19365 = _12298 ? coded_block[1263] : r1263;
  wire _19366 = _12296 ? _19364 : _19365;
  always @ (posedge reset or posedge clock) if (reset) r1263 <= 1'd0; else if (_12300) r1263 <= _19366;
  wire [1:0] _19367 = {_0, _608} + {_0, _2430};
  wire [1:0] _19368 = {_0, _4574} + {_0, _8092};
  wire [2:0] _19369 = {_0, _19367} + {_0, _19368};
  wire [1:0] _19370 = {_0, _8383} + {_0, _11326};
  wire [3:0] _19371 = {_0, _19369} + {_0, _0, _19370};
  wire _19372 = _12301 < _19371;
  wire _19373 = r1262 ^ _19372;
  wire _19374 = _12298 ? coded_block[1262] : r1262;
  wire _19375 = _12296 ? _19373 : _19374;
  always @ (posedge reset or posedge clock) if (reset) r1262 <= 1'd0; else if (_12300) r1262 <= _19375;
  wire [1:0] _19376 = {_0, _639} + {_0, _3549};
  wire [1:0] _19377 = {_0, _4511} + {_0, _6652};
  wire [2:0] _19378 = {_0, _19376} + {_0, _19377};
  wire [1:0] _19379 = {_0, _10172} + {_0, _10462};
  wire [3:0] _19380 = {_0, _19378} + {_0, _0, _19379};
  wire _19381 = _12301 < _19380;
  wire _19382 = r1261 ^ _19381;
  wire _19383 = _12298 ? coded_block[1261] : r1261;
  wire _19384 = _12296 ? _19382 : _19383;
  always @ (posedge reset or posedge clock) if (reset) r1261 <= 1'd0; else if (_12300) r1261 <= _19384;
  wire [1:0] _19385 = {_0, _672} + {_0, _2208};
  wire [1:0] _19386 = {_0, _5628} + {_0, _6589};
  wire [2:0] _19387 = {_0, _19385} + {_0, _19386};
  wire [1:0] _19388 = {_0, _8736} + {_0, _12251};
  wire [3:0] _19389 = {_0, _19387} + {_0, _0, _19388};
  wire _19390 = _12301 < _19389;
  wire _19391 = r1260 ^ _19390;
  wire _19392 = _12298 ? coded_block[1260] : r1260;
  wire _19393 = _12296 ? _19391 : _19392;
  always @ (posedge reset or posedge clock) if (reset) r1260 <= 1'd0; else if (_12300) r1260 <= _19393;
  wire [1:0] _19394 = {_0, _703} + {_0, _3805};
  wire [1:0] _19395 = {_0, _4287} + {_0, _7710};
  wire [2:0] _19396 = {_0, _19394} + {_0, _19395};
  wire [1:0] _19397 = {_0, _8670} + {_0, _10814};
  wire [3:0] _19398 = {_0, _19396} + {_0, _0, _19397};
  wire _19399 = _12301 < _19398;
  wire _19400 = r1259 ^ _19399;
  wire _19401 = _12298 ? coded_block[1259] : r1259;
  wire _19402 = _12296 ? _19400 : _19401;
  always @ (posedge reset or posedge clock) if (reset) r1259 <= 1'd0; else if (_12300) r1259 <= _19402;
  wire [1:0] _19403 = {_0, _735} + {_0, _3517};
  wire [1:0] _19404 = {_0, _5884} + {_0, _6366};
  wire [2:0] _19405 = {_0, _19403} + {_0, _19404};
  wire [1:0] _19406 = {_0, _9790} + {_0, _10748};
  wire [3:0] _19407 = {_0, _19405} + {_0, _0, _19406};
  wire _19408 = _12301 < _19407;
  wire _19409 = r1258 ^ _19408;
  wire _19410 = _12298 ? coded_block[1258] : r1258;
  wire _19411 = _12296 ? _19409 : _19410;
  always @ (posedge reset or posedge clock) if (reset) r1258 <= 1'd0; else if (_12300) r1258 <= _19411;
  wire [1:0] _19412 = {_0, _766} + {_0, _2463};
  wire [1:0] _19413 = {_0, _5597} + {_0, _7965};
  wire [2:0] _19414 = {_0, _19412} + {_0, _19413};
  wire [1:0] _19415 = {_0, _8446} + {_0, _11869};
  wire [3:0] _19416 = {_0, _19414} + {_0, _0, _19415};
  wire _19417 = _12301 < _19416;
  wire _19418 = r1257 ^ _19417;
  wire _19419 = _12298 ? coded_block[1257] : r1257;
  wire _19420 = _12296 ? _19418 : _19419;
  always @ (posedge reset or posedge clock) if (reset) r1257 <= 1'd0; else if (_12300) r1257 <= _19420;
  wire [1:0] _19421 = {_0, _831} + {_0, _2941};
  wire [1:0] _19422 = {_0, _6045} + {_0, _6621};
  wire [2:0] _19423 = {_0, _19421} + {_0, _19422};
  wire [1:0] _19424 = {_0, _9759} + {_0, _12124};
  wire [3:0] _19425 = {_0, _19423} + {_0, _0, _19424};
  wire _19426 = _12301 < _19425;
  wire _19427 = r1256 ^ _19426;
  wire _19428 = _12298 ? coded_block[1256] : r1256;
  wire _19429 = _12296 ? _19427 : _19428;
  always @ (posedge reset or posedge clock) if (reset) r1256 <= 1'd0; else if (_12300) r1256 <= _19429;
  wire [1:0] _19430 = {_0, _863} + {_0, _3709};
  wire [1:0] _19431 = {_0, _5022} + {_0, _8123};
  wire [2:0] _19432 = {_0, _19430} + {_0, _19431};
  wire [1:0] _19433 = {_0, _8701} + {_0, _11837};
  wire [3:0] _19434 = {_0, _19432} + {_0, _0, _19433};
  wire _19435 = _12301 < _19434;
  wire _19436 = r1255 ^ _19435;
  wire _19437 = _12298 ? coded_block[1255] : r1255;
  wire _19438 = _12296 ? _19436 : _19437;
  always @ (posedge reset or posedge clock) if (reset) r1255 <= 1'd0; else if (_12300) r1255 <= _19438;
  wire [1:0] _19439 = {_0, _927} + {_0, _2399};
  wire [1:0] _19440 = {_0, _4958} + {_0, _7868};
  wire [2:0] _19441 = {_0, _19439} + {_0, _19440};
  wire [1:0] _19442 = {_0, _9181} + {_0, _12282};
  wire [3:0] _19443 = {_0, _19441} + {_0, _0, _19442};
  wire _19444 = _12301 < _19443;
  wire _19445 = r1254 ^ _19444;
  wire _19446 = _12298 ? coded_block[1254] : r1254;
  wire _19447 = _12296 ? _19445 : _19446;
  always @ (posedge reset or posedge clock) if (reset) r1254 <= 1'd0; else if (_12300) r1254 <= _19447;
  wire [1:0] _19448 = {_0, _958} + {_0, _2526};
  wire [1:0] _19449 = {_0, _4478} + {_0, _7036};
  wire [2:0] _19450 = {_0, _19448} + {_0, _19449};
  wire [1:0] _19451 = {_0, _9949} + {_0, _11259};
  wire [3:0] _19452 = {_0, _19450} + {_0, _0, _19451};
  wire _19453 = _12301 < _19452;
  wire _19454 = r1253 ^ _19453;
  wire _19455 = _12298 ? coded_block[1253] : r1253;
  wire _19456 = _12296 ? _19454 : _19455;
  always @ (posedge reset or posedge clock) if (reset) r1253 <= 1'd0; else if (_12300) r1253 <= _19456;
  wire [1:0] _19457 = {_0, _990} + {_0, _3870};
  wire [1:0] _19458 = {_0, _4605} + {_0, _6558};
  wire [2:0] _19459 = {_0, _19457} + {_0, _19458};
  wire [1:0] _19460 = {_0, _9118} + {_0, _12027};
  wire [3:0] _19461 = {_0, _19459} + {_0, _0, _19460};
  wire _19462 = _12301 < _19461;
  wire _19463 = r1252 ^ _19462;
  wire _19464 = _12298 ? coded_block[1252] : r1252;
  wire _19465 = _12296 ? _19463 : _19464;
  always @ (posedge reset or posedge clock) if (reset) r1252 <= 1'd0; else if (_12300) r1252 <= _19465;
  wire [1:0] _19466 = {_0, _1021} + {_0, _3104};
  wire [1:0] _19467 = {_0, _5949} + {_0, _6687};
  wire [2:0] _19468 = {_0, _19466} + {_0, _19467};
  wire [1:0] _19469 = {_0, _8638} + {_0, _11196};
  wire [3:0] _19470 = {_0, _19468} + {_0, _0, _19469};
  wire _19471 = _12301 < _19470;
  wire _19472 = r1251 ^ _19471;
  wire _19473 = _12298 ? coded_block[1251] : r1251;
  wire _19474 = _12296 ? _19472 : _19473;
  always @ (posedge reset or posedge clock) if (reset) r1251 <= 1'd0; else if (_12300) r1251 <= _19474;
  wire [1:0] _19475 = {_0, _1057} + {_0, _3068};
  wire [1:0] _19476 = {_0, _5183} + {_0, _8028};
  wire [2:0] _19477 = {_0, _19475} + {_0, _19476};
  wire [1:0] _19478 = {_0, _8767} + {_0, _10717};
  wire [3:0] _19479 = {_0, _19477} + {_0, _0, _19478};
  wire _19480 = _12301 < _19479;
  wire _19481 = r1250 ^ _19480;
  wire _19482 = _12298 ? coded_block[1250] : r1250;
  wire _19483 = _12296 ? _19481 : _19482;
  always @ (posedge reset or posedge clock) if (reset) r1250 <= 1'd0; else if (_12300) r1250 <= _19483;
  wire [1:0] _19484 = {_0, _1088} + {_0, _3901};
  wire [1:0] _19485 = {_0, _5152} + {_0, _7262};
  wire [2:0] _19486 = {_0, _19484} + {_0, _19485};
  wire [1:0] _19487 = {_0, _10108} + {_0, _10846};
  wire [3:0] _19488 = {_0, _19486} + {_0, _0, _19487};
  wire _19489 = _12301 < _19488;
  wire _19490 = r1249 ^ _19489;
  wire _19491 = _12298 ? coded_block[1249] : r1249;
  wire _19492 = _12296 ? _19490 : _19491;
  always @ (posedge reset or posedge clock) if (reset) r1249 <= 1'd0; else if (_12300) r1249 <= _19492;
  wire [1:0] _19493 = {_0, _1120} + {_0, _2175};
  wire [1:0] _19494 = {_0, _5981} + {_0, _7230};
  wire [2:0] _19495 = {_0, _19493} + {_0, _19494};
  wire [1:0] _19496 = {_0, _9342} + {_0, _12188};
  wire [3:0] _19497 = {_0, _19495} + {_0, _0, _19496};
  wire _19498 = _12301 < _19497;
  wire _19499 = r1248 ^ _19498;
  wire _19500 = _12298 ? coded_block[1248] : r1248;
  wire _19501 = _12296 ? _19499 : _19500;
  always @ (posedge reset or posedge clock) if (reset) r1248 <= 1'd0; else if (_12300) r1248 <= _19501;
  wire [1:0] _19502 = {_0, _1151} + {_0, _3580};
  wire [1:0] _19503 = {_0, _4256} + {_0, _8059};
  wire [2:0] _19504 = {_0, _19502} + {_0, _19503};
  wire [1:0] _19505 = {_0, _9311} + {_0, _11422};
  wire [3:0] _19506 = {_0, _19504} + {_0, _0, _19505};
  wire _19507 = _12301 < _19506;
  wire _19508 = r1247 ^ _19507;
  wire _19509 = _12298 ? coded_block[1247] : r1247;
  wire _19510 = _12296 ? _19508 : _19509;
  always @ (posedge reset or posedge clock) if (reset) r1247 <= 1'd0; else if (_12300) r1247 <= _19510;
  wire [1:0] _19511 = {_0, _1184} + {_0, _3422};
  wire [1:0] _19512 = {_0, _5663} + {_0, _6334};
  wire [2:0] _19513 = {_0, _19511} + {_0, _19512};
  wire [1:0] _19514 = {_0, _10141} + {_0, _11389};
  wire [3:0] _19515 = {_0, _19513} + {_0, _0, _19514};
  wire _19516 = _12301 < _19515;
  wire _19517 = r1246 ^ _19516;
  wire _19518 = _12298 ? coded_block[1246] : r1246;
  wire _19519 = _12296 ? _19517 : _19518;
  always @ (posedge reset or posedge clock) if (reset) r1246 <= 1'd0; else if (_12300) r1246 <= _19519;
  wire [1:0] _19520 = {_0, _1215} + {_0, _2081};
  wire [1:0] _19521 = {_0, _5501} + {_0, _7741};
  wire [2:0] _19522 = {_0, _19520} + {_0, _19521};
  wire [1:0] _19523 = {_0, _8415} + {_0, _12219};
  wire [3:0] _19524 = {_0, _19522} + {_0, _0, _19523};
  wire _19525 = _12301 < _19524;
  wire _19526 = r1245 ^ _19525;
  wire _19527 = _12298 ? coded_block[1245] : r1245;
  wire _19528 = _12296 ? _19526 : _19527;
  always @ (posedge reset or posedge clock) if (reset) r1245 <= 1'd0; else if (_12300) r1245 <= _19528;
  wire [1:0] _19529 = {_0, _1247} + {_0, _3453};
  wire [1:0] _19530 = {_0, _4129} + {_0, _7581};
  wire [2:0] _19531 = {_0, _19529} + {_0, _19530};
  wire [1:0] _19532 = {_0, _9822} + {_0, _10493};
  wire [3:0] _19533 = {_0, _19531} + {_0, _0, _19532};
  wire _19534 = _12301 < _19533;
  wire _19535 = r1244 ^ _19534;
  wire _19536 = _12298 ? coded_block[1244] : r1244;
  wire _19537 = _12296 ? _19535 : _19536;
  always @ (posedge reset or posedge clock) if (reset) r1244 <= 1'd0; else if (_12300) r1244 <= _19537;
  wire [1:0] _19538 = {_0, _1278} + {_0, _3646};
  wire [1:0] _19539 = {_0, _5534} + {_0, _6176};
  wire [2:0] _19540 = {_0, _19538} + {_0, _19539};
  wire [1:0] _19541 = {_0, _9661} + {_0, _11900};
  wire [3:0] _19542 = {_0, _19540} + {_0, _0, _19541};
  wire _19543 = _12301 < _19542;
  wire _19544 = r1243 ^ _19543;
  wire _19545 = _12298 ? coded_block[1243] : r1243;
  wire _19546 = _12296 ? _19544 : _19545;
  always @ (posedge reset or posedge clock) if (reset) r1243 <= 1'd0; else if (_12300) r1243 <= _19546;
  wire [1:0] _19547 = {_0, _1312} + {_0, _2271};
  wire [1:0] _19548 = {_0, _5726} + {_0, _7612};
  wire [2:0] _19549 = {_0, _19547} + {_0, _19548};
  wire [1:0] _19550 = {_0, _8225} + {_0, _11740};
  wire [3:0] _19551 = {_0, _19549} + {_0, _0, _19550};
  wire _19552 = _12301 < _19551;
  wire _19553 = r1242 ^ _19552;
  wire _19554 = _12298 ? coded_block[1242] : r1242;
  wire _19555 = _12296 ? _19553 : _19554;
  always @ (posedge reset or posedge clock) if (reset) r1242 <= 1'd0; else if (_12300) r1242 <= _19555;
  wire [1:0] _19556 = {_0, _1375} + {_0, _3231};
  wire [1:0] _19557 = {_0, _6108} + {_0, _6431};
  wire [2:0] _19558 = {_0, _19556} + {_0, _19557};
  wire [1:0] _19559 = {_0, _9886} + {_0, _11771};
  wire [3:0] _19560 = {_0, _19558} + {_0, _0, _19559};
  wire _19561 = _12301 < _19560;
  wire _19562 = r1241 ^ _19561;
  wire _19563 = _12298 ? coded_block[1241] : r1241;
  wire _19564 = _12296 ? _19562 : _19563;
  always @ (posedge reset or posedge clock) if (reset) r1241 <= 1'd0; else if (_12300) r1241 <= _19564;
  wire [1:0] _19565 = {_0, _1439} + {_0, _4091};
  wire [1:0] _19566 = {_0, _5373} + {_0, _7389};
  wire [2:0] _19567 = {_0, _19565} + {_0, _19566};
  wire [1:0] _19568 = {_0, _8256} + {_0, _10590};
  wire [3:0] _19569 = {_0, _19567} + {_0, _0, _19568};
  wire _19570 = _12301 < _19569;
  wire _19571 = r1240 ^ _19570;
  wire _19572 = _12298 ? coded_block[1240] : r1240;
  wire _19573 = _12296 ? _19571 : _19572;
  always @ (posedge reset or posedge clock) if (reset) r1240 <= 1'd0; else if (_12300) r1240 <= _19573;
  wire [1:0] _19574 = {_0, _1502} + {_0, _2686};
  wire [1:0] _19575 = {_0, _4861} + {_0, _6239};
  wire [2:0] _19576 = {_0, _19574} + {_0, _19575};
  wire [1:0] _19577 = {_0, _9534} + {_0, _11550};
  wire [3:0] _19578 = {_0, _19576} + {_0, _0, _19577};
  wire _19579 = _12301 < _19578;
  wire _19580 = r1239 ^ _19579;
  wire _19581 = _12298 ? coded_block[1239] : r1239;
  wire _19582 = _12296 ? _19580 : _19581;
  always @ (posedge reset or posedge clock) if (reset) r1239 <= 1'd0; else if (_12300) r1239 <= _19582;
  wire [1:0] _19583 = {_0, _1533} + {_0, _3198};
  wire [1:0] _19584 = {_0, _4767} + {_0, _6942};
  wire [2:0] _19585 = {_0, _19583} + {_0, _19584};
  wire [1:0] _19586 = {_0, _8319} + {_0, _11613};
  wire [3:0] _19587 = {_0, _19585} + {_0, _0, _19586};
  wire _19588 = _12301 < _19587;
  wire _19589 = r1238 ^ _19588;
  wire _19590 = _12298 ? coded_block[1238] : r1238;
  wire _19591 = _12296 ? _19589 : _19590;
  always @ (posedge reset or posedge clock) if (reset) r1238 <= 1'd0; else if (_12300) r1238 <= _19591;
  wire [1:0] _19592 = {_0, _1568} + {_0, _4060};
  wire [1:0] _19593 = {_0, _5279} + {_0, _6845};
  wire [2:0] _19594 = {_0, _19592} + {_0, _19593};
  wire [1:0] _19595 = {_0, _9022} + {_0, _10399};
  wire [3:0] _19596 = {_0, _19594} + {_0, _0, _19595};
  wire _19597 = _12301 < _19596;
  wire _19598 = r1237 ^ _19597;
  wire _19599 = _12298 ? coded_block[1237] : r1237;
  wire _19600 = _12296 ? _19598 : _19599;
  always @ (posedge reset or posedge clock) if (reset) r1237 <= 1'd0; else if (_12300) r1237 <= _19600;
  wire [1:0] _19601 = {_0, _1599} + {_0, _3325};
  wire [1:0] _19602 = {_0, _6139} + {_0, _7357};
  wire [2:0] _19603 = {_0, _19601} + {_0, _19602};
  wire [1:0] _19604 = {_0, _8926} + {_0, _11101};
  wire [3:0] _19605 = {_0, _19603} + {_0, _0, _19604};
  wire _19606 = _12301 < _19605;
  wire _19607 = r1236 ^ _19606;
  wire _19608 = _12298 ? coded_block[1236] : r1236;
  wire _19609 = _12296 ? _19607 : _19608;
  always @ (posedge reset or posedge clock) if (reset) r1236 <= 1'd0; else if (_12300) r1236 <= _19609;
  wire [1:0] _19610 = {_0, _1631} + {_0, _2367};
  wire [1:0] _19611 = {_0, _5407} + {_0, _6207};
  wire [2:0] _19612 = {_0, _19610} + {_0, _19611};
  wire [1:0] _19613 = {_0, _9438} + {_0, _11004};
  wire [3:0] _19614 = {_0, _19612} + {_0, _0, _19613};
  wire _19615 = _12301 < _19614;
  wire _19616 = r1235 ^ _19615;
  wire _19617 = _12298 ? coded_block[1235] : r1235;
  wire _19618 = _12296 ? _19616 : _19617;
  always @ (posedge reset or posedge clock) if (reset) r1235 <= 1'd0; else if (_12300) r1235 <= _19618;
  wire [1:0] _19619 = {_0, _1695} + {_0, _3997};
  wire [1:0] _19620 = {_0, _4989} + {_0, _6525};
  wire [2:0] _19621 = {_0, _19619} + {_0, _19620};
  wire [1:0] _19622 = {_0, _9566} + {_0, _10366};
  wire [3:0] _19623 = {_0, _19621} + {_0, _0, _19622};
  wire _19624 = _12301 < _19623;
  wire _19625 = r1234 ^ _19624;
  wire _19626 = _12298 ? coded_block[1234] : r1234;
  wire _19627 = _12296 ? _19625 : _19626;
  always @ (posedge reset or posedge clock) if (reset) r1234 <= 1'd0; else if (_12300) r1234 <= _19627;
  wire [1:0] _19628 = {_0, _1726} + {_0, _2302};
  wire [1:0] _19629 = {_0, _6076} + {_0, _7069};
  wire [2:0] _19630 = {_0, _19628} + {_0, _19629};
  wire [1:0] _19631 = {_0, _8607} + {_0, _11644};
  wire [3:0] _19632 = {_0, _19630} + {_0, _0, _19631};
  wire _19633 = _12301 < _19632;
  wire _19634 = r1233 ^ _19633;
  wire _19635 = _12298 ? coded_block[1233] : r1233;
  wire _19636 = _12296 ? _19634 : _19635;
  always @ (posedge reset or posedge clock) if (reset) r1233 <= 1'd0; else if (_12300) r1233 <= _19636;
  wire [1:0] _19637 = {_0, _1758} + {_0, _2750};
  wire [1:0] _19638 = {_0, _4384} + {_0, _8155};
  wire [2:0] _19639 = {_0, _19637} + {_0, _19638};
  wire [1:0] _19640 = {_0, _9149} + {_0, _10685};
  wire [3:0] _19641 = {_0, _19639} + {_0, _0, _19640};
  wire _19642 = _12301 < _19641;
  wire _19643 = r1232 ^ _19642;
  wire _19644 = _12298 ? coded_block[1232] : r1232;
  wire _19645 = _12296 ? _19643 : _19644;
  always @ (posedge reset or posedge clock) if (reset) r1232 <= 1'd0; else if (_12300) r1232 <= _19645;
  wire [1:0] _19646 = {_0, _1789} + {_0, _2112};
  wire [1:0] _19647 = {_0, _4830} + {_0, _6462};
  wire [2:0] _19648 = {_0, _19646} + {_0, _19647};
  wire [1:0] _19649 = {_0, _10235} + {_0, _11228};
  wire [3:0] _19650 = {_0, _19648} + {_0, _0, _19649};
  wire _19651 = _12301 < _19650;
  wire _19652 = r1231 ^ _19651;
  wire _19653 = _12298 ? coded_block[1231] : r1231;
  wire _19654 = _12296 ? _19652 : _19653;
  always @ (posedge reset or posedge clock) if (reset) r1231 <= 1'd0; else if (_12300) r1231 <= _19654;
  wire [1:0] _19655 = {_0, _1823} + {_0, _3037};
  wire [1:0] _19656 = {_0, _4192} + {_0, _6908};
  wire [2:0] _19657 = {_0, _19655} + {_0, _19656};
  wire [1:0] _19658 = {_0, _8543} + {_0, _10303};
  wire [3:0] _19659 = {_0, _19657} + {_0, _0, _19658};
  wire _19660 = _12301 < _19659;
  wire _19661 = r1230 ^ _19660;
  wire _19662 = _12298 ? coded_block[1230] : r1230;
  wire _19663 = _12296 ? _19661 : _19662;
  always @ (posedge reset or posedge clock) if (reset) r1230 <= 1'd0; else if (_12300) r1230 <= _19663;
  wire [1:0] _19664 = {_0, _1854} + {_0, _3135};
  wire [1:0] _19665 = {_0, _5116} + {_0, _6270};
  wire [2:0] _19666 = {_0, _19664} + {_0, _19665};
  wire [1:0] _19667 = {_0, _8991} + {_0, _10621};
  wire [3:0] _19668 = {_0, _19666} + {_0, _0, _19667};
  wire _19669 = _12301 < _19668;
  wire _19670 = r1229 ^ _19669;
  wire _19671 = _12298 ? coded_block[1229] : r1229;
  wire _19672 = _12296 ? _19670 : _19671;
  always @ (posedge reset or posedge clock) if (reset) r1229 <= 1'd0; else if (_12300) r1229 <= _19672;
  wire [1:0] _19673 = {_0, _1886} + {_0, _2592};
  wire [1:0] _19674 = {_0, _5215} + {_0, _7199};
  wire [2:0] _19675 = {_0, _19673} + {_0, _19674};
  wire [1:0] _19676 = {_0, _8352} + {_0, _11069};
  wire [3:0] _19677 = {_0, _19675} + {_0, _0, _19676};
  wire _19678 = _12301 < _19677;
  wire _19679 = r1228 ^ _19678;
  wire _19680 = _12298 ? coded_block[1228] : r1228;
  wire _19681 = _12296 ? _19679 : _19680;
  always @ (posedge reset or posedge clock) if (reset) r1228 <= 1'd0; else if (_12300) r1228 <= _19681;
  wire [1:0] _19682 = {_0, _1917} + {_0, _2847};
  wire [1:0] _19683 = {_0, _4671} + {_0, _7293};
  wire [2:0] _19684 = {_0, _19682} + {_0, _19683};
  wire [1:0] _19685 = {_0, _9279} + {_0, _10430};
  wire [3:0] _19686 = {_0, _19684} + {_0, _0, _19685};
  wire _19687 = _12301 < _19686;
  wire _19688 = r1227 ^ _19687;
  wire _19689 = _12298 ? coded_block[1227] : r1227;
  wire _19690 = _12296 ? _19688 : _19689;
  always @ (posedge reset or posedge clock) if (reset) r1227 <= 1'd0; else if (_12300) r1227 <= _19690;
  wire [1:0] _19691 = {_0, _1950} + {_0, _3742};
  wire [1:0] _19692 = {_0, _4926} + {_0, _6750};
  wire [2:0] _19693 = {_0, _19691} + {_0, _19692};
  wire [1:0] _19694 = {_0, _9375} + {_0, _11358};
  wire [3:0] _19695 = {_0, _19693} + {_0, _0, _19694};
  wire _19696 = _12301 < _19695;
  wire _19697 = r1226 ^ _19696;
  wire _19698 = _12298 ? coded_block[1226] : r1226;
  wire _19699 = _12296 ? _19697 : _19698;
  always @ (posedge reset or posedge clock) if (reset) r1226 <= 1'd0; else if (_12300) r1226 <= _19699;
  wire [1:0] _19700 = {_0, _1981} + {_0, _3390};
  wire [1:0] _19701 = {_0, _5821} + {_0, _7005};
  wire [2:0] _19702 = {_0, _19700} + {_0, _19701};
  wire [1:0] _19703 = {_0, _8830} + {_0, _11453};
  wire [3:0] _19704 = {_0, _19702} + {_0, _0, _19703};
  wire _19705 = _12301 < _19704;
  wire _19706 = r1225 ^ _19705;
  wire _19707 = _12298 ? coded_block[1225] : r1225;
  wire _19708 = _12296 ? _19706 : _19707;
  always @ (posedge reset or posedge clock) if (reset) r1225 <= 1'd0; else if (_12300) r1225 <= _19708;
  wire [1:0] _19709 = {_0, _1470} + {_0, _3742};
  wire [1:0] _19710 = {_0, _6139} + {_0, _6908};
  wire [2:0] _19711 = {_0, _19709} + {_0, _19710};
  wire [1:0] _19712 = {_0, _9566} + {_0, _11165};
  wire [3:0] _19713 = {_0, _19711} + {_0, _0, _19712};
  wire _19714 = _12301 < _19713;
  wire _19715 = r1224 ^ _19714;
  wire _19716 = _12298 ? coded_block[1224] : r1224;
  wire _19717 = _12296 ? _19715 : _19716;
  always @ (posedge reset or posedge clock) if (reset) r1224 <= 1'd0; else if (_12300) r1224 <= _19717;
  wire [1:0] _19718 = {_0, _1502} + {_0, _3901};
  wire [1:0] _19719 = {_0, _5821} + {_0, _6207};
  wire [2:0] _19720 = {_0, _19718} + {_0, _19719};
  wire [1:0] _19721 = {_0, _8991} + {_0, _11644};
  wire [3:0] _19722 = {_0, _19720} + {_0, _0, _19721};
  wire _19723 = _12301 < _19722;
  wire _19724 = r1223 ^ _19723;
  wire _19725 = _12298 ? coded_block[1223] : r1223;
  wire _19726 = _12296 ? _19724 : _19725;
  always @ (posedge reset or posedge clock) if (reset) r1223 <= 1'd0; else if (_12300) r1223 <= _19726;
  wire [1:0] _19727 = {_0, _1533} + {_0, _3709};
  wire [1:0] _19728 = {_0, _5981} + {_0, _7900};
  wire [2:0] _19729 = {_0, _19727} + {_0, _19728};
  wire [1:0] _19730 = {_0, _8288} + {_0, _11069};
  wire [3:0] _19731 = {_0, _19729} + {_0, _0, _19730};
  wire _19732 = _12301 < _19731;
  wire _19733 = r1222 ^ _19732;
  wire _19734 = _12298 ? coded_block[1222] : r1222;
  wire _19735 = _12296 ? _19733 : _19734;
  always @ (posedge reset or posedge clock) if (reset) r1222 <= 1'd0; else if (_12300) r1222 <= _19735;
  wire [1:0] _19736 = {_0, _1568} + {_0, _4091};
  wire [1:0] _19737 = {_0, _5790} + {_0, _8059};
  wire [2:0] _19738 = {_0, _19736} + {_0, _19737};
  wire [1:0] _19739 = {_0, _9980} + {_0, _10366};
  wire [3:0] _19740 = {_0, _19738} + {_0, _0, _19739};
  wire _19741 = _12301 < _19740;
  wire _19742 = r1221 ^ _19741;
  wire _19743 = _12298 ? coded_block[1221] : r1221;
  wire _19744 = _12296 ? _19742 : _19743;
  always @ (posedge reset or posedge clock) if (reset) r1221 <= 1'd0; else if (_12300) r1221 <= _19744;
  wire [1:0] _19745 = {_0, _1599} + {_0, _3231};
  wire [1:0] _19746 = {_0, _4160} + {_0, _7868};
  wire [2:0] _19747 = {_0, _19745} + {_0, _19746};
  wire [1:0] _19748 = {_0, _10141} + {_0, _12061};
  wire [3:0] _19749 = {_0, _19747} + {_0, _0, _19748};
  wire _19750 = _12301 < _19749;
  wire _19751 = r1220 ^ _19750;
  wire _19752 = _12298 ? coded_block[1220] : r1220;
  wire _19753 = _12296 ? _19751 : _19752;
  always @ (posedge reset or posedge clock) if (reset) r1220 <= 1'd0; else if (_12300) r1220 <= _19753;
  wire [1:0] _19754 = {_0, _1631} + {_0, _3005};
  wire [1:0] _19755 = {_0, _5310} + {_0, _6239};
  wire [2:0] _19756 = {_0, _19754} + {_0, _19755};
  wire [1:0] _19757 = {_0, _9949} + {_0, _12219};
  wire [3:0] _19758 = {_0, _19756} + {_0, _0, _19757};
  wire _19759 = _12301 < _19758;
  wire _19760 = r1219 ^ _19759;
  wire _19761 = _12298 ? coded_block[1219] : r1219;
  wire _19762 = _12296 ? _19760 : _19761;
  always @ (posedge reset or posedge clock) if (reset) r1219 <= 1'd0; else if (_12300) r1219 <= _19762;
  wire [1:0] _19763 = {_0, _1662} + {_0, _3580};
  wire [1:0] _19764 = {_0, _5085} + {_0, _7389};
  wire [2:0] _19765 = {_0, _19763} + {_0, _19764};
  wire [1:0] _19766 = {_0, _8319} + {_0, _12027};
  wire [3:0] _19767 = {_0, _19765} + {_0, _0, _19766};
  wire _19768 = _12301 < _19767;
  wire _19769 = r1218 ^ _19768;
  wire _19770 = _12298 ? coded_block[1218] : r1218;
  wire _19771 = _12296 ? _19769 : _19770;
  always @ (posedge reset or posedge clock) if (reset) r1218 <= 1'd0; else if (_12300) r1218 <= _19771;
  wire [1:0] _19772 = {_0, _1439} + {_0, _2750};
  wire [1:0] _19773 = {_0, _6139} + {_0, _7420};
  wire [2:0] _19774 = {_0, _19772} + {_0, _19773};
  wire [1:0] _19775 = {_0, _9438} + {_0, _10303};
  wire [3:0] _19776 = {_0, _19774} + {_0, _0, _19775};
  wire _19777 = _12301 < _19776;
  wire _19778 = r1217 ^ _19777;
  wire _19779 = _12298 ? coded_block[1217] : r1217;
  wire _19780 = _12296 ? _19778 : _19779;
  always @ (posedge reset or posedge clock) if (reset) r1217 <= 1'd0; else if (_12300) r1217 <= _19780;
  wire [1:0] _19781 = {_0, _1470} + {_0, _2655};
  wire [1:0] _19782 = {_0, _4830} + {_0, _6207};
  wire [2:0] _19783 = {_0, _19781} + {_0, _19782};
  wire [1:0] _19784 = {_0, _9503} + {_0, _11516};
  wire [3:0] _19785 = {_0, _19783} + {_0, _0, _19784};
  wire _19786 = _12301 < _19785;
  wire _19787 = r1216 ^ _19786;
  wire _19788 = _12298 ? coded_block[1216] : r1216;
  wire _19789 = _12296 ? _19787 : _19788;
  always @ (posedge reset or posedge clock) if (reset) r1216 <= 1'd0; else if (_12300) r1216 <= _19789;
  wire [1:0] _19790 = {_0, _1502} + {_0, _3167};
  wire [1:0] _19791 = {_0, _4734} + {_0, _6908};
  wire [2:0] _19792 = {_0, _19790} + {_0, _19791};
  wire [1:0] _19793 = {_0, _8288} + {_0, _11581};
  wire [3:0] _19794 = {_0, _19792} + {_0, _0, _19793};
  wire _19795 = _12301 < _19794;
  wire _19796 = r1215 ^ _19795;
  wire _19797 = _12298 ? coded_block[1215] : r1215;
  wire _19798 = _12296 ? _19796 : _19797;
  always @ (posedge reset or posedge clock) if (reset) r1215 <= 1'd0; else if (_12300) r1215 <= _19798;
  wire [1:0] _19799 = {_0, _1599} + {_0, _2336};
  wire [1:0] _19800 = {_0, _5373} + {_0, _8186};
  wire [2:0] _19801 = {_0, _19799} + {_0, _19800};
  wire [1:0] _19802 = {_0, _9406} + {_0, _10973};
  wire [3:0] _19803 = {_0, _19801} + {_0, _0, _19802};
  wire _19804 = _12301 < _19803;
  wire _19805 = r1214 ^ _19804;
  wire _19806 = _12298 ? coded_block[1214] : r1214;
  wire _19807 = _12296 ? _19805 : _19806;
  always @ (posedge reset or posedge clock) if (reset) r1214 <= 1'd0; else if (_12300) r1214 <= _19807;
  wire [1:0] _19808 = {_0, _1631} + {_0, _2878};
  wire [1:0] _19809 = {_0, _4415} + {_0, _7454};
  wire [2:0] _19810 = {_0, _19808} + {_0, _19809};
  wire [1:0] _19811 = {_0, _8256} + {_0, _11485};
  wire [3:0] _19812 = {_0, _19810} + {_0, _0, _19811};
  wire _19813 = _12301 < _19812;
  wire _19814 = r1213 ^ _19813;
  wire _19815 = _12298 ? coded_block[1213] : r1213;
  wire _19816 = _12296 ? _19814 : _19815;
  always @ (posedge reset or posedge clock) if (reset) r1213 <= 1'd0; else if (_12300) r1213 <= _19816;
  wire [1:0] _19817 = {_0, _1695} + {_0, _2271};
  wire [1:0] _19818 = {_0, _6045} + {_0, _7036};
  wire [2:0] _19819 = {_0, _19817} + {_0, _19818};
  wire [1:0] _19820 = {_0, _8574} + {_0, _11613};
  wire [3:0] _19821 = {_0, _19819} + {_0, _0, _19820};
  wire _19822 = _12301 < _19821;
  wire _19823 = r1212 ^ _19822;
  wire _19824 = _12298 ? coded_block[1212] : r1212;
  wire _19825 = _12296 ? _19823 : _19824;
  always @ (posedge reset or posedge clock) if (reset) r1212 <= 1'd0; else if (_12300) r1212 <= _19825;
  wire [1:0] _19826 = {_0, _1726} + {_0, _2719};
  wire [1:0] _19827 = {_0, _4350} + {_0, _8123};
  wire [2:0] _19828 = {_0, _19826} + {_0, _19827};
  wire [1:0] _19829 = {_0, _9118} + {_0, _10654};
  wire [3:0] _19830 = {_0, _19828} + {_0, _0, _19829};
  wire _19831 = _12301 < _19830;
  wire _19832 = r1211 ^ _19831;
  wire _19833 = _12298 ? coded_block[1211] : r1211;
  wire _19834 = _12296 ? _19832 : _19833;
  always @ (posedge reset or posedge clock) if (reset) r1211 <= 1'd0; else if (_12300) r1211 <= _19834;
  wire [1:0] _19835 = {_0, _1758} + {_0, _4091};
  wire [1:0] _19836 = {_0, _4798} + {_0, _6431};
  wire [2:0] _19837 = {_0, _19835} + {_0, _19836};
  wire [1:0] _19838 = {_0, _10204} + {_0, _11196};
  wire [3:0] _19839 = {_0, _19837} + {_0, _0, _19838};
  wire _19840 = _12301 < _19839;
  wire _19841 = r1210 ^ _19840;
  wire _19842 = _12298 ? coded_block[1210] : r1210;
  wire _19843 = _12296 ? _19841 : _19842;
  always @ (posedge reset or posedge clock) if (reset) r1210 <= 1'd0; else if (_12300) r1210 <= _19843;
  wire [1:0] _19844 = {_0, _1789} + {_0, _3005};
  wire [1:0] _19845 = {_0, _4160} + {_0, _6877};
  wire [2:0] _19846 = {_0, _19844} + {_0, _19845};
  wire [1:0] _19847 = {_0, _8511} + {_0, _12282};
  wire [3:0] _19848 = {_0, _19846} + {_0, _0, _19847};
  wire _19849 = _12301 < _19848;
  wire _19850 = r1209 ^ _19849;
  wire _19851 = _12298 ? coded_block[1209] : r1209;
  wire _19852 = _12296 ? _19850 : _19851;
  always @ (posedge reset or posedge clock) if (reset) r1209 <= 1'd0; else if (_12300) r1209 <= _19852;
  wire [1:0] _19853 = {_0, _1823} + {_0, _3104};
  wire [1:0] _19854 = {_0, _5085} + {_0, _6239};
  wire [2:0] _19855 = {_0, _19853} + {_0, _19854};
  wire [1:0] _19856 = {_0, _8957} + {_0, _10590};
  wire [3:0] _19857 = {_0, _19855} + {_0, _0, _19856};
  wire _19858 = _12301 < _19857;
  wire _19859 = r1208 ^ _19858;
  wire _19860 = _12298 ? coded_block[1208] : r1208;
  wire _19861 = _12296 ? _19859 : _19860;
  always @ (posedge reset or posedge clock) if (reset) r1208 <= 1'd0; else if (_12300) r1208 <= _19861;
  wire [1:0] _19862 = {_0, _1854} + {_0, _2557};
  wire [1:0] _19863 = {_0, _5183} + {_0, _7163};
  wire [2:0] _19864 = {_0, _19862} + {_0, _19863};
  wire [1:0] _19865 = {_0, _8319} + {_0, _11038};
  wire [3:0] _19866 = {_0, _19864} + {_0, _0, _19865};
  wire _19867 = _12301 < _19866;
  wire _19868 = r1207 ^ _19867;
  wire _19869 = _12298 ? coded_block[1207] : r1207;
  wire _19870 = _12296 ? _19868 : _19869;
  always @ (posedge reset or posedge clock) if (reset) r1207 <= 1'd0; else if (_12300) r1207 <= _19870;
  wire [1:0] _19871 = {_0, _1886} + {_0, _2813};
  wire [1:0] _19872 = {_0, _4640} + {_0, _7262};
  wire [2:0] _19873 = {_0, _19871} + {_0, _19872};
  wire [1:0] _19874 = {_0, _9248} + {_0, _10399};
  wire [3:0] _19875 = {_0, _19873} + {_0, _0, _19874};
  wire _19876 = _12301 < _19875;
  wire _19877 = r1206 ^ _19876;
  wire _19878 = _12298 ? coded_block[1206] : r1206;
  wire _19879 = _12296 ? _19877 : _19878;
  always @ (posedge reset or posedge clock) if (reset) r1206 <= 1'd0; else if (_12300) r1206 <= _19879;
  wire [1:0] _19880 = {_0, _1917} + {_0, _3709};
  wire [1:0] _19881 = {_0, _4895} + {_0, _6718};
  wire [2:0] _19882 = {_0, _19880} + {_0, _19881};
  wire [1:0] _19883 = {_0, _9342} + {_0, _11326};
  wire [3:0] _19884 = {_0, _19882} + {_0, _0, _19883};
  wire _19885 = _12301 < _19884;
  wire _19886 = r1205 ^ _19885;
  wire _19887 = _12298 ? coded_block[1205] : r1205;
  wire _19888 = _12296 ? _19886 : _19887;
  always @ (posedge reset or posedge clock) if (reset) r1205 <= 1'd0; else if (_12300) r1205 <= _19888;
  wire [1:0] _19889 = {_0, _1950} + {_0, _3359};
  wire [1:0] _19890 = {_0, _5790} + {_0, _6973};
  wire [2:0] _19891 = {_0, _19889} + {_0, _19890};
  wire [1:0] _19892 = {_0, _8799} + {_0, _11422};
  wire [3:0] _19893 = {_0, _19891} + {_0, _0, _19892};
  wire _19894 = _12301 < _19893;
  wire _19895 = r1204 ^ _19894;
  wire _19896 = _12298 ? coded_block[1204] : r1204;
  wire _19897 = _12296 ? _19895 : _19896;
  always @ (posedge reset or posedge clock) if (reset) r1204 <= 1'd0; else if (_12300) r1204 <= _19897;
  wire [1:0] _19898 = {_0, _1981} + {_0, _3580};
  wire [1:0] _19899 = {_0, _5438} + {_0, _7868};
  wire [2:0] _19900 = {_0, _19898} + {_0, _19899};
  wire [1:0] _19901 = {_0, _9054} + {_0, _10877};
  wire [3:0] _19902 = {_0, _19900} + {_0, _0, _19901};
  wire _19903 = _12301 < _19902;
  wire _19904 = r1203 ^ _19903;
  wire _19905 = _12298 ? coded_block[1203] : r1203;
  wire _19906 = _12296 ? _19904 : _19905;
  always @ (posedge reset or posedge clock) if (reset) r1203 <= 1'd0; else if (_12300) r1203 <= _19906;
  wire [1:0] _19907 = {_0, _2013} + {_0, _3453};
  wire [1:0] _19908 = {_0, _5663} + {_0, _7517};
  wire [2:0] _19909 = {_0, _19907} + {_0, _19908};
  wire [1:0] _19910 = {_0, _9949} + {_0, _11132};
  wire [3:0] _19911 = {_0, _19909} + {_0, _0, _19910};
  wire _19912 = _12301 < _19911;
  wire _19913 = r1202 ^ _19912;
  wire _19914 = _12298 ? coded_block[1202] : r1202;
  wire _19915 = _12296 ? _19913 : _19914;
  always @ (posedge reset or posedge clock) if (reset) r1202 <= 1'd0; else if (_12300) r1202 <= _19915;
  wire [1:0] _19916 = {_0, _2044} + {_0, _3805};
  wire [1:0] _19917 = {_0, _5534} + {_0, _7741};
  wire [2:0] _19918 = {_0, _19916} + {_0, _19917};
  wire [1:0] _19919 = {_0, _9597} + {_0, _12027};
  wire [3:0] _19920 = {_0, _19918} + {_0, _0, _19919};
  wire _19921 = _12301 < _19920;
  wire _19922 = r1201 ^ _19921;
  wire _19923 = _12298 ? coded_block[1201] : r1201;
  wire _19924 = _12296 ? _19922 : _19923;
  always @ (posedge reset or posedge clock) if (reset) r1201 <= 1'd0; else if (_12300) r1201 <= _19924;
  wire [1:0] _19925 = {_0, _65} + {_0, _2526};
  wire [1:0] _19926 = {_0, _5884} + {_0, _7612};
  wire [2:0] _19927 = {_0, _19925} + {_0, _19926};
  wire [1:0] _19928 = {_0, _9822} + {_0, _11677};
  wire [3:0] _19929 = {_0, _19927} + {_0, _0, _19928};
  wire _19930 = _12301 < _19929;
  wire _19931 = r1200 ^ _19930;
  wire _19932 = _12298 ? coded_block[1200] : r1200;
  wire _19933 = _12296 ? _19931 : _19932;
  always @ (posedge reset or posedge clock) if (reset) r1200 <= 1'd0; else if (_12300) r1200 <= _19933;
  wire [1:0] _19934 = {_0, _97} + {_0, _3135};
  wire [1:0] _19935 = {_0, _4605} + {_0, _7965};
  wire [2:0] _19936 = {_0, _19934} + {_0, _19935};
  wire [1:0] _19937 = {_0, _9693} + {_0, _11900};
  wire [3:0] _19938 = {_0, _19936} + {_0, _0, _19937};
  wire _19939 = _12301 < _19938;
  wire _19940 = r1199 ^ _19939;
  wire _19941 = _12298 ? coded_block[1199] : r1199;
  wire _19942 = _12296 ? _19940 : _19941;
  always @ (posedge reset or posedge clock) if (reset) r1199 <= 1'd0; else if (_12300) r1199 <= _19942;
  wire [1:0] _19943 = {_0, _161} + {_0, _2302};
  wire [1:0] _19944 = {_0, _4767} + {_0, _7293};
  wire [2:0] _19945 = {_0, _19943} + {_0, _19944};
  wire [1:0] _19946 = {_0, _8767} + {_0, _12124};
  wire [3:0] _19947 = {_0, _19945} + {_0, _0, _19946};
  wire _19948 = _12301 < _19947;
  wire _19949 = r1198 ^ _19948;
  wire _19950 = _12298 ? coded_block[1198] : r1198;
  wire _19951 = _12296 ? _19949 : _19950;
  always @ (posedge reset or posedge clock) if (reset) r1198 <= 1'd0; else if (_12300) r1198 <= _19951;
  wire [1:0] _19952 = {_0, _192} + {_0, _3325};
  wire [1:0] _19953 = {_0, _4384} + {_0, _6845};
  wire [2:0] _19954 = {_0, _19952} + {_0, _19953};
  wire [1:0] _19955 = {_0, _9375} + {_0, _10846};
  wire [3:0] _19956 = {_0, _19954} + {_0, _0, _19955};
  wire _19957 = _12301 < _19956;
  wire _19958 = r1197 ^ _19957;
  wire _19959 = _12298 ? coded_block[1197] : r1197;
  wire _19960 = _12296 ? _19958 : _19959;
  always @ (posedge reset or posedge clock) if (reset) r1197 <= 1'd0; else if (_12300) r1197 <= _19960;
  wire [1:0] _19961 = {_0, _224} + {_0, _3742};
  wire [1:0] _19962 = {_0, _5407} + {_0, _6462};
  wire [2:0] _19963 = {_0, _19961} + {_0, _19962};
  wire [1:0] _19964 = {_0, _8926} + {_0, _11453};
  wire [3:0] _19965 = {_0, _19963} + {_0, _0, _19964};
  wire _19966 = _12301 < _19965;
  wire _19967 = r1196 ^ _19966;
  wire _19968 = _12298 ? coded_block[1196] : r1196;
  wire _19969 = _12296 ? _19967 : _19968;
  always @ (posedge reset or posedge clock) if (reset) r1196 <= 1'd0; else if (_12300) r1196 <= _19969;
  wire [1:0] _19970 = {_0, _255} + {_0, _2208};
  wire [1:0] _19971 = {_0, _5821} + {_0, _7485};
  wire [2:0] _19972 = {_0, _19970} + {_0, _19971};
  wire [1:0] _19973 = {_0, _8543} + {_0, _11004};
  wire [3:0] _19974 = {_0, _19972} + {_0, _0, _19973};
  wire _19975 = _12301 < _19974;
  wire _19976 = r1195 ^ _19975;
  wire _19977 = _12298 ? coded_block[1195] : r1195;
  wire _19978 = _12296 ? _19976 : _19977;
  always @ (posedge reset or posedge clock) if (reset) r1195 <= 1'd0; else if (_12300) r1195 <= _19978;
  wire [1:0] _19979 = {_0, _289} + {_0, _3646};
  wire [1:0] _19980 = {_0, _4287} + {_0, _7900};
  wire [2:0] _19981 = {_0, _19979} + {_0, _19980};
  wire [1:0] _19982 = {_0, _9566} + {_0, _10621};
  wire [3:0] _19983 = {_0, _19981} + {_0, _0, _19982};
  wire _19984 = _12301 < _19983;
  wire _19985 = r1194 ^ _19984;
  wire _19986 = _12298 ? coded_block[1194] : r1194;
  wire _19987 = _12296 ? _19985 : _19986;
  always @ (posedge reset or posedge clock) if (reset) r1194 <= 1'd0; else if (_12300) r1194 <= _19987;
  wire [1:0] _19988 = {_0, _320} + {_0, _2941};
  wire [1:0] _19989 = {_0, _5726} + {_0, _6366};
  wire [2:0] _19990 = {_0, _19988} + {_0, _19989};
  wire [1:0] _19991 = {_0, _9980} + {_0, _11644};
  wire [3:0] _19992 = {_0, _19990} + {_0, _0, _19991};
  wire _19993 = _12301 < _19992;
  wire _19994 = r1193 ^ _19993;
  wire _19995 = _12298 ? coded_block[1193] : r1193;
  wire _19996 = _12296 ? _19994 : _19995;
  always @ (posedge reset or posedge clock) if (reset) r1193 <= 1'd0; else if (_12300) r1193 <= _19996;
  wire [1:0] _19997 = {_0, _416} + {_0, _2592};
  wire [1:0] _19998 = {_0, _4861} + {_0, _6781};
  wire [2:0] _19999 = {_0, _19997} + {_0, _19998};
  wire [1:0] _20000 = {_0, _9181} + {_0, _11964};
  wire [3:0] _20001 = {_0, _19999} + {_0, _0, _20000};
  wire _20002 = _12301 < _20001;
  wire _20003 = r1192 ^ _20002;
  wire _20004 = _12298 ? coded_block[1192] : r1192;
  wire _20005 = _12296 ? _20003 : _20004;
  always @ (posedge reset or posedge clock) if (reset) r1192 <= 1'd0; else if (_12300) r1192 <= _20005;
  wire [1:0] _20006 = {_0, _447} + {_0, _2974};
  wire [1:0] _20007 = {_0, _4671} + {_0, _6942};
  wire [2:0] _20008 = {_0, _20006} + {_0, _20007};
  wire [1:0] _20009 = {_0, _8863} + {_0, _11259};
  wire [3:0] _20010 = {_0, _20008} + {_0, _0, _20009};
  wire _20011 = _12301 < _20010;
  wire _20012 = r1191 ^ _20011;
  wire _20013 = _12298 ? coded_block[1191] : r1191;
  wire _20014 = _12296 ? _20012 : _20013;
  always @ (posedge reset or posedge clock) if (reset) r1191 <= 1'd0; else if (_12300) r1191 <= _20014;
  wire [1:0] _20015 = {_0, _479} + {_0, _2112};
  wire [1:0] _20016 = {_0, _5053} + {_0, _6750};
  wire [2:0] _20017 = {_0, _20015} + {_0, _20016};
  wire [1:0] _20018 = {_0, _9022} + {_0, _10941};
  wire [3:0] _20019 = {_0, _20017} + {_0, _0, _20018};
  wire _20020 = _12301 < _20019;
  wire _20021 = r1190 ^ _20020;
  wire _20022 = _12298 ? coded_block[1190] : r1190;
  wire _20023 = _12296 ? _20021 : _20022;
  always @ (posedge reset or posedge clock) if (reset) r1190 <= 1'd0; else if (_12300) r1190 <= _20023;
  wire [1:0] _20024 = {_0, _510} + {_0, _3901};
  wire [1:0] _20025 = {_0, _4192} + {_0, _7132};
  wire [2:0] _20026 = {_0, _20024} + {_0, _20025};
  wire [1:0] _20027 = {_0, _8830} + {_0, _11101};
  wire [3:0] _20028 = {_0, _20026} + {_0, _0, _20027};
  wire _20029 = _12301 < _20028;
  wire _20030 = r1189 ^ _20029;
  wire _20031 = _12298 ? coded_block[1189] : r1189;
  wire _20032 = _12296 ? _20030 : _20031;
  always @ (posedge reset or posedge clock) if (reset) r1189 <= 1'd0; else if (_12300) r1189 <= _20032;
  wire [1:0] _20033 = {_0, _545} + {_0, _2463};
  wire [1:0] _20034 = {_0, _5981} + {_0, _6270};
  wire [2:0] _20035 = {_0, _20033} + {_0, _20034};
  wire [1:0] _20036 = {_0, _9212} + {_0, _10910};
  wire [3:0] _20037 = {_0, _20035} + {_0, _0, _20036};
  wire _20038 = _12301 < _20037;
  wire _20039 = r1188 ^ _20038;
  wire _20040 = _12298 ? coded_block[1188] : r1188;
  wire _20041 = _12296 ? _20039 : _20040;
  always @ (posedge reset or posedge clock) if (reset) r1188 <= 1'd0; else if (_12300) r1188 <= _20041;
  wire [1:0] _20042 = {_0, _576} + {_0, _2399};
  wire [1:0] _20043 = {_0, _4542} + {_0, _8059};
  wire [2:0] _20044 = {_0, _20042} + {_0, _20043};
  wire [1:0] _20045 = {_0, _8352} + {_0, _11295};
  wire [3:0] _20046 = {_0, _20044} + {_0, _0, _20045};
  wire _20047 = _12301 < _20046;
  wire _20048 = r1187 ^ _20047;
  wire _20049 = _12298 ? coded_block[1187] : r1187;
  wire _20050 = _12296 ? _20048 : _20049;
  always @ (posedge reset or posedge clock) if (reset) r1187 <= 1'd0; else if (_12300) r1187 <= _20050;
  wire [1:0] _20051 = {_0, _608} + {_0, _3517};
  wire [1:0] _20052 = {_0, _4478} + {_0, _6621};
  wire [2:0] _20053 = {_0, _20051} + {_0, _20052};
  wire [1:0] _20054 = {_0, _10141} + {_0, _10430};
  wire [3:0] _20055 = {_0, _20053} + {_0, _0, _20054};
  wire _20056 = _12301 < _20055;
  wire _20057 = r1186 ^ _20056;
  wire _20058 = _12298 ? coded_block[1186] : r1186;
  wire _20059 = _12296 ? _20057 : _20058;
  always @ (posedge reset or posedge clock) if (reset) r1186 <= 1'd0; else if (_12300) r1186 <= _20059;
  wire [1:0] _20060 = {_0, _672} + {_0, _3773};
  wire [1:0] _20061 = {_0, _4256} + {_0, _7675};
  wire [2:0] _20062 = {_0, _20060} + {_0, _20061};
  wire [1:0] _20063 = {_0, _8638} + {_0, _10783};
  wire [3:0] _20064 = {_0, _20062} + {_0, _0, _20063};
  wire _20065 = _12301 < _20064;
  wire _20066 = r1185 ^ _20065;
  wire _20067 = _12298 ? coded_block[1185] : r1185;
  wire _20068 = _12296 ? _20066 : _20067;
  always @ (posedge reset or posedge clock) if (reset) r1185 <= 1'd0; else if (_12300) r1185 <= _20068;
  wire [1:0] _20069 = {_0, _703} + {_0, _3486};
  wire [1:0] _20070 = {_0, _5853} + {_0, _6334};
  wire [2:0] _20071 = {_0, _20069} + {_0, _20070};
  wire [1:0] _20072 = {_0, _9759} + {_0, _10717};
  wire [3:0] _20073 = {_0, _20071} + {_0, _0, _20072};
  wire _20074 = _12301 < _20073;
  wire _20075 = r1184 ^ _20074;
  wire _20076 = _12298 ? coded_block[1184] : r1184;
  wire _20077 = _12296 ? _20075 : _20076;
  always @ (posedge reset or posedge clock) if (reset) r1184 <= 1'd0; else if (_12300) r1184 <= _20077;
  wire [1:0] _20078 = {_0, _735} + {_0, _2430};
  wire [1:0] _20079 = {_0, _5565} + {_0, _7931};
  wire [2:0] _20080 = {_0, _20078} + {_0, _20079};
  wire [1:0] _20081 = {_0, _8415} + {_0, _11837};
  wire [3:0] _20082 = {_0, _20080} + {_0, _0, _20081};
  wire _20083 = _12301 < _20082;
  wire _20084 = r1183 ^ _20083;
  wire _20085 = _12298 ? coded_block[1183] : r1183;
  wire _20086 = _12296 ? _20084 : _20085;
  always @ (posedge reset or posedge clock) if (reset) r1183 <= 1'd0; else if (_12300) r1183 <= _20086;
  wire [1:0] _20087 = {_0, _766} + {_0, _3933};
  wire [1:0] _20088 = {_0, _4511} + {_0, _7644};
  wire [2:0] _20089 = {_0, _20087} + {_0, _20088};
  wire [1:0] _20090 = {_0, _10014} + {_0, _10493};
  wire [3:0] _20091 = {_0, _20089} + {_0, _0, _20090};
  wire _20092 = _12301 < _20091;
  wire _20093 = r1182 ^ _20092;
  wire _20094 = _12298 ? coded_block[1182] : r1182;
  wire _20095 = _12296 ? _20093 : _20094;
  always @ (posedge reset or posedge clock) if (reset) r1182 <= 1'd0; else if (_12300) r1182 <= _20095;
  wire [1:0] _20096 = {_0, _800} + {_0, _2910};
  wire [1:0] _20097 = {_0, _6012} + {_0, _6589};
  wire [2:0] _20098 = {_0, _20096} + {_0, _20097};
  wire [1:0] _20099 = {_0, _9724} + {_0, _12092};
  wire [3:0] _20100 = {_0, _20098} + {_0, _0, _20099};
  wire _20101 = _12301 < _20100;
  wire _20102 = r1181 ^ _20101;
  wire _20103 = _12298 ? coded_block[1181] : r1181;
  wire _20104 = _12296 ? _20102 : _20103;
  always @ (posedge reset or posedge clock) if (reset) r1181 <= 1'd0; else if (_12300) r1181 <= _20104;
  wire [1:0] _20105 = {_0, _831} + {_0, _3678};
  wire [1:0] _20106 = {_0, _4989} + {_0, _8092};
  wire [2:0] _20107 = {_0, _20105} + {_0, _20106};
  wire [1:0] _20108 = {_0, _8670} + {_0, _11806};
  wire [3:0] _20109 = {_0, _20107} + {_0, _0, _20108};
  wire _20110 = _12301 < _20109;
  wire _20111 = r1180 ^ _20110;
  wire _20112 = _12298 ? coded_block[1180] : r1180;
  wire _20113 = _12296 ? _20111 : _20112;
  always @ (posedge reset or posedge clock) if (reset) r1180 <= 1'd0; else if (_12300) r1180 <= _20113;
  wire [1:0] _20114 = {_0, _863} + {_0, _2847};
  wire [1:0] _20115 = {_0, _5757} + {_0, _7069};
  wire [2:0] _20116 = {_0, _20114} + {_0, _20115};
  wire [1:0] _20117 = {_0, _10172} + {_0, _10748};
  wire [3:0] _20118 = {_0, _20116} + {_0, _0, _20117};
  wire _20119 = _12301 < _20118;
  wire _20120 = r1179 ^ _20119;
  wire _20121 = _12298 ? coded_block[1179] : r1179;
  wire _20122 = _12296 ? _20120 : _20121;
  always @ (posedge reset or posedge clock) if (reset) r1179 <= 1'd0; else if (_12300) r1179 <= _20122;
  wire [1:0] _20123 = {_0, _894} + {_0, _2367};
  wire [1:0] _20124 = {_0, _4926} + {_0, _7837};
  wire [2:0] _20125 = {_0, _20123} + {_0, _20124};
  wire [1:0] _20126 = {_0, _9149} + {_0, _12251};
  wire [3:0] _20127 = {_0, _20125} + {_0, _0, _20126};
  wire _20128 = _12301 < _20127;
  wire _20129 = r1178 ^ _20128;
  wire _20130 = _12298 ? coded_block[1178] : r1178;
  wire _20131 = _12296 ? _20129 : _20130;
  always @ (posedge reset or posedge clock) if (reset) r1178 <= 1'd0; else if (_12300) r1178 <= _20131;
  wire [1:0] _20132 = {_0, _927} + {_0, _2494};
  wire [1:0] _20133 = {_0, _4447} + {_0, _7005};
  wire [2:0] _20134 = {_0, _20132} + {_0, _20133};
  wire [1:0] _20135 = {_0, _9917} + {_0, _11228};
  wire [3:0] _20136 = {_0, _20134} + {_0, _0, _20135};
  wire _20137 = _12301 < _20136;
  wire _20138 = r1177 ^ _20137;
  wire _20139 = _12298 ? coded_block[1177] : r1177;
  wire _20140 = _12296 ? _20138 : _20139;
  always @ (posedge reset or posedge clock) if (reset) r1177 <= 1'd0; else if (_12300) r1177 <= _20140;
  wire [1:0] _20141 = {_0, _990} + {_0, _3068};
  wire [1:0] _20142 = {_0, _5918} + {_0, _6652};
  wire [2:0] _20143 = {_0, _20141} + {_0, _20142};
  wire [1:0] _20144 = {_0, _8607} + {_0, _11165};
  wire [3:0] _20145 = {_0, _20143} + {_0, _0, _20144};
  wire _20146 = _12301 < _20145;
  wire _20147 = r1176 ^ _20146;
  wire _20148 = _12298 ? coded_block[1176] : r1176;
  wire _20149 = _12296 ? _20147 : _20148;
  always @ (posedge reset or posedge clock) if (reset) r1176 <= 1'd0; else if (_12300) r1176 <= _20149;
  wire [1:0] _20150 = {_0, _1021} + {_0, _3037};
  wire [1:0] _20151 = {_0, _5152} + {_0, _7996};
  wire [2:0] _20152 = {_0, _20150} + {_0, _20151};
  wire [1:0] _20153 = {_0, _8736} + {_0, _10685};
  wire [3:0] _20154 = {_0, _20152} + {_0, _0, _20153};
  wire _20155 = _12301 < _20154;
  wire _20156 = r1175 ^ _20155;
  wire _20157 = _12298 ? coded_block[1175] : r1175;
  wire _20158 = _12296 ? _20156 : _20157;
  always @ (posedge reset or posedge clock) if (reset) r1175 <= 1'd0; else if (_12300) r1175 <= _20158;
  wire [1:0] _20159 = {_0, _1088} + {_0, _2144};
  wire [1:0] _20160 = {_0, _5949} + {_0, _7199};
  wire [2:0] _20161 = {_0, _20159} + {_0, _20160};
  wire [1:0] _20162 = {_0, _9311} + {_0, _12155};
  wire [3:0] _20163 = {_0, _20161} + {_0, _0, _20162};
  wire _20164 = _12301 < _20163;
  wire _20165 = r1174 ^ _20164;
  wire _20166 = _12298 ? coded_block[1174] : r1174;
  wire _20167 = _12296 ? _20165 : _20166;
  always @ (posedge reset or posedge clock) if (reset) r1174 <= 1'd0; else if (_12300) r1174 <= _20167;
  wire [1:0] _20168 = {_0, _1120} + {_0, _3549};
  wire [1:0] _20169 = {_0, _4223} + {_0, _8028};
  wire [2:0] _20170 = {_0, _20168} + {_0, _20169};
  wire [1:0] _20171 = {_0, _9279} + {_0, _11389};
  wire [3:0] _20172 = {_0, _20170} + {_0, _0, _20171};
  wire _20173 = _12301 < _20172;
  wire _20174 = r1173 ^ _20173;
  wire _20175 = _12298 ? coded_block[1173] : r1173;
  wire _20176 = _12296 ? _20174 : _20175;
  always @ (posedge reset or posedge clock) if (reset) r1173 <= 1'd0; else if (_12300) r1173 <= _20176;
  wire [1:0] _20177 = {_0, _1151} + {_0, _3390};
  wire [1:0] _20178 = {_0, _5628} + {_0, _6303};
  wire [2:0] _20179 = {_0, _20177} + {_0, _20178};
  wire [1:0] _20180 = {_0, _10108} + {_0, _11358};
  wire [3:0] _20181 = {_0, _20179} + {_0, _0, _20180};
  wire _20182 = _12301 < _20181;
  wire _20183 = r1172 ^ _20182;
  wire _20184 = _12298 ? coded_block[1172] : r1172;
  wire _20185 = _12296 ? _20183 : _20184;
  always @ (posedge reset or posedge clock) if (reset) r1172 <= 1'd0; else if (_12300) r1172 <= _20185;
  wire [1:0] _20186 = {_0, _1184} + {_0, _2081};
  wire [1:0] _20187 = {_0, _5470} + {_0, _7710};
  wire [2:0] _20188 = {_0, _20186} + {_0, _20187};
  wire [1:0] _20189 = {_0, _8383} + {_0, _12188};
  wire [3:0] _20190 = {_0, _20188} + {_0, _0, _20189};
  wire _20191 = _12301 < _20190;
  wire _20192 = r1171 ^ _20191;
  wire _20193 = _12298 ? coded_block[1171] : r1171;
  wire _20194 = _12296 ? _20192 : _20193;
  always @ (posedge reset or posedge clock) if (reset) r1171 <= 1'd0; else if (_12300) r1171 <= _20194;
  wire [1:0] _20195 = {_0, _1215} + {_0, _3422};
  wire [1:0] _20196 = {_0, _4129} + {_0, _7548};
  wire [2:0] _20197 = {_0, _20195} + {_0, _20196};
  wire [1:0] _20198 = {_0, _9790} + {_0, _10462};
  wire [3:0] _20199 = {_0, _20197} + {_0, _0, _20198};
  wire _20200 = _12301 < _20199;
  wire _20201 = r1170 ^ _20200;
  wire _20202 = _12298 ? coded_block[1170] : r1170;
  wire _20203 = _12296 ? _20201 : _20202;
  always @ (posedge reset or posedge clock) if (reset) r1170 <= 1'd0; else if (_12300) r1170 <= _20203;
  wire [1:0] _20204 = {_0, _1695} + {_0, _3517};
  wire [1:0] _20205 = {_0, _5663} + {_0, _7163};
  wire [2:0] _20206 = {_0, _20204} + {_0, _20205};
  wire [1:0] _20207 = {_0, _9469} + {_0, _10399};
  wire [3:0] _20208 = {_0, _20206} + {_0, _0, _20207};
  wire _20209 = _12301 < _20208;
  wire _20210 = r1169 ^ _20209;
  wire _20211 = _12298 ? coded_block[1169] : r1169;
  wire _20212 = _12296 ? _20210 : _20211;
  always @ (posedge reset or posedge clock) if (reset) r1169 <= 1'd0; else if (_12300) r1169 <= _20212;
  wire [1:0] _20213 = {_0, _1726} + {_0, _2623};
  wire [1:0] _20214 = {_0, _5597} + {_0, _7741};
  wire [2:0] _20215 = {_0, _20213} + {_0, _20214};
  wire [1:0] _20216 = {_0, _9248} + {_0, _11550};
  wire [3:0] _20217 = {_0, _20215} + {_0, _0, _20216};
  wire _20218 = _12301 < _20217;
  wire _20219 = r1168 ^ _20218;
  wire _20220 = _12298 ? coded_block[1168] : r1168;
  wire _20221 = _12296 ? _20219 : _20220;
  always @ (posedge reset or posedge clock) if (reset) r1168 <= 1'd0; else if (_12300) r1168 <= _20221;
  wire [1:0] _20222 = {_0, _1789} + {_0, _2878};
  wire [1:0] _20223 = {_0, _5373} + {_0, _6781};
  wire [2:0] _20224 = {_0, _20222} + {_0, _20223};
  wire [1:0] _20225 = {_0, _9759} + {_0, _11900};
  wire [3:0] _20226 = {_0, _20224} + {_0, _0, _20225};
  wire _20227 = _12301 < _20226;
  wire _20228 = r1167 ^ _20227;
  wire _20229 = _12298 ? coded_block[1167] : r1167;
  wire _20230 = _12296 ? _20228 : _20229;
  always @ (posedge reset or posedge clock) if (reset) r1167 <= 1'd0; else if (_12300) r1167 <= _20230;
  wire [1:0] _20231 = {_0, _1823} + {_0, _2592};
  wire [1:0] _20232 = {_0, _4958} + {_0, _7454};
  wire [2:0] _20233 = {_0, _20231} + {_0, _20232};
  wire [1:0] _20234 = {_0, _8863} + {_0, _11837};
  wire [3:0] _20235 = {_0, _20233} + {_0, _0, _20234};
  wire _20236 = _12301 < _20235;
  wire _20237 = r1166 ^ _20236;
  wire _20238 = _12298 ? coded_block[1166] : r1166;
  wire _20239 = _12296 ? _20237 : _20238;
  always @ (posedge reset or posedge clock) if (reset) r1166 <= 1'd0; else if (_12300) r1166 <= _20239;
  wire [1:0] _20240 = {_0, _1854} + {_0, _3549};
  wire [1:0] _20241 = {_0, _4671} + {_0, _7036};
  wire [2:0] _20242 = {_0, _20240} + {_0, _20241};
  wire [1:0] _20243 = {_0, _9534} + {_0, _10941};
  wire [3:0] _20244 = {_0, _20242} + {_0, _0, _20243};
  wire _20245 = _12301 < _20244;
  wire _20246 = r1165 ^ _20245;
  wire _20247 = _12298 ? coded_block[1165] : r1165;
  wire _20248 = _12296 ? _20246 : _20247;
  always @ (posedge reset or posedge clock) if (reset) r1165 <= 1'd0; else if (_12300) r1165 <= _20248;
  wire [1:0] _20249 = {_0, _1886} + {_0, _3037};
  wire [1:0] _20250 = {_0, _5628} + {_0, _6750};
  wire [2:0] _20251 = {_0, _20249} + {_0, _20250};
  wire [1:0] _20252 = {_0, _9118} + {_0, _11613};
  wire [3:0] _20253 = {_0, _20251} + {_0, _0, _20252};
  wire _20254 = _12301 < _20253;
  wire _20255 = r1164 ^ _20254;
  wire _20256 = _12298 ? coded_block[1164] : r1164;
  wire _20257 = _12296 ? _20255 : _20256;
  always @ (posedge reset or posedge clock) if (reset) r1164 <= 1'd0; else if (_12300) r1164 <= _20257;
  wire [1:0] _20258 = {_0, _1215} + {_0, _3231};
  wire [1:0] _20259 = {_0, _5342} + {_0, _8186};
  wire [2:0] _20260 = {_0, _20258} + {_0, _20259};
  wire [1:0] _20261 = {_0, _8926} + {_0, _10877};
  wire [3:0] _20262 = {_0, _20260} + {_0, _0, _20261};
  wire _20263 = _12301 < _20262;
  wire _20264 = r1163 ^ _20263;
  wire _20265 = _12298 ? coded_block[1163] : r1163;
  wire _20266 = _12296 ? _20264 : _20265;
  always @ (posedge reset or posedge clock) if (reset) r1163 <= 1'd0; else if (_12300) r1163 <= _20266;
  wire [1:0] _20267 = {_0, _1247} + {_0, _4060};
  wire [1:0] _20268 = {_0, _5310} + {_0, _7420};
  wire [2:0] _20269 = {_0, _20267} + {_0, _20268};
  wire [1:0] _20270 = {_0, _8256} + {_0, _11004};
  wire [3:0] _20271 = {_0, _20269} + {_0, _0, _20270};
  wire _20272 = _12301 < _20271;
  wire _20273 = r1162 ^ _20272;
  wire _20274 = _12298 ? coded_block[1162] : r1162;
  wire _20275 = _12296 ? _20273 : _20274;
  always @ (posedge reset or posedge clock) if (reset) r1162 <= 1'd0; else if (_12300) r1162 <= _20275;
  wire [1:0] _20276 = {_0, _1278} + {_0, _2336};
  wire [1:0] _20277 = {_0, _6139} + {_0, _7389};
  wire [2:0] _20278 = {_0, _20276} + {_0, _20277};
  wire [1:0] _20279 = {_0, _9503} + {_0, _10335};
  wire [3:0] _20280 = {_0, _20278} + {_0, _0, _20279};
  wire _20281 = _12301 < _20280;
  wire _20282 = r1161 ^ _20281;
  wire _20283 = _12298 ? coded_block[1161] : r1161;
  wire _20284 = _12296 ? _20282 : _20283;
  always @ (posedge reset or posedge clock) if (reset) r1161 <= 1'd0; else if (_12300) r1161 <= _20284;
  wire [1:0] _20285 = {_0, _1312} + {_0, _3742};
  wire [1:0] _20286 = {_0, _4415} + {_0, _6207};
  wire [2:0] _20287 = {_0, _20285} + {_0, _20286};
  wire [1:0] _20288 = {_0, _9469} + {_0, _11581};
  wire [3:0] _20289 = {_0, _20287} + {_0, _0, _20288};
  wire _20290 = _12301 < _20289;
  wire _20291 = r1160 ^ _20290;
  wire _20292 = _12298 ? coded_block[1160] : r1160;
  wire _20293 = _12296 ? _20291 : _20292;
  always @ (posedge reset or posedge clock) if (reset) r1160 <= 1'd0; else if (_12300) r1160 <= _20293;
  wire [1:0] _20294 = {_0, _1343} + {_0, _3580};
  wire [1:0] _20295 = {_0, _5821} + {_0, _6494};
  wire [2:0] _20296 = {_0, _20294} + {_0, _20295};
  wire [1:0] _20297 = {_0, _8288} + {_0, _11550};
  wire [3:0] _20298 = {_0, _20296} + {_0, _0, _20297};
  wire _20299 = _12301 < _20298;
  wire _20300 = r1159 ^ _20299;
  wire _20301 = _12298 ? coded_block[1159] : r1159;
  wire _20302 = _12296 ? _20300 : _20301;
  always @ (posedge reset or posedge clock) if (reset) r1159 <= 1'd0; else if (_12300) r1159 <= _20302;
  wire [1:0] _20303 = {_0, _1375} + {_0, _2081};
  wire [1:0] _20304 = {_0, _5663} + {_0, _7900};
  wire [2:0] _20305 = {_0, _20303} + {_0, _20304};
  wire [1:0] _20306 = {_0, _8574} + {_0, _10366};
  wire [3:0] _20307 = {_0, _20305} + {_0, _0, _20306};
  wire _20308 = _12301 < _20307;
  wire _20309 = r1158 ^ _20308;
  wire _20310 = _12298 ? coded_block[1158] : r1158;
  wire _20311 = _12296 ? _20309 : _20310;
  always @ (posedge reset or posedge clock) if (reset) r1158 <= 1'd0; else if (_12300) r1158 <= _20311;
  wire [1:0] _20312 = {_0, _1406} + {_0, _3615};
  wire [1:0] _20313 = {_0, _4129} + {_0, _7741};
  wire [2:0] _20314 = {_0, _20312} + {_0, _20313};
  wire [1:0] _20315 = {_0, _9980} + {_0, _10654};
  wire [3:0] _20316 = {_0, _20314} + {_0, _0, _20315};
  wire _20317 = _12301 < _20316;
  wire _20318 = r1157 ^ _20317;
  wire _20319 = _12298 ? coded_block[1157] : r1157;
  wire _20320 = _12296 ? _20318 : _20319;
  always @ (posedge reset or posedge clock) if (reset) r1157 <= 1'd0; else if (_12300) r1157 <= _20320;
  wire [1:0] _20321 = {_0, _1439} + {_0, _3805};
  wire [1:0] _20322 = {_0, _5694} + {_0, _6176};
  wire [2:0] _20323 = {_0, _20321} + {_0, _20322};
  wire [1:0] _20324 = {_0, _9822} + {_0, _12061};
  wire [3:0] _20325 = {_0, _20323} + {_0, _0, _20324};
  wire _20326 = _12301 < _20325;
  wire _20327 = r1156 ^ _20326;
  wire _20328 = _12298 ? coded_block[1156] : r1156;
  wire _20329 = _12296 ? _20327 : _20328;
  always @ (posedge reset or posedge clock) if (reset) r1156 <= 1'd0; else if (_12300) r1156 <= _20329;
  wire [1:0] _20330 = {_0, _1470} + {_0, _2430};
  wire [1:0] _20331 = {_0, _5884} + {_0, _7773};
  wire [2:0] _20332 = {_0, _20330} + {_0, _20331};
  wire [1:0] _20333 = {_0, _8225} + {_0, _11900};
  wire [3:0] _20334 = {_0, _20332} + {_0, _0, _20333};
  wire _20335 = _12301 < _20334;
  wire _20336 = r1155 ^ _20335;
  wire _20337 = _12298 ? coded_block[1155] : r1155;
  wire _20338 = _12296 ? _20336 : _20337;
  always @ (posedge reset or posedge clock) if (reset) r1155 <= 1'd0; else if (_12300) r1155 <= _20338;
  wire [1:0] _20339 = {_0, _1502} + {_0, _2175};
  wire [1:0] _20340 = {_0, _4511} + {_0, _7965};
  wire [2:0] _20341 = {_0, _20339} + {_0, _20340};
  wire [1:0] _20342 = {_0, _9853} + {_0, _10272};
  wire [3:0] _20343 = {_0, _20341} + {_0, _0, _20342};
  wire _20344 = _12301 < _20343;
  wire _20345 = r1154 ^ _20344;
  wire _20346 = _12298 ? coded_block[1154] : r1154;
  wire _20347 = _12296 ? _20345 : _20346;
  always @ (posedge reset or posedge clock) if (reset) r1154 <= 1'd0; else if (_12300) r1154 <= _20347;
  wire [1:0] _20348 = {_0, _1568} + {_0, _3453};
  wire [1:0] _20349 = {_0, _5470} + {_0, _6334};
  wire [2:0] _20350 = {_0, _20348} + {_0, _20349};
  wire [1:0] _20351 = {_0, _8670} + {_0, _12124};
  wire [3:0] _20352 = {_0, _20350} + {_0, _0, _20351};
  wire _20353 = _12301 < _20352;
  wire _20354 = r1153 ^ _20353;
  wire _20355 = _12298 ? coded_block[1153] : r1153;
  wire _20356 = _12296 ? _20354 : _20355;
  always @ (posedge reset or posedge clock) if (reset) r1153 <= 1'd0; else if (_12300) r1153 <= _20356;
  wire [1:0] _20357 = {_0, _1599} + {_0, _2239};
  wire [1:0] _20358 = {_0, _5534} + {_0, _7548};
  wire [2:0] _20359 = {_0, _20357} + {_0, _20358};
  wire [1:0] _20360 = {_0, _8415} + {_0, _10748};
  wire [3:0] _20361 = {_0, _20359} + {_0, _0, _20360};
  wire _20362 = _12301 < _20361;
  wire _20363 = r1152 ^ _20362;
  wire _20364 = _12298 ? coded_block[1152] : r1152;
  wire _20365 = _12296 ? _20363 : _20364;
  always @ (posedge reset or posedge clock) if (reset) r1152 <= 1'd0; else if (_12300) r1152 <= _20365;
  wire [1:0] _20366 = {_0, _1631} + {_0, _2941};
  wire [1:0] _20367 = {_0, _4319} + {_0, _7612};
  wire [2:0] _20368 = {_0, _20366} + {_0, _20367};
  wire [1:0] _20369 = {_0, _9630} + {_0, _10493};
  wire [3:0] _20370 = {_0, _20368} + {_0, _0, _20369};
  wire _20371 = _12301 < _20370;
  wire _20372 = r1151 ^ _20371;
  wire _20373 = _12298 ? coded_block[1151] : r1151;
  wire _20374 = _12296 ? _20372 : _20373;
  always @ (posedge reset or posedge clock) if (reset) r1151 <= 1'd0; else if (_12300) r1151 <= _20374;
  wire [1:0] _20375 = {_0, _1662} + {_0, _2847};
  wire [1:0] _20376 = {_0, _5022} + {_0, _6397};
  wire [2:0] _20377 = {_0, _20375} + {_0, _20376};
  wire [1:0] _20378 = {_0, _9693} + {_0, _11708};
  wire [3:0] _20379 = {_0, _20377} + {_0, _0, _20378};
  wire _20380 = _12301 < _20379;
  wire _20381 = r1150 ^ _20380;
  wire _20382 = _12298 ? coded_block[1150] : r1150;
  wire _20383 = _12296 ? _20381 : _20382;
  always @ (posedge reset or posedge clock) if (reset) r1150 <= 1'd0; else if (_12300) r1150 <= _20383;
  wire [1:0] _20384 = {_0, _1695} + {_0, _3359};
  wire [1:0] _20385 = {_0, _4926} + {_0, _7100};
  wire [2:0] _20386 = {_0, _20384} + {_0, _20385};
  wire [1:0] _20387 = {_0, _8480} + {_0, _11771};
  wire [3:0] _20388 = {_0, _20386} + {_0, _0, _20387};
  wire _20389 = _12301 < _20388;
  wire _20390 = r1149 ^ _20389;
  wire _20391 = _12298 ? coded_block[1149] : r1149;
  wire _20392 = _12296 ? _20390 : _20391;
  always @ (posedge reset or posedge clock) if (reset) r1149 <= 1'd0; else if (_12300) r1149 <= _20392;
  wire [1:0] _20393 = {_0, _1726} + {_0, _2208};
  wire [1:0] _20394 = {_0, _5438} + {_0, _7005};
  wire [2:0] _20395 = {_0, _20393} + {_0, _20394};
  wire [1:0] _20396 = {_0, _9181} + {_0, _10558};
  wire [3:0] _20397 = {_0, _20395} + {_0, _0, _20396};
  wire _20398 = _12301 < _20397;
  wire _20399 = r1148 ^ _20398;
  wire _20400 = _12298 ? coded_block[1148] : r1148;
  wire _20401 = _12296 ? _20399 : _20400;
  always @ (posedge reset or posedge clock) if (reset) r1148 <= 1'd0; else if (_12300) r1148 <= _20401;
  wire [1:0] _20402 = {_0, _1758} + {_0, _3486};
  wire [1:0] _20403 = {_0, _4287} + {_0, _7517};
  wire [2:0] _20404 = {_0, _20402} + {_0, _20403};
  wire [1:0] _20405 = {_0, _9085} + {_0, _11259};
  wire [3:0] _20406 = {_0, _20404} + {_0, _0, _20405};
  wire _20407 = _12301 < _20406;
  wire _20408 = r1147 ^ _20407;
  wire _20409 = _12298 ? coded_block[1147] : r1147;
  wire _20410 = _12296 ? _20408 : _20409;
  always @ (posedge reset or posedge clock) if (reset) r1147 <= 1'd0; else if (_12300) r1147 <= _20410;
  wire [1:0] _20411 = {_0, _1789} + {_0, _2526};
  wire [1:0] _20412 = {_0, _5565} + {_0, _6366};
  wire [2:0] _20413 = {_0, _20411} + {_0, _20412};
  wire [1:0] _20414 = {_0, _9597} + {_0, _11165};
  wire [3:0] _20415 = {_0, _20413} + {_0, _0, _20414};
  wire _20416 = _12301 < _20415;
  wire _20417 = r1146 ^ _20416;
  wire _20418 = _12298 ? coded_block[1146] : r1146;
  wire _20419 = _12296 ? _20417 : _20418;
  always @ (posedge reset or posedge clock) if (reset) r1146 <= 1'd0; else if (_12300) r1146 <= _20419;
  wire [1:0] _20420 = {_0, _1823} + {_0, _3068};
  wire [1:0] _20421 = {_0, _4605} + {_0, _7644};
  wire [2:0] _20422 = {_0, _20420} + {_0, _20421};
  wire [1:0] _20423 = {_0, _8446} + {_0, _11677};
  wire [3:0] _20424 = {_0, _20422} + {_0, _0, _20423};
  wire _20425 = _12301 < _20424;
  wire _20426 = r1145 ^ _20425;
  wire _20427 = _12298 ? coded_block[1145] : r1145;
  wire _20428 = _12296 ? _20426 : _20427;
  always @ (posedge reset or posedge clock) if (reset) r1145 <= 1'd0; else if (_12300) r1145 <= _20428;
  wire [1:0] _20429 = {_0, _1854} + {_0, _2144};
  wire [1:0] _20430 = {_0, _5152} + {_0, _6687};
  wire [2:0] _20431 = {_0, _20429} + {_0, _20430};
  wire [1:0] _20432 = {_0, _9724} + {_0, _10527};
  wire [3:0] _20433 = {_0, _20431} + {_0, _0, _20432};
  wire _20434 = _12301 < _20433;
  wire _20435 = r1144 ^ _20434;
  wire _20436 = _12298 ? coded_block[1144] : r1144;
  wire _20437 = _12296 ? _20435 : _20436;
  always @ (posedge reset or posedge clock) if (reset) r1144 <= 1'd0; else if (_12300) r1144 <= _20437;
  wire [1:0] _20438 = {_0, _1886} + {_0, _2463};
  wire [1:0] _20439 = {_0, _4223} + {_0, _7230};
  wire [2:0] _20440 = {_0, _20438} + {_0, _20439};
  wire [1:0] _20441 = {_0, _8767} + {_0, _11806};
  wire [3:0] _20442 = {_0, _20440} + {_0, _0, _20441};
  wire _20443 = _12301 < _20442;
  wire _20444 = r1143 ^ _20443;
  wire _20445 = _12298 ? coded_block[1143] : r1143;
  wire _20446 = _12296 ? _20444 : _20445;
  always @ (posedge reset or posedge clock) if (reset) r1143 <= 1'd0; else if (_12300) r1143 <= _20446;
  wire [1:0] _20447 = {_0, _1917} + {_0, _2910};
  wire [1:0] _20448 = {_0, _4542} + {_0, _6303};
  wire [2:0] _20449 = {_0, _20447} + {_0, _20448};
  wire [1:0] _20450 = {_0, _9311} + {_0, _10846};
  wire [3:0] _20451 = {_0, _20449} + {_0, _0, _20450};
  wire _20452 = _12301 < _20451;
  wire _20453 = r1142 ^ _20452;
  wire _20454 = _12298 ? coded_block[1142] : r1142;
  wire _20455 = _12296 ? _20453 : _20454;
  always @ (posedge reset or posedge clock) if (reset) r1142 <= 1'd0; else if (_12300) r1142 <= _20455;
  wire [1:0] _20456 = {_0, _1950} + {_0, _2271};
  wire [1:0] _20457 = {_0, _4989} + {_0, _6621};
  wire [2:0] _20458 = {_0, _20456} + {_0, _20457};
  wire [1:0] _20459 = {_0, _8383} + {_0, _11389};
  wire [3:0] _20460 = {_0, _20458} + {_0, _0, _20459};
  wire _20461 = _12301 < _20460;
  wire _20462 = r1141 ^ _20461;
  wire _20463 = _12298 ? coded_block[1141] : r1141;
  wire _20464 = _12296 ? _20462 : _20463;
  always @ (posedge reset or posedge clock) if (reset) r1141 <= 1'd0; else if (_12300) r1141 <= _20464;
  wire [1:0] _20465 = {_0, _1981} + {_0, _3198};
  wire [1:0] _20466 = {_0, _4350} + {_0, _7069};
  wire [2:0] _20467 = {_0, _20465} + {_0, _20466};
  wire [1:0] _20468 = {_0, _8701} + {_0, _10462};
  wire [3:0] _20469 = {_0, _20467} + {_0, _0, _20468};
  wire _20470 = _12301 < _20469;
  wire _20471 = r1140 ^ _20470;
  wire _20472 = _12298 ? coded_block[1140] : r1140;
  wire _20473 = _12296 ? _20471 : _20472;
  always @ (posedge reset or posedge clock) if (reset) r1140 <= 1'd0; else if (_12300) r1140 <= _20473;
  wire [1:0] _20474 = {_0, _2013} + {_0, _3294};
  wire [1:0] _20475 = {_0, _5279} + {_0, _6431};
  wire [2:0] _20476 = {_0, _20474} + {_0, _20475};
  wire [1:0] _20477 = {_0, _9149} + {_0, _10783};
  wire [3:0] _20478 = {_0, _20476} + {_0, _0, _20477};
  wire _20479 = _12301 < _20478;
  wire _20480 = r1139 ^ _20479;
  wire _20481 = _12298 ? coded_block[1139] : r1139;
  wire _20482 = _12296 ? _20480 : _20481;
  always @ (posedge reset or posedge clock) if (reset) r1139 <= 1'd0; else if (_12300) r1139 <= _20482;
  wire [1:0] _20483 = {_0, _65} + {_0, _3005};
  wire [1:0] _20484 = {_0, _4830} + {_0, _7454};
  wire [2:0] _20485 = {_0, _20483} + {_0, _20484};
  wire [1:0] _20486 = {_0, _9438} + {_0, _10590};
  wire [3:0] _20487 = {_0, _20485} + {_0, _0, _20486};
  wire _20488 = _12301 < _20487;
  wire _20489 = r1138 ^ _20488;
  wire _20490 = _12298 ? coded_block[1138] : r1138;
  wire _20491 = _12296 ? _20489 : _20490;
  always @ (posedge reset or posedge clock) if (reset) r1138 <= 1'd0; else if (_12300) r1138 <= _20491;
  wire [1:0] _20492 = {_0, _97} + {_0, _3901};
  wire [1:0] _20493 = {_0, _5085} + {_0, _6908};
  wire [2:0] _20494 = {_0, _20492} + {_0, _20493};
  wire [1:0] _20495 = {_0, _9534} + {_0, _11516};
  wire [3:0] _20496 = {_0, _20494} + {_0, _0, _20495};
  wire _20497 = _12301 < _20496;
  wire _20498 = r1137 ^ _20497;
  wire _20499 = _12298 ? coded_block[1137] : r1137;
  wire _20500 = _12296 ? _20498 : _20499;
  always @ (posedge reset or posedge clock) if (reset) r1137 <= 1'd0; else if (_12300) r1137 <= _20500;
  wire [1:0] _20501 = {_0, _128} + {_0, _3549};
  wire [1:0] _20502 = {_0, _5981} + {_0, _7163};
  wire [2:0] _20503 = {_0, _20501} + {_0, _20502};
  wire [1:0] _20504 = {_0, _8991} + {_0, _11613};
  wire [3:0] _20505 = {_0, _20503} + {_0, _0, _20504};
  wire _20506 = _12301 < _20505;
  wire _20507 = r1136 ^ _20506;
  wire _20508 = _12298 ? coded_block[1136] : r1136;
  wire _20509 = _12296 ? _20507 : _20508;
  always @ (posedge reset or posedge clock) if (reset) r1136 <= 1'd0; else if (_12300) r1136 <= _20509;
  wire [1:0] _20510 = {_0, _161} + {_0, _3773};
  wire [1:0] _20511 = {_0, _5628} + {_0, _8059};
  wire [2:0] _20512 = {_0, _20510} + {_0, _20511};
  wire [1:0] _20513 = {_0, _9248} + {_0, _11069};
  wire [3:0] _20514 = {_0, _20512} + {_0, _0, _20513};
  wire _20515 = _12301 < _20514;
  wire _20516 = r1135 ^ _20515;
  wire _20517 = _12298 ? coded_block[1135] : r1135;
  wire _20518 = _12296 ? _20516 : _20517;
  always @ (posedge reset or posedge clock) if (reset) r1135 <= 1'd0; else if (_12300) r1135 <= _20518;
  wire [1:0] _20519 = {_0, _192} + {_0, _3646};
  wire [1:0] _20520 = {_0, _5853} + {_0, _7710};
  wire [2:0] _20521 = {_0, _20519} + {_0, _20520};
  wire [1:0] _20522 = {_0, _10141} + {_0, _11326};
  wire [3:0] _20523 = {_0, _20521} + {_0, _0, _20522};
  wire _20524 = _12301 < _20523;
  wire _20525 = r1134 ^ _20524;
  wire _20526 = _12298 ? coded_block[1134] : r1134;
  wire _20527 = _12296 ? _20525 : _20526;
  always @ (posedge reset or posedge clock) if (reset) r1134 <= 1'd0; else if (_12300) r1134 <= _20527;
  wire [1:0] _20528 = {_0, _224} + {_0, _3997};
  wire [1:0] _20529 = {_0, _5726} + {_0, _7931};
  wire [2:0] _20530 = {_0, _20528} + {_0, _20529};
  wire [1:0] _20531 = {_0, _9790} + {_0, _12219};
  wire [3:0] _20532 = {_0, _20530} + {_0, _0, _20531};
  wire _20533 = _12301 < _20532;
  wire _20534 = r1133 ^ _20533;
  wire _20535 = _12298 ? coded_block[1133] : r1133;
  wire _20536 = _12296 ? _20534 : _20535;
  always @ (posedge reset or posedge clock) if (reset) r1133 <= 1'd0; else if (_12300) r1133 <= _20536;
  wire [1:0] _20537 = {_0, _255} + {_0, _2719};
  wire [1:0] _20538 = {_0, _6076} + {_0, _7804};
  wire [2:0] _20539 = {_0, _20537} + {_0, _20538};
  wire [1:0] _20540 = {_0, _10014} + {_0, _11869};
  wire [3:0] _20541 = {_0, _20539} + {_0, _0, _20540};
  wire _20542 = _12301 < _20541;
  wire _20543 = r1132 ^ _20542;
  wire _20544 = _12298 ? coded_block[1132] : r1132;
  wire _20545 = _12296 ? _20543 : _20544;
  always @ (posedge reset or posedge clock) if (reset) r1132 <= 1'd0; else if (_12300) r1132 <= _20545;
  wire [1:0] _20546 = {_0, _289} + {_0, _3325};
  wire [1:0] _20547 = {_0, _4798} + {_0, _8155};
  wire [2:0] _20548 = {_0, _20546} + {_0, _20547};
  wire [1:0] _20549 = {_0, _9886} + {_0, _12092};
  wire [3:0] _20550 = {_0, _20548} + {_0, _0, _20549};
  wire _20551 = _12301 < _20550;
  wire _20552 = r1131 ^ _20551;
  wire _20553 = _12298 ? coded_block[1131] : r1131;
  wire _20554 = _12296 ? _20552 : _20553;
  always @ (posedge reset or posedge clock) if (reset) r1131 <= 1'd0; else if (_12300) r1131 <= _20554;
  wire [1:0] _20555 = {_0, _320} + {_0, _2878};
  wire [1:0] _20556 = {_0, _5407} + {_0, _6877};
  wire [2:0] _20557 = {_0, _20555} + {_0, _20556};
  wire [1:0] _20558 = {_0, _10235} + {_0, _11964};
  wire [3:0] _20559 = {_0, _20557} + {_0, _0, _20558};
  wire _20560 = _12301 < _20559;
  wire _20561 = r1130 ^ _20560;
  wire _20562 = _12298 ? coded_block[1130] : r1130;
  wire _20563 = _12296 ? _20561 : _20562;
  always @ (posedge reset or posedge clock) if (reset) r1130 <= 1'd0; else if (_12300) r1130 <= _20563;
  wire [1:0] _20564 = {_0, _383} + {_0, _3517};
  wire [1:0] _20565 = {_0, _4574} + {_0, _7036};
  wire [2:0] _20566 = {_0, _20564} + {_0, _20565};
  wire [1:0] _20567 = {_0, _9566} + {_0, _11038};
  wire [3:0] _20568 = {_0, _20566} + {_0, _0, _20567};
  wire _20569 = _12301 < _20568;
  wire _20570 = r1129 ^ _20569;
  wire _20571 = _12298 ? coded_block[1129] : r1129;
  wire _20572 = _12296 ? _20570 : _20571;
  always @ (posedge reset or posedge clock) if (reset) r1129 <= 1'd0; else if (_12300) r1129 <= _20572;
  wire [1:0] _20573 = {_0, _416} + {_0, _3933};
  wire [1:0] _20574 = {_0, _5597} + {_0, _6652};
  wire [2:0] _20575 = {_0, _20573} + {_0, _20574};
  wire [1:0] _20576 = {_0, _9118} + {_0, _11644};
  wire [3:0] _20577 = {_0, _20575} + {_0, _0, _20576};
  wire _20578 = _12301 < _20577;
  wire _20579 = r1128 ^ _20578;
  wire _20580 = _12298 ? coded_block[1128] : r1128;
  wire _20581 = _12296 ? _20579 : _20580;
  always @ (posedge reset or posedge clock) if (reset) r1128 <= 1'd0; else if (_12300) r1128 <= _20581;
  wire [1:0] _20582 = {_0, _447} + {_0, _2399};
  wire [1:0] _20583 = {_0, _6012} + {_0, _7675};
  wire [2:0] _20584 = {_0, _20582} + {_0, _20583};
  wire [1:0] _20585 = {_0, _8736} + {_0, _11196};
  wire [3:0] _20586 = {_0, _20584} + {_0, _0, _20585};
  wire _20587 = _12301 < _20586;
  wire _20588 = r1127 ^ _20587;
  wire _20589 = _12298 ? coded_block[1127] : r1127;
  wire _20590 = _12296 ? _20588 : _20589;
  always @ (posedge reset or posedge clock) if (reset) r1127 <= 1'd0; else if (_12300) r1127 <= _20590;
  wire [1:0] _20591 = {_0, _479} + {_0, _3836};
  wire [1:0] _20592 = {_0, _4478} + {_0, _8092};
  wire [2:0] _20593 = {_0, _20591} + {_0, _20592};
  wire [1:0] _20594 = {_0, _9759} + {_0, _10814};
  wire [3:0] _20595 = {_0, _20593} + {_0, _0, _20594};
  wire _20596 = _12301 < _20595;
  wire _20597 = r1126 ^ _20596;
  wire _20598 = _12298 ? coded_block[1126] : r1126;
  wire _20599 = _12296 ? _20597 : _20598;
  always @ (posedge reset or posedge clock) if (reset) r1126 <= 1'd0; else if (_12300) r1126 <= _20599;
  wire [1:0] _20600 = {_0, _510} + {_0, _3135};
  wire [1:0] _20601 = {_0, _5918} + {_0, _6558};
  wire [2:0] _20602 = {_0, _20600} + {_0, _20601};
  wire [1:0] _20603 = {_0, _10172} + {_0, _11837};
  wire [3:0] _20604 = {_0, _20602} + {_0, _0, _20603};
  wire _20605 = _12301 < _20604;
  wire _20606 = r1125 ^ _20605;
  wire _20607 = _12298 ? coded_block[1125] : r1125;
  wire _20608 = _12296 ? _20606 : _20607;
  always @ (posedge reset or posedge clock) if (reset) r1125 <= 1'd0; else if (_12300) r1125 <= _20608;
  wire [1:0] _20609 = {_0, _545} + {_0, _2813};
  wire [1:0] _20610 = {_0, _5215} + {_0, _7996};
  wire [2:0] _20611 = {_0, _20609} + {_0, _20610};
  wire [1:0] _20612 = {_0, _8638} + {_0, _12251};
  wire [3:0] _20613 = {_0, _20611} + {_0, _0, _20612};
  wire _20614 = _12301 < _20613;
  wire _20615 = r1124 ^ _20614;
  wire _20616 = _12298 ? coded_block[1124] : r1124;
  wire _20617 = _12296 ? _20615 : _20616;
  always @ (posedge reset or posedge clock) if (reset) r1124 <= 1'd0; else if (_12300) r1124 <= _20617;
  wire [1:0] _20618 = {_0, _576} + {_0, _2974};
  wire [1:0] _20619 = {_0, _4895} + {_0, _7293};
  wire [2:0] _20620 = {_0, _20618} + {_0, _20619};
  wire [1:0] _20621 = {_0, _10077} + {_0, _10717};
  wire [3:0] _20622 = {_0, _20620} + {_0, _0, _20621};
  wire _20623 = _12301 < _20622;
  wire _20624 = r1123 ^ _20623;
  wire _20625 = _12298 ? coded_block[1123] : r1123;
  wire _20626 = _12296 ? _20624 : _20625;
  always @ (posedge reset or posedge clock) if (reset) r1123 <= 1'd0; else if (_12300) r1123 <= _20626;
  wire [1:0] _20627 = {_0, _608} + {_0, _2782};
  wire [1:0] _20628 = {_0, _5053} + {_0, _6973};
  wire [2:0] _20629 = {_0, _20627} + {_0, _20628};
  wire [1:0] _20630 = {_0, _9375} + {_0, _12155};
  wire [3:0] _20631 = {_0, _20629} + {_0, _0, _20630};
  wire _20632 = _12301 < _20631;
  wire _20633 = r1122 ^ _20632;
  wire _20634 = _12298 ? coded_block[1122] : r1122;
  wire _20635 = _12296 ? _20633 : _20634;
  always @ (posedge reset or posedge clock) if (reset) r1122 <= 1'd0; else if (_12300) r1122 <= _20635;
  wire [1:0] _20636 = {_0, _672} + {_0, _2302};
  wire [1:0] _20637 = {_0, _5246} + {_0, _6942};
  wire [2:0] _20638 = {_0, _20636} + {_0, _20637};
  wire [1:0] _20639 = {_0, _9212} + {_0, _11132};
  wire [3:0] _20640 = {_0, _20638} + {_0, _0, _20639};
  wire _20641 = _12301 < _20640;
  wire _20642 = r1121 ^ _20641;
  wire _20643 = _12298 ? coded_block[1121] : r1121;
  wire _20644 = _12296 ? _20642 : _20643;
  always @ (posedge reset or posedge clock) if (reset) r1121 <= 1'd0; else if (_12300) r1121 <= _20644;
  wire [1:0] _20645 = {_0, _703} + {_0, _4091};
  wire [1:0] _20646 = {_0, _4384} + {_0, _7326};
  wire [2:0] _20647 = {_0, _20645} + {_0, _20646};
  wire [1:0] _20648 = {_0, _9022} + {_0, _11295};
  wire [3:0] _20649 = {_0, _20647} + {_0, _0, _20648};
  wire _20650 = _12301 < _20649;
  wire _20651 = r1120 ^ _20650;
  wire _20652 = _12298 ? coded_block[1120] : r1120;
  wire _20653 = _12296 ? _20651 : _20652;
  always @ (posedge reset or posedge clock) if (reset) r1120 <= 1'd0; else if (_12300) r1120 <= _20653;
  wire [1:0] _20654 = {_0, _735} + {_0, _2655};
  wire [1:0] _20655 = {_0, _4160} + {_0, _6462};
  wire [2:0] _20656 = {_0, _20654} + {_0, _20655};
  wire [1:0] _20657 = {_0, _9406} + {_0, _11101};
  wire [3:0] _20658 = {_0, _20656} + {_0, _0, _20657};
  wire _20659 = _12301 < _20658;
  wire _20660 = r1119 ^ _20659;
  wire _20661 = _12298 ? coded_block[1119] : r1119;
  wire _20662 = _12296 ? _20660 : _20661;
  always @ (posedge reset or posedge clock) if (reset) r1119 <= 1'd0; else if (_12300) r1119 <= _20662;
  wire [1:0] _20663 = {_0, _766} + {_0, _2592};
  wire [1:0] _20664 = {_0, _4734} + {_0, _6239};
  wire [2:0] _20665 = {_0, _20663} + {_0, _20664};
  wire [1:0] _20666 = {_0, _8543} + {_0, _11485};
  wire [3:0] _20667 = {_0, _20665} + {_0, _0, _20666};
  wire _20668 = _12301 < _20667;
  wire _20669 = r1118 ^ _20668;
  wire _20670 = _12298 ? coded_block[1118] : r1118;
  wire _20671 = _12296 ? _20669 : _20670;
  always @ (posedge reset or posedge clock) if (reset) r1118 <= 1'd0; else if (_12300) r1118 <= _20671;
  wire [1:0] _20672 = {_0, _800} + {_0, _3709};
  wire [1:0] _20673 = {_0, _4671} + {_0, _6814};
  wire [2:0] _20674 = {_0, _20672} + {_0, _20673};
  wire [1:0] _20675 = {_0, _8319} + {_0, _10621};
  wire [3:0] _20676 = {_0, _20674} + {_0, _0, _20675};
  wire _20677 = _12301 < _20676;
  wire _20678 = r1117 ^ _20677;
  wire _20679 = _12298 ? coded_block[1117] : r1117;
  wire _20680 = _12296 ? _20678 : _20679;
  always @ (posedge reset or posedge clock) if (reset) r1117 <= 1'd0; else if (_12300) r1117 <= _20680;
  wire [1:0] _20681 = {_0, _831} + {_0, _2367};
  wire [1:0] _20682 = {_0, _5790} + {_0, _6750};
  wire [2:0] _20683 = {_0, _20681} + {_0, _20682};
  wire [1:0] _20684 = {_0, _8894} + {_0, _10399};
  wire [3:0] _20685 = {_0, _20683} + {_0, _0, _20684};
  wire _20686 = _12301 < _20685;
  wire _20687 = r1116 ^ _20686;
  wire _20688 = _12298 ? coded_block[1116] : r1116;
  wire _20689 = _12296 ? _20687 : _20688;
  always @ (posedge reset or posedge clock) if (reset) r1116 <= 1'd0; else if (_12300) r1116 <= _20689;
  wire [1:0] _20690 = {_0, _863} + {_0, _3964};
  wire [1:0] _20691 = {_0, _4447} + {_0, _7868};
  wire [2:0] _20692 = {_0, _20690} + {_0, _20691};
  wire [1:0] _20693 = {_0, _8830} + {_0, _10973};
  wire [3:0] _20694 = {_0, _20692} + {_0, _0, _20693};
  wire _20695 = _12301 < _20694;
  wire _20696 = r1115 ^ _20695;
  wire _20697 = _12298 ? coded_block[1115] : r1115;
  wire _20698 = _12296 ? _20696 : _20697;
  always @ (posedge reset or posedge clock) if (reset) r1115 <= 1'd0; else if (_12300) r1115 <= _20698;
  wire [1:0] _20699 = {_0, _927} + {_0, _2623};
  wire [1:0] _20700 = {_0, _5757} + {_0, _8123};
  wire [2:0] _20701 = {_0, _20699} + {_0, _20700};
  wire [1:0] _20702 = {_0, _8607} + {_0, _12027};
  wire [3:0] _20703 = {_0, _20701} + {_0, _0, _20702};
  wire _20704 = _12301 < _20703;
  wire _20705 = r1114 ^ _20704;
  wire _20706 = _12298 ? coded_block[1114] : r1114;
  wire _20707 = _12296 ? _20705 : _20706;
  always @ (posedge reset or posedge clock) if (reset) r1114 <= 1'd0; else if (_12300) r1114 <= _20707;
  wire [1:0] _20708 = {_0, _1917} + {_0, _4028};
  wire [1:0] _20709 = {_0, _5116} + {_0, _7710};
  wire [2:0] _20710 = {_0, _20708} + {_0, _20709};
  wire [1:0] _20711 = {_0, _8830} + {_0, _11196};
  wire [3:0] _20712 = {_0, _20710} + {_0, _0, _20711};
  wire _20713 = _12301 < _20712;
  wire _20714 = r1113 ^ _20713;
  wire _20715 = _12298 ? coded_block[1113] : r1113;
  wire _20716 = _12296 ? _20714 : _20715;
  always @ (posedge reset or posedge clock) if (reset) r1113 <= 1'd0; else if (_12300) r1113 <= _20716;
  wire [1:0] _20717 = {_0, _1950} + {_0, _2782};
  wire [1:0] _20718 = {_0, _6108} + {_0, _7199};
  wire [2:0] _20719 = {_0, _20717} + {_0, _20718};
  wire [1:0] _20720 = {_0, _9790} + {_0, _10910};
  wire [3:0] _20721 = {_0, _20719} + {_0, _0, _20720};
  wire _20722 = _12301 < _20721;
  wire _20723 = r1112 ^ _20722;
  wire _20724 = _12298 ? coded_block[1112] : r1112;
  wire _20725 = _12296 ? _20723 : _20724;
  always @ (posedge reset or posedge clock) if (reset) r1112 <= 1'd0; else if (_12300) r1112 <= _20725;
  wire [1:0] _20726 = {_0, _703} + {_0, _3709};
  wire [1:0] _20727 = {_0, _5342} + {_0, _7100};
  wire [2:0] _20728 = {_0, _20726} + {_0, _20727};
  wire [1:0] _20729 = {_0, _10108} + {_0, _11644};
  wire [3:0] _20730 = {_0, _20728} + {_0, _0, _20729};
  wire _20731 = _12301 < _20730;
  wire _20732 = r1111 ^ _20731;
  wire _20733 = _12298 ? coded_block[1111] : r1111;
  wire _20734 = _12296 ? _20732 : _20733;
  always @ (posedge reset or posedge clock) if (reset) r1111 <= 1'd0; else if (_12300) r1111 <= _20734;
  wire [1:0] _20735 = {_0, _1981} + {_0, _3964};
  wire [1:0] _20736 = {_0, _4861} + {_0, _8186};
  wire [2:0] _20737 = {_0, _20735} + {_0, _20736};
  wire [1:0] _20738 = {_0, _9279} + {_0, _11869};
  wire [3:0] _20739 = {_0, _20737} + {_0, _0, _20738};
  wire _20740 = _12301 < _20739;
  wire _20741 = r1110 ^ _20740;
  wire _20742 = _12298 ? coded_block[1110] : r1110;
  wire _20743 = _12296 ? _20741 : _20742;
  always @ (posedge reset or posedge clock) if (reset) r1110 <= 1'd0; else if (_12300) r1110 <= _20743;
  wire [1:0] _20744 = {_0, _766} + {_0, _3997};
  wire [1:0] _20745 = {_0, _5152} + {_0, _7868};
  wire [2:0] _20746 = {_0, _20744} + {_0, _20745};
  wire [1:0] _20747 = {_0, _9503} + {_0, _11259};
  wire [3:0] _20748 = {_0, _20746} + {_0, _0, _20747};
  wire _20749 = _12301 < _20748;
  wire _20750 = r1109 ^ _20749;
  wire _20751 = _12298 ? coded_block[1109] : r1109;
  wire _20752 = _12296 ? _20750 : _20751;
  always @ (posedge reset or posedge clock) if (reset) r1109 <= 1'd0; else if (_12300) r1109 <= _20752;
  wire [1:0] _20753 = {_0, _2013} + {_0, _3486};
  wire [1:0] _20754 = {_0, _6045} + {_0, _6942};
  wire [2:0] _20755 = {_0, _20753} + {_0, _20754};
  wire [1:0] _20756 = {_0, _8256} + {_0, _11358};
  wire [3:0] _20757 = {_0, _20755} + {_0, _0, _20756};
  wire _20758 = _12301 < _20757;
  wire _20759 = r1108 ^ _20758;
  wire _20760 = _12298 ? coded_block[1108] : r1108;
  wire _20761 = _12296 ? _20759 : _20760;
  always @ (posedge reset or posedge clock) if (reset) r1108 <= 1'd0; else if (_12300) r1108 <= _20761;
  wire [1:0] _20762 = {_0, _831} + {_0, _3549};
  wire [1:0] _20763 = {_0, _4160} + {_0, _8155};
  wire [2:0] _20764 = {_0, _20762} + {_0, _20763};
  wire [1:0] _20765 = {_0, _9311} + {_0, _12027};
  wire [3:0] _20766 = {_0, _20764} + {_0, _0, _20765};
  wire _20767 = _12301 < _20766;
  wire _20768 = r1107 ^ _20767;
  wire _20769 = _12298 ? coded_block[1107] : r1107;
  wire _20770 = _12296 ? _20768 : _20769;
  always @ (posedge reset or posedge clock) if (reset) r1107 <= 1'd0; else if (_12300) r1107 <= _20770;
  wire [1:0] _20771 = {_0, _863} + {_0, _3805};
  wire [1:0] _20772 = {_0, _5628} + {_0, _6239};
  wire [2:0] _20773 = {_0, _20771} + {_0, _20772};
  wire [1:0] _20774 = {_0, _10235} + {_0, _11389};
  wire [3:0] _20775 = {_0, _20773} + {_0, _0, _20774};
  wire _20776 = _12301 < _20775;
  wire _20777 = r1106 ^ _20776;
  wire _20778 = _12298 ? coded_block[1106] : r1106;
  wire _20779 = _12296 ? _20777 : _20778;
  always @ (posedge reset or posedge clock) if (reset) r1106 <= 1'd0; else if (_12300) r1106 <= _20779;
  wire [1:0] _20780 = {_0, _894} + {_0, _2686};
  wire [1:0] _20781 = {_0, _5884} + {_0, _7710};
  wire [2:0] _20782 = {_0, _20780} + {_0, _20781};
  wire [1:0] _20783 = {_0, _8319} + {_0, _10303};
  wire [3:0] _20784 = {_0, _20782} + {_0, _0, _20783};
  wire _20785 = _12301 < _20784;
  wire _20786 = r1105 ^ _20785;
  wire _20787 = _12298 ? coded_block[1105] : r1105;
  wire _20788 = _12296 ? _20786 : _20787;
  always @ (posedge reset or posedge clock) if (reset) r1105 <= 1'd0; else if (_12300) r1105 <= _20788;
  wire [1:0] _20789 = {_0, _927} + {_0, _2336};
  wire [1:0] _20790 = {_0, _4767} + {_0, _7965};
  wire [2:0] _20791 = {_0, _20789} + {_0, _20790};
  wire [1:0] _20792 = {_0, _9790} + {_0, _10399};
  wire [3:0] _20793 = {_0, _20791} + {_0, _0, _20792};
  wire _20794 = _12301 < _20793;
  wire _20795 = r1104 ^ _20794;
  wire _20796 = _12298 ? coded_block[1104] : r1104;
  wire _20797 = _12296 ? _20795 : _20796;
  always @ (posedge reset or posedge clock) if (reset) r1104 <= 1'd0; else if (_12300) r1104 <= _20797;
  wire [1:0] _20798 = {_0, _958} + {_0, _2557};
  wire [1:0] _20799 = {_0, _4415} + {_0, _6845};
  wire [2:0] _20800 = {_0, _20798} + {_0, _20799};
  wire [1:0] _20801 = {_0, _10045} + {_0, _11869};
  wire [3:0] _20802 = {_0, _20800} + {_0, _0, _20801};
  wire _20803 = _12301 < _20802;
  wire _20804 = r1103 ^ _20803;
  wire _20805 = _12298 ? coded_block[1103] : r1103;
  wire _20806 = _12296 ? _20804 : _20805;
  always @ (posedge reset or posedge clock) if (reset) r1103 <= 1'd0; else if (_12300) r1103 <= _20806;
  wire [1:0] _20807 = {_0, _990} + {_0, _2430};
  wire [1:0] _20808 = {_0, _4640} + {_0, _6494};
  wire [2:0] _20809 = {_0, _20807} + {_0, _20808};
  wire [1:0] _20810 = {_0, _8926} + {_0, _12124};
  wire [3:0] _20811 = {_0, _20809} + {_0, _0, _20810};
  wire _20812 = _12301 < _20811;
  wire _20813 = r1102 ^ _20812;
  wire _20814 = _12298 ? coded_block[1102] : r1102;
  wire _20815 = _12296 ? _20813 : _20814;
  always @ (posedge reset or posedge clock) if (reset) r1102 <= 1'd0; else if (_12300) r1102 <= _20815;
  wire [1:0] _20816 = {_0, _1021} + {_0, _2782};
  wire [1:0] _20817 = {_0, _4511} + {_0, _6718};
  wire [2:0] _20818 = {_0, _20816} + {_0, _20817};
  wire [1:0] _20819 = {_0, _8574} + {_0, _11004};
  wire [3:0] _20820 = {_0, _20818} + {_0, _0, _20819};
  wire _20821 = _12301 < _20820;
  wire _20822 = r1101 ^ _20821;
  wire _20823 = _12298 ? coded_block[1101] : r1101;
  wire _20824 = _12296 ? _20822 : _20823;
  always @ (posedge reset or posedge clock) if (reset) r1101 <= 1'd0; else if (_12300) r1101 <= _20824;
  wire [1:0] _20825 = {_0, _1088} + {_0, _2112};
  wire [1:0] _20826 = {_0, _5597} + {_0, _6942};
  wire [2:0] _20827 = {_0, _20825} + {_0, _20826};
  wire [1:0] _20828 = {_0, _8670} + {_0, _10877};
  wire [3:0] _20829 = {_0, _20827} + {_0, _0, _20828};
  wire _20830 = _12301 < _20829;
  wire _20831 = r1100 ^ _20830;
  wire _20832 = _12298 ? coded_block[1100] : r1100;
  wire _20833 = _12296 ? _20831 : _20832;
  always @ (posedge reset or posedge clock) if (reset) r1100 <= 1'd0; else if (_12300) r1100 <= _20833;
  wire [1:0] _20834 = {_0, _1120} + {_0, _3678};
  wire [1:0] _20835 = {_0, _4192} + {_0, _7675};
  wire [2:0] _20836 = {_0, _20834} + {_0, _20835};
  wire [1:0] _20837 = {_0, _9022} + {_0, _10748};
  wire [3:0] _20838 = {_0, _20836} + {_0, _0, _20837};
  wire _20839 = _12301 < _20838;
  wire _20840 = r1099 ^ _20839;
  wire _20841 = _12298 ? coded_block[1099] : r1099;
  wire _20842 = _12296 ? _20840 : _20841;
  always @ (posedge reset or posedge clock) if (reset) r1099 <= 1'd0; else if (_12300) r1099 <= _20842;
  wire [1:0] _20843 = {_0, _1151} + {_0, _3294};
  wire [1:0] _20844 = {_0, _5757} + {_0, _6270};
  wire [2:0] _20845 = {_0, _20843} + {_0, _20844};
  wire [1:0] _20846 = {_0, _9759} + {_0, _11101};
  wire [3:0] _20847 = {_0, _20845} + {_0, _0, _20846};
  wire _20848 = _12301 < _20847;
  wire _20849 = r1098 ^ _20848;
  wire _20850 = _12298 ? coded_block[1098] : r1098;
  wire _20851 = _12296 ? _20849 : _20850;
  always @ (posedge reset or posedge clock) if (reset) r1098 <= 1'd0; else if (_12300) r1098 <= _20851;
  wire [1:0] _20852 = {_0, _1215} + {_0, _2719};
  wire [1:0] _20853 = {_0, _4384} + {_0, _7454};
  wire [2:0] _20854 = {_0, _20852} + {_0, _20853};
  wire [1:0] _20855 = {_0, _9917} + {_0, _10430};
  wire [3:0] _20856 = {_0, _20854} + {_0, _0, _20855};
  wire _20857 = _12301 < _20856;
  wire _20858 = r1097 ^ _20857;
  wire _20859 = _12298 ? coded_block[1097] : r1097;
  wire _20860 = _12296 ? _20858 : _20859;
  always @ (posedge reset or posedge clock) if (reset) r1097 <= 1'd0; else if (_12300) r1097 <= _20860;
  wire [1:0] _20861 = {_0, _1247} + {_0, _3198};
  wire [1:0] _20862 = {_0, _4798} + {_0, _6462};
  wire [2:0] _20863 = {_0, _20861} + {_0, _20862};
  wire [1:0] _20864 = {_0, _9534} + {_0, _11996};
  wire [3:0] _20865 = {_0, _20863} + {_0, _0, _20864};
  wire _20866 = _12301 < _20865;
  wire _20867 = r1096 ^ _20866;
  wire _20868 = _12298 ? coded_block[1096] : r1096;
  wire _20869 = _12296 ? _20867 : _20868;
  always @ (posedge reset or posedge clock) if (reset) r1096 <= 1'd0; else if (_12300) r1096 <= _20869;
  wire [1:0] _20870 = {_0, _1278} + {_0, _2623};
  wire [1:0] _20871 = {_0, _5279} + {_0, _6877};
  wire [2:0] _20872 = {_0, _20870} + {_0, _20871};
  wire [1:0] _20873 = {_0, _8543} + {_0, _11613};
  wire [3:0] _20874 = {_0, _20872} + {_0, _0, _20873};
  wire _20875 = _12301 < _20874;
  wire _20876 = r1095 ^ _20875;
  wire _20877 = _12298 ? coded_block[1095] : r1095;
  wire _20878 = _12296 ? _20876 : _20877;
  always @ (posedge reset or posedge clock) if (reset) r1095 <= 1'd0; else if (_12300) r1095 <= _20878;
  wire [1:0] _20879 = {_0, _1343} + {_0, _3615};
  wire [1:0] _20880 = {_0, _6012} + {_0, _6781};
  wire [2:0] _20881 = {_0, _20879} + {_0, _20880};
  wire [1:0] _20882 = {_0, _9438} + {_0, _11038};
  wire [3:0] _20883 = {_0, _20881} + {_0, _0, _20882};
  wire _20884 = _12301 < _20883;
  wire _20885 = r1094 ^ _20884;
  wire _20886 = _12298 ? coded_block[1094] : r1094;
  wire _20887 = _12296 ? _20885 : _20886;
  always @ (posedge reset or posedge clock) if (reset) r1094 <= 1'd0; else if (_12300) r1094 <= _20887;
  wire [1:0] _20888 = {_0, _1375} + {_0, _3773};
  wire [1:0] _20889 = {_0, _5694} + {_0, _8092};
  wire [2:0] _20890 = {_0, _20888} + {_0, _20889};
  wire [1:0] _20891 = {_0, _8863} + {_0, _11516};
  wire [3:0] _20892 = {_0, _20890} + {_0, _0, _20891};
  wire _20893 = _12301 < _20892;
  wire _20894 = r1093 ^ _20893;
  wire _20895 = _12298 ? coded_block[1093] : r1093;
  wire _20896 = _12296 ? _20894 : _20895;
  always @ (posedge reset or posedge clock) if (reset) r1093 <= 1'd0; else if (_12300) r1093 <= _20896;
  wire [1:0] _20897 = {_0, _1406} + {_0, _3580};
  wire [1:0] _20898 = {_0, _5853} + {_0, _7773};
  wire [2:0] _20899 = {_0, _20897} + {_0, _20898};
  wire [1:0] _20900 = {_0, _10172} + {_0, _10941};
  wire [3:0] _20901 = {_0, _20899} + {_0, _0, _20900};
  wire _20902 = _12301 < _20901;
  wire _20903 = r1092 ^ _20902;
  wire _20904 = _12298 ? coded_block[1092] : r1092;
  wire _20905 = _12296 ? _20903 : _20904;
  always @ (posedge reset or posedge clock) if (reset) r1092 <= 1'd0; else if (_12300) r1092 <= _20905;
  wire [1:0] _20906 = {_0, _1439} + {_0, _3964};
  wire [1:0] _20907 = {_0, _5663} + {_0, _7931};
  wire [2:0] _20908 = {_0, _20906} + {_0, _20907};
  wire [1:0] _20909 = {_0, _9853} + {_0, _12251};
  wire [3:0] _20910 = {_0, _20908} + {_0, _0, _20909};
  wire _20911 = _12301 < _20910;
  wire _20912 = r1091 ^ _20911;
  wire _20913 = _12298 ? coded_block[1091] : r1091;
  wire _20914 = _12296 ? _20912 : _20913;
  always @ (posedge reset or posedge clock) if (reset) r1091 <= 1'd0; else if (_12300) r1091 <= _20914;
  wire [1:0] _20915 = {_0, _1470} + {_0, _3104};
  wire [1:0] _20916 = {_0, _6045} + {_0, _7741};
  wire [2:0] _20917 = {_0, _20915} + {_0, _20916};
  wire [1:0] _20918 = {_0, _10014} + {_0, _11933};
  wire [3:0] _20919 = {_0, _20917} + {_0, _0, _20918};
  wire _20920 = _12301 < _20919;
  wire _20921 = r1090 ^ _20920;
  wire _20922 = _12298 ? coded_block[1090] : r1090;
  wire _20923 = _12296 ? _20921 : _20922;
  always @ (posedge reset or posedge clock) if (reset) r1090 <= 1'd0; else if (_12300) r1090 <= _20923;
  wire [1:0] _20924 = {_0, _1568} + {_0, _3390};
  wire [1:0] _20925 = {_0, _5534} + {_0, _7036};
  wire [2:0] _20926 = {_0, _20924} + {_0, _20925};
  wire [1:0] _20927 = {_0, _9342} + {_0, _12282};
  wire [3:0] _20928 = {_0, _20926} + {_0, _0, _20927};
  wire _20929 = _12301 < _20928;
  wire _20930 = r1089 ^ _20929;
  wire _20931 = _12298 ? coded_block[1089] : r1089;
  wire _20932 = _12296 ? _20930 : _20931;
  always @ (posedge reset or posedge clock) if (reset) r1089 <= 1'd0; else if (_12300) r1089 <= _20932;
  wire [1:0] _20933 = {_0, _1599} + {_0, _2494};
  wire [1:0] _20934 = {_0, _5470} + {_0, _7612};
  wire [2:0] _20935 = {_0, _20933} + {_0, _20934};
  wire [1:0] _20936 = {_0, _9118} + {_0, _11422};
  wire [3:0] _20937 = {_0, _20935} + {_0, _0, _20936};
  wire _20938 = _12301 < _20937;
  wire _20939 = r1088 ^ _20938;
  wire _20940 = _12298 ? coded_block[1088] : r1088;
  wire _20941 = _12296 ? _20939 : _20940;
  always @ (posedge reset or posedge clock) if (reset) r1088 <= 1'd0; else if (_12300) r1088 <= _20941;
  wire [1:0] _20942 = {_0, _1662} + {_0, _2750};
  wire [1:0] _20943 = {_0, _5246} + {_0, _6652};
  wire [2:0] _20944 = {_0, _20942} + {_0, _20943};
  wire [1:0] _20945 = {_0, _9630} + {_0, _11771};
  wire [3:0] _20946 = {_0, _20944} + {_0, _0, _20945};
  wire _20947 = _12301 < _20946;
  wire _20948 = r1087 ^ _20947;
  wire _20949 = _12298 ? coded_block[1087] : r1087;
  wire _20950 = _12296 ? _20948 : _20949;
  always @ (posedge reset or posedge clock) if (reset) r1087 <= 1'd0; else if (_12300) r1087 <= _20950;
  wire [1:0] _20951 = {_0, _1695} + {_0, _2463};
  wire [1:0] _20952 = {_0, _4830} + {_0, _7326};
  wire [2:0] _20953 = {_0, _20951} + {_0, _20952};
  wire [1:0] _20954 = {_0, _8736} + {_0, _11708};
  wire [3:0] _20955 = {_0, _20953} + {_0, _0, _20954};
  wire _20956 = _12301 < _20955;
  wire _20957 = r1086 ^ _20956;
  wire _20958 = _12298 ? coded_block[1086] : r1086;
  wire _20959 = _12296 ? _20957 : _20958;
  always @ (posedge reset or posedge clock) if (reset) r1086 <= 1'd0; else if (_12300) r1086 <= _20959;
  wire [1:0] _20960 = {_0, _1726} + {_0, _3422};
  wire [1:0] _20961 = {_0, _4542} + {_0, _6908};
  wire [2:0] _20962 = {_0, _20960} + {_0, _20961};
  wire [1:0] _20963 = {_0, _9406} + {_0, _10814};
  wire [3:0] _20964 = {_0, _20962} + {_0, _0, _20963};
  wire _20965 = _12301 < _20964;
  wire _20966 = r1085 ^ _20965;
  wire _20967 = _12298 ? coded_block[1085] : r1085;
  wire _20968 = _12296 ? _20966 : _20967;
  always @ (posedge reset or posedge clock) if (reset) r1085 <= 1'd0; else if (_12300) r1085 <= _20968;
  wire [1:0] _20969 = {_0, _1758} + {_0, _2910};
  wire [1:0] _20970 = {_0, _5501} + {_0, _6621};
  wire [2:0] _20971 = {_0, _20969} + {_0, _20970};
  wire [1:0] _20972 = {_0, _8991} + {_0, _11485};
  wire [3:0] _20973 = {_0, _20971} + {_0, _0, _20972};
  wire _20974 = _12301 < _20973;
  wire _20975 = r1084 ^ _20974;
  wire _20976 = _12298 ? coded_block[1084] : r1084;
  wire _20977 = _12296 ? _20975 : _20976;
  always @ (posedge reset or posedge clock) if (reset) r1084 <= 1'd0; else if (_12300) r1084 <= _20977;
  wire [1:0] _20978 = {_0, _1789} + {_0, _3901};
  wire [1:0] _20979 = {_0, _4989} + {_0, _7581};
  wire [2:0] _20980 = {_0, _20978} + {_0, _20979};
  wire [1:0] _20981 = {_0, _8701} + {_0, _11069};
  wire [3:0] _20982 = {_0, _20980} + {_0, _0, _20981};
  wire _20983 = _12301 < _20982;
  wire _20984 = r1083 ^ _20983;
  wire _20985 = _12298 ? coded_block[1083] : r1083;
  wire _20986 = _12296 ? _20984 : _20985;
  always @ (posedge reset or posedge clock) if (reset) r1083 <= 1'd0; else if (_12300) r1083 <= _20986;
  wire [1:0] _20987 = {_0, _1823} + {_0, _2655};
  wire [1:0] _20988 = {_0, _5981} + {_0, _7069};
  wire [2:0] _20989 = {_0, _20987} + {_0, _20988};
  wire [1:0] _20990 = {_0, _9661} + {_0, _10783};
  wire [3:0] _20991 = {_0, _20989} + {_0, _0, _20990};
  wire _20992 = _12301 < _20991;
  wire _20993 = r1082 ^ _20992;
  wire _20994 = _12298 ? coded_block[1082] : r1082;
  wire _20995 = _12296 ? _20993 : _20994;
  always @ (posedge reset or posedge clock) if (reset) r1082 <= 1'd0; else if (_12300) r1082 <= _20995;
  wire [1:0] _20996 = {_0, _1854} + {_0, _3836};
  wire [1:0] _20997 = {_0, _4734} + {_0, _8059};
  wire [2:0] _20998 = {_0, _20996} + {_0, _20997};
  wire [1:0] _20999 = {_0, _9149} + {_0, _11740};
  wire [3:0] _21000 = {_0, _20998} + {_0, _0, _20999};
  wire _21001 = _12301 < _21000;
  wire _21002 = r1081 ^ _21001;
  wire _21003 = _12298 ? coded_block[1081] : r1081;
  wire _21004 = _12296 ? _21002 : _21003;
  always @ (posedge reset or posedge clock) if (reset) r1081 <= 1'd0; else if (_12300) r1081 <= _21004;
  wire [1:0] _21005 = {_0, _1886} + {_0, _3359};
  wire [1:0] _21006 = {_0, _5918} + {_0, _6814};
  wire [2:0] _21007 = {_0, _21005} + {_0, _21006};
  wire [1:0] _21008 = {_0, _10141} + {_0, _11228};
  wire [3:0] _21009 = {_0, _21007} + {_0, _0, _21008};
  wire _21010 = _12301 < _21009;
  wire _21011 = r1080 ^ _21010;
  wire _21012 = _12298 ? coded_block[1080] : r1080;
  wire _21013 = _12296 ? _21011 : _21012;
  always @ (posedge reset or posedge clock) if (reset) r1080 <= 1'd0; else if (_12300) r1080 <= _21013;
  wire [1:0] _21014 = {_0, _1981} + {_0, _4060};
  wire [1:0] _21015 = {_0, _4895} + {_0, _7644};
  wire [2:0] _21016 = {_0, _21014} + {_0, _21015};
  wire [1:0] _21017 = {_0, _9597} + {_0, _12155};
  wire [3:0] _21018 = {_0, _21016} + {_0, _0, _21017};
  wire _21019 = _12301 < _21018;
  wire _21020 = r1079 ^ _21019;
  wire _21021 = _12298 ? coded_block[1079] : r1079;
  wire _21022 = _12296 ? _21020 : _21021;
  always @ (posedge reset or posedge clock) if (reset) r1079 <= 1'd0; else if (_12300) r1079 <= _21022;
  wire [1:0] _21023 = {_0, _2013} + {_0, _4028};
  wire [1:0] _21024 = {_0, _6139} + {_0, _6973};
  wire [2:0] _21025 = {_0, _21023} + {_0, _21024};
  wire [1:0] _21026 = {_0, _9724} + {_0, _11677};
  wire [3:0] _21027 = {_0, _21025} + {_0, _0, _21026};
  wire _21028 = _12301 < _21027;
  wire _21029 = r1078 ^ _21028;
  wire _21030 = _12298 ? coded_block[1078] : r1078;
  wire _21031 = _12296 ? _21029 : _21030;
  always @ (posedge reset or posedge clock) if (reset) r1078 <= 1'd0; else if (_12300) r1078 <= _21031;
  wire [1:0] _21032 = {_0, _65} + {_0, _3135};
  wire [1:0] _21033 = {_0, _4926} + {_0, _8186};
  wire [2:0] _21034 = {_0, _21032} + {_0, _21033};
  wire [1:0] _21035 = {_0, _8288} + {_0, _11132};
  wire [3:0] _21036 = {_0, _21034} + {_0, _0, _21035};
  wire _21037 = _12301 < _21036;
  wire _21038 = r1077 ^ _21037;
  wire _21039 = _12298 ? coded_block[1077] : r1077;
  wire _21040 = _12296 ? _21038 : _21039;
  always @ (posedge reset or posedge clock) if (reset) r1077 <= 1'd0; else if (_12300) r1077 <= _21040;
  wire [1:0] _21041 = {_0, _97} + {_0, _2526};
  wire [1:0] _21042 = {_0, _5215} + {_0, _7005};
  wire [2:0] _21043 = {_0, _21041} + {_0, _21042};
  wire [1:0] _21044 = {_0, _8256} + {_0, _10366};
  wire [3:0] _21045 = {_0, _21043} + {_0, _0, _21044};
  wire _21046 = _12301 < _21045;
  wire _21047 = r1076 ^ _21046;
  wire _21048 = _12298 ? coded_block[1076] : r1076;
  wire _21049 = _12296 ? _21047 : _21048;
  always @ (posedge reset or posedge clock) if (reset) r1076 <= 1'd0; else if (_12300) r1076 <= _21049;
  wire [1:0] _21050 = {_0, _128} + {_0, _2367};
  wire [1:0] _21051 = {_0, _4605} + {_0, _7293};
  wire [2:0] _21052 = {_0, _21050} + {_0, _21051};
  wire [1:0] _21053 = {_0, _9085} + {_0, _10335};
  wire [3:0] _21054 = {_0, _21052} + {_0, _0, _21053};
  wire _21055 = _12301 < _21054;
  wire _21056 = r1075 ^ _21055;
  wire _21057 = _12298 ? coded_block[1075] : r1075;
  wire _21058 = _12296 ? _21056 : _21057;
  always @ (posedge reset or posedge clock) if (reset) r1075 <= 1'd0; else if (_12300) r1075 <= _21058;
  wire [1:0] _21059 = {_0, _161} + {_0, _2081};
  wire [1:0] _21060 = {_0, _4447} + {_0, _6687};
  wire [2:0] _21061 = {_0, _21059} + {_0, _21060};
  wire [1:0] _21062 = {_0, _9375} + {_0, _11165};
  wire [3:0] _21063 = {_0, _21061} + {_0, _0, _21062};
  wire _21064 = _12301 < _21063;
  wire _21065 = r1074 ^ _21064;
  wire _21066 = _12298 ? coded_block[1074] : r1074;
  wire _21067 = _12296 ? _21065 : _21066;
  always @ (posedge reset or posedge clock) if (reset) r1074 <= 1'd0; else if (_12300) r1074 <= _21067;
  wire [1:0] _21068 = {_0, _192} + {_0, _2399};
  wire [1:0] _21069 = {_0, _4129} + {_0, _6525};
  wire [2:0] _21070 = {_0, _21068} + {_0, _21069};
  wire [1:0] _21071 = {_0, _8767} + {_0, _11453};
  wire [3:0] _21072 = {_0, _21070} + {_0, _0, _21071};
  wire _21073 = _12301 < _21072;
  wire _21074 = r1073 ^ _21073;
  wire _21075 = _12298 ? coded_block[1073] : r1073;
  wire _21076 = _12296 ? _21074 : _21075;
  always @ (posedge reset or posedge clock) if (reset) r1073 <= 1'd0; else if (_12300) r1073 <= _21076;
  wire [1:0] _21077 = {_0, _224} + {_0, _2592};
  wire [1:0] _21078 = {_0, _4478} + {_0, _6176};
  wire [2:0] _21079 = {_0, _21077} + {_0, _21078};
  wire [1:0] _21080 = {_0, _8607} + {_0, _10846};
  wire [3:0] _21081 = {_0, _21079} + {_0, _0, _21080};
  wire _21082 = _12301 < _21081;
  wire _21083 = r1072 ^ _21082;
  wire _21084 = _12298 ? coded_block[1072] : r1072;
  wire _21085 = _12296 ? _21083 : _21084;
  always @ (posedge reset or posedge clock) if (reset) r1072 <= 1'd0; else if (_12300) r1072 <= _21085;
  wire [1:0] _21086 = {_0, _255} + {_0, _3231};
  wire [1:0] _21087 = {_0, _4671} + {_0, _6558};
  wire [2:0] _21088 = {_0, _21086} + {_0, _21087};
  wire [1:0] _21089 = {_0, _8225} + {_0, _10685};
  wire [3:0] _21090 = {_0, _21088} + {_0, _0, _21089};
  wire _21091 = _12301 < _21090;
  wire _21092 = r1071 ^ _21091;
  wire _21093 = _12298 ? coded_block[1071] : r1071;
  wire _21094 = _12296 ? _21092 : _21093;
  always @ (posedge reset or posedge clock) if (reset) r1071 <= 1'd0; else if (_12300) r1071 <= _21094;
  wire [1:0] _21095 = {_0, _289} + {_0, _2974};
  wire [1:0] _21096 = {_0, _5310} + {_0, _6750};
  wire [2:0] _21097 = {_0, _21095} + {_0, _21096};
  wire [1:0] _21098 = {_0, _8638} + {_0, _10272};
  wire [3:0] _21099 = {_0, _21097} + {_0, _0, _21098};
  wire _21100 = _12301 < _21099;
  wire _21101 = r1070 ^ _21100;
  wire _21102 = _12298 ? coded_block[1070] : r1070;
  wire _21103 = _12296 ? _21101 : _21102;
  always @ (posedge reset or posedge clock) if (reset) r1070 <= 1'd0; else if (_12300) r1070 <= _21103;
  wire [1:0] _21104 = {_0, _320} + {_0, _2175};
  wire [1:0] _21105 = {_0, _5053} + {_0, _7389};
  wire [2:0] _21106 = {_0, _21104} + {_0, _21105};
  wire [1:0] _21107 = {_0, _8830} + {_0, _10717};
  wire [3:0] _21108 = {_0, _21106} + {_0, _0, _21107};
  wire _21109 = _12301 < _21108;
  wire _21110 = r1069 ^ _21109;
  wire _21111 = _12298 ? coded_block[1069] : r1069;
  wire _21112 = _12296 ? _21110 : _21111;
  always @ (posedge reset or posedge clock) if (reset) r1069 <= 1'd0; else if (_12300) r1069 <= _21112;
  wire [1:0] _21113 = {_0, _383} + {_0, _3037};
  wire [1:0] _21114 = {_0, _4319} + {_0, _6334};
  wire [2:0] _21115 = {_0, _21113} + {_0, _21114};
  wire [1:0] _21116 = {_0, _9212} + {_0, _11550};
  wire [3:0] _21117 = {_0, _21115} + {_0, _0, _21116};
  wire _21118 = _12301 < _21117;
  wire _21119 = r1068 ^ _21118;
  wire _21120 = _12298 ? coded_block[1068] : r1068;
  wire _21121 = _12296 ? _21119 : _21120;
  always @ (posedge reset or posedge clock) if (reset) r1068 <= 1'd0; else if (_12300) r1068 <= _21121;
  wire [1:0] _21122 = {_0, _416} + {_0, _3742};
  wire [1:0] _21123 = {_0, _5116} + {_0, _6397};
  wire [2:0] _21124 = {_0, _21122} + {_0, _21123};
  wire [1:0] _21125 = {_0, _8415} + {_0, _11295};
  wire [3:0] _21126 = {_0, _21124} + {_0, _0, _21125};
  wire _21127 = _12301 < _21126;
  wire _21128 = r1067 ^ _21127;
  wire _21129 = _12298 ? coded_block[1067] : r1067;
  wire _21130 = _12296 ? _21128 : _21129;
  always @ (posedge reset or posedge clock) if (reset) r1067 <= 1'd0; else if (_12300) r1067 <= _21130;
  wire [1:0] _21131 = {_0, _447} + {_0, _3646};
  wire [1:0] _21132 = {_0, _5821} + {_0, _7199};
  wire [2:0] _21133 = {_0, _21131} + {_0, _21132};
  wire [1:0] _21134 = {_0, _8480} + {_0, _10493};
  wire [3:0] _21135 = {_0, _21133} + {_0, _0, _21134};
  wire _21136 = _12301 < _21135;
  wire _21137 = r1066 ^ _21136;
  wire _21138 = _12298 ? coded_block[1066] : r1066;
  wire _21139 = _12296 ? _21137 : _21138;
  always @ (posedge reset or posedge clock) if (reset) r1066 <= 1'd0; else if (_12300) r1066 <= _21139;
  wire [1:0] _21140 = {_0, _479} + {_0, _2144};
  wire [1:0] _21141 = {_0, _5726} + {_0, _7900};
  wire [2:0] _21142 = {_0, _21140} + {_0, _21141};
  wire [1:0] _21143 = {_0, _9279} + {_0, _10558};
  wire [3:0] _21144 = {_0, _21142} + {_0, _0, _21143};
  wire _21145 = _12301 < _21144;
  wire _21146 = r1065 ^ _21145;
  wire _21147 = _12298 ? coded_block[1065] : r1065;
  wire _21148 = _12296 ? _21146 : _21147;
  always @ (posedge reset or posedge clock) if (reset) r1065 <= 1'd0; else if (_12300) r1065 <= _21148;
  wire [1:0] _21149 = {_0, _510} + {_0, _3005};
  wire [1:0] _21150 = {_0, _4223} + {_0, _7804};
  wire [2:0] _21151 = {_0, _21149} + {_0, _21150};
  wire [1:0] _21152 = {_0, _9980} + {_0, _11358};
  wire [3:0] _21153 = {_0, _21151} + {_0, _0, _21152};
  wire _21154 = _12301 < _21153;
  wire _21155 = r1064 ^ _21154;
  wire _21156 = _12298 ? coded_block[1064] : r1064;
  wire _21157 = _12296 ? _21155 : _21156;
  always @ (posedge reset or posedge clock) if (reset) r1064 <= 1'd0; else if (_12300) r1064 <= _21157;
  wire [1:0] _21158 = {_0, _545} + {_0, _2271};
  wire [1:0] _21159 = {_0, _5085} + {_0, _6303};
  wire [2:0] _21160 = {_0, _21158} + {_0, _21159};
  wire [1:0] _21161 = {_0, _9886} + {_0, _12061};
  wire [3:0] _21162 = {_0, _21160} + {_0, _0, _21161};
  wire _21163 = _12301 < _21162;
  wire _21164 = r1063 ^ _21163;
  wire _21165 = _12298 ? coded_block[1063] : r1063;
  wire _21166 = _12296 ? _21164 : _21165;
  always @ (posedge reset or posedge clock) if (reset) r1063 <= 1'd0; else if (_12300) r1063 <= _21166;
  wire [1:0] _21167 = {_0, _576} + {_0, _3325};
  wire [1:0] _21168 = {_0, _4350} + {_0, _7163};
  wire [2:0] _21169 = {_0, _21167} + {_0, _21168};
  wire [1:0] _21170 = {_0, _8383} + {_0, _11964};
  wire [3:0] _21171 = {_0, _21169} + {_0, _0, _21170};
  wire _21172 = _12301 < _21171;
  wire _21173 = r1062 ^ _21172;
  wire _21174 = _12298 ? coded_block[1062] : r1062;
  wire _21175 = _12296 ? _21173 : _21174;
  always @ (posedge reset or posedge clock) if (reset) r1062 <= 1'd0; else if (_12300) r1062 <= _21175;
  wire [1:0] _21176 = {_0, _608} + {_0, _3870};
  wire [1:0] _21177 = {_0, _5407} + {_0, _6431};
  wire [2:0] _21178 = {_0, _21176} + {_0, _21177};
  wire [1:0] _21179 = {_0, _9248} + {_0, _10462};
  wire [3:0] _21180 = {_0, _21178} + {_0, _0, _21179};
  wire _21181 = _12301 < _21180;
  wire _21182 = r1061 ^ _21181;
  wire _21183 = _12298 ? coded_block[1061] : r1061;
  wire _21184 = _12296 ? _21182 : _21183;
  always @ (posedge reset or posedge clock) if (reset) r1061 <= 1'd0; else if (_12300) r1061 <= _21184;
  wire [1:0] _21185 = {_0, _2044} + {_0, _3615};
  wire [1:0] _21186 = {_0, _5565} + {_0, _8123};
  wire [2:0] _21187 = {_0, _21185} + {_0, _21186};
  wire [1:0] _21188 = {_0, _9022} + {_0, _10335};
  wire [3:0] _21189 = {_0, _21187} + {_0, _0, _21188};
  wire _21190 = _12301 < _21189;
  wire _21191 = r1060 ^ _21190;
  wire _21192 = _12298 ? coded_block[1060] : r1060;
  wire _21193 = _12296 ? _21191 : _21192;
  always @ (posedge reset or posedge clock) if (reset) r1060 <= 1'd0; else if (_12300) r1060 <= _21193;
  wire [1:0] _21194 = {_0, _65} + {_0, _2941};
  wire [1:0] _21195 = {_0, _5694} + {_0, _7644};
  wire [2:0] _21196 = {_0, _21194} + {_0, _21195};
  wire [1:0] _21197 = {_0, _10204} + {_0, _11101};
  wire [3:0] _21198 = {_0, _21196} + {_0, _0, _21197};
  wire _21199 = _12301 < _21198;
  wire _21200 = r1059 ^ _21199;
  wire _21201 = _12298 ? coded_block[1059] : r1059;
  wire _21202 = _12296 ? _21200 : _21201;
  always @ (posedge reset or posedge clock) if (reset) r1059 <= 1'd0; else if (_12300) r1059 <= _21202;
  wire [1:0] _21203 = {_0, _863} + {_0, _2782};
  wire [1:0] _21204 = {_0, _4287} + {_0, _6589};
  wire [2:0] _21205 = {_0, _21203} + {_0, _21204};
  wire [1:0] _21206 = {_0, _9534} + {_0, _11228};
  wire [3:0] _21207 = {_0, _21205} + {_0, _0, _21206};
  wire _21208 = _12301 < _21207;
  wire _21209 = r1058 ^ _21208;
  wire _21210 = _12298 ? coded_block[1058] : r1058;
  wire _21211 = _12296 ? _21209 : _21210;
  always @ (posedge reset or posedge clock) if (reset) r1058 <= 1'd0; else if (_12300) r1058 <= _21211;
  wire [1:0] _21212 = {_0, _894} + {_0, _2719};
  wire [1:0] _21213 = {_0, _4861} + {_0, _6366};
  wire [2:0] _21214 = {_0, _21212} + {_0, _21213};
  wire [1:0] _21215 = {_0, _8670} + {_0, _11613};
  wire [3:0] _21216 = {_0, _21214} + {_0, _0, _21215};
  wire _21217 = _12301 < _21216;
  wire _21218 = r1057 ^ _21217;
  wire _21219 = _12298 ? coded_block[1057] : r1057;
  wire _21220 = _12296 ? _21218 : _21219;
  always @ (posedge reset or posedge clock) if (reset) r1057 <= 1'd0; else if (_12300) r1057 <= _21220;
  wire [1:0] _21221 = {_0, _927} + {_0, _3836};
  wire [1:0] _21222 = {_0, _4798} + {_0, _6942};
  wire [2:0] _21223 = {_0, _21221} + {_0, _21222};
  wire [1:0] _21224 = {_0, _8446} + {_0, _10748};
  wire [3:0] _21225 = {_0, _21223} + {_0, _0, _21224};
  wire _21226 = _12301 < _21225;
  wire _21227 = r1056 ^ _21226;
  wire _21228 = _12298 ? coded_block[1056] : r1056;
  wire _21229 = _12296 ? _21227 : _21228;
  always @ (posedge reset or posedge clock) if (reset) r1056 <= 1'd0; else if (_12300) r1056 <= _21229;
  wire [1:0] _21230 = {_0, _958} + {_0, _2494};
  wire [1:0] _21231 = {_0, _5918} + {_0, _6877};
  wire [2:0] _21232 = {_0, _21230} + {_0, _21231};
  wire [1:0] _21233 = {_0, _9022} + {_0, _10527};
  wire [3:0] _21234 = {_0, _21232} + {_0, _0, _21233};
  wire _21235 = _12301 < _21234;
  wire _21236 = r1055 ^ _21235;
  wire _21237 = _12298 ? coded_block[1055] : r1055;
  wire _21238 = _12296 ? _21236 : _21237;
  always @ (posedge reset or posedge clock) if (reset) r1055 <= 1'd0; else if (_12300) r1055 <= _21238;
  wire [1:0] _21239 = {_0, _990} + {_0, _4091};
  wire [1:0] _21240 = {_0, _4574} + {_0, _7996};
  wire [2:0] _21241 = {_0, _21239} + {_0, _21240};
  wire [1:0] _21242 = {_0, _8957} + {_0, _11101};
  wire [3:0] _21243 = {_0, _21241} + {_0, _0, _21242};
  wire _21244 = _12301 < _21243;
  wire _21245 = r1054 ^ _21244;
  wire _21246 = _12298 ? coded_block[1054] : r1054;
  wire _21247 = _12296 ? _21245 : _21246;
  always @ (posedge reset or posedge clock) if (reset) r1054 <= 1'd0; else if (_12300) r1054 <= _21247;
  wire [1:0] _21248 = {_0, _1021} + {_0, _3805};
  wire [1:0] _21249 = {_0, _4160} + {_0, _6652};
  wire [2:0] _21250 = {_0, _21248} + {_0, _21249};
  wire [1:0] _21251 = {_0, _10077} + {_0, _11038};
  wire [3:0] _21252 = {_0, _21250} + {_0, _0, _21251};
  wire _21253 = _12301 < _21252;
  wire _21254 = r1053 ^ _21253;
  wire _21255 = _12298 ? coded_block[1053] : r1053;
  wire _21256 = _12296 ? _21254 : _21255;
  always @ (posedge reset or posedge clock) if (reset) r1053 <= 1'd0; else if (_12300) r1053 <= _21256;
  wire [1:0] _21257 = {_0, _1057} + {_0, _2750};
  wire [1:0] _21258 = {_0, _5884} + {_0, _6239};
  wire [2:0] _21259 = {_0, _21257} + {_0, _21258};
  wire [1:0] _21260 = {_0, _8736} + {_0, _12155};
  wire [3:0] _21261 = {_0, _21259} + {_0, _0, _21260};
  wire _21262 = _12301 < _21261;
  wire _21263 = r1052 ^ _21262;
  wire _21264 = _12298 ? coded_block[1052] : r1052;
  wire _21265 = _12296 ? _21263 : _21264;
  always @ (posedge reset or posedge clock) if (reset) r1052 <= 1'd0; else if (_12300) r1052 <= _21265;
  wire [1:0] _21266 = {_0, _1088} + {_0, _2239};
  wire [1:0] _21267 = {_0, _4830} + {_0, _7965};
  wire [2:0] _21268 = {_0, _21266} + {_0, _21267};
  wire [1:0] _21269 = {_0, _8319} + {_0, _10814};
  wire [3:0] _21270 = {_0, _21268} + {_0, _0, _21269};
  wire _21271 = _12301 < _21270;
  wire _21272 = r1051 ^ _21271;
  wire _21273 = _12298 ? coded_block[1051] : r1051;
  wire _21274 = _12296 ? _21272 : _21273;
  always @ (posedge reset or posedge clock) if (reset) r1051 <= 1'd0; else if (_12300) r1051 <= _21274;
  wire [1:0] _21275 = {_0, _1120} + {_0, _3231};
  wire [1:0] _21276 = {_0, _4319} + {_0, _6908};
  wire [2:0] _21277 = {_0, _21275} + {_0, _21276};
  wire [1:0] _21278 = {_0, _10045} + {_0, _10399};
  wire [3:0] _21279 = {_0, _21277} + {_0, _0, _21278};
  wire _21280 = _12301 < _21279;
  wire _21281 = r1050 ^ _21280;
  wire _21282 = _12298 ? coded_block[1050] : r1050;
  wire _21283 = _12296 ? _21281 : _21282;
  always @ (posedge reset or posedge clock) if (reset) r1050 <= 1'd0; else if (_12300) r1050 <= _21283;
  wire [1:0] _21284 = {_0, _1151} + {_0, _3997};
  wire [1:0] _21285 = {_0, _5310} + {_0, _6397};
  wire [2:0] _21286 = {_0, _21284} + {_0, _21285};
  wire [1:0] _21287 = {_0, _8991} + {_0, _12124};
  wire [3:0] _21288 = {_0, _21286} + {_0, _0, _21287};
  wire _21289 = _12301 < _21288;
  wire _21290 = r1049 ^ _21289;
  wire _21291 = _12298 ? coded_block[1049] : r1049;
  wire _21292 = _12296 ? _21290 : _21291;
  always @ (posedge reset or posedge clock) if (reset) r1049 <= 1'd0; else if (_12300) r1049 <= _21292;
  wire [1:0] _21293 = {_0, _1184} + {_0, _3167};
  wire [1:0] _21294 = {_0, _6076} + {_0, _7389};
  wire [2:0] _21295 = {_0, _21293} + {_0, _21294};
  wire [1:0] _21296 = {_0, _8480} + {_0, _11069};
  wire [3:0] _21297 = {_0, _21295} + {_0, _0, _21296};
  wire _21298 = _12301 < _21297;
  wire _21299 = r1048 ^ _21298;
  wire _21300 = _12298 ? coded_block[1048] : r1048;
  wire _21301 = _12296 ? _21299 : _21300;
  always @ (posedge reset or posedge clock) if (reset) r1048 <= 1'd0; else if (_12300) r1048 <= _21301;
  wire [1:0] _21302 = {_0, _1215} + {_0, _2686};
  wire [1:0] _21303 = {_0, _5246} + {_0, _8155};
  wire [2:0] _21304 = {_0, _21302} + {_0, _21303};
  wire [1:0] _21305 = {_0, _9469} + {_0, _10558};
  wire [3:0] _21306 = {_0, _21304} + {_0, _0, _21305};
  wire _21307 = _12301 < _21306;
  wire _21308 = r1047 ^ _21307;
  wire _21309 = _12298 ? coded_block[1047] : r1047;
  wire _21310 = _12296 ? _21308 : _21309;
  always @ (posedge reset or posedge clock) if (reset) r1047 <= 1'd0; else if (_12300) r1047 <= _21310;
  wire [1:0] _21311 = {_0, _1247} + {_0, _2813};
  wire [1:0] _21312 = {_0, _4767} + {_0, _7326};
  wire [2:0] _21313 = {_0, _21311} + {_0, _21312};
  wire [1:0] _21314 = {_0, _10235} + {_0, _11550};
  wire [3:0] _21315 = {_0, _21313} + {_0, _0, _21314};
  wire _21316 = _12301 < _21315;
  wire _21317 = r1046 ^ _21316;
  wire _21318 = _12298 ? coded_block[1046] : r1046;
  wire _21319 = _12296 ? _21317 : _21318;
  always @ (posedge reset or posedge clock) if (reset) r1046 <= 1'd0; else if (_12300) r1046 <= _21319;
  wire [1:0] _21320 = {_0, _1278} + {_0, _2144};
  wire [1:0] _21321 = {_0, _4895} + {_0, _6845};
  wire [2:0] _21322 = {_0, _21320} + {_0, _21321};
  wire [1:0] _21323 = {_0, _9406} + {_0, _10303};
  wire [3:0] _21324 = {_0, _21322} + {_0, _0, _21323};
  wire _21325 = _12301 < _21324;
  wire _21326 = r1045 ^ _21325;
  wire _21327 = _12298 ? coded_block[1045] : r1045;
  wire _21328 = _12296 ? _21326 : _21327;
  always @ (posedge reset or posedge clock) if (reset) r1045 <= 1'd0; else if (_12300) r1045 <= _21328;
  wire [1:0] _21329 = {_0, _1312} + {_0, _3390};
  wire [1:0] _21330 = {_0, _4223} + {_0, _6973};
  wire [2:0] _21331 = {_0, _21329} + {_0, _21330};
  wire [1:0] _21332 = {_0, _8926} + {_0, _11485};
  wire [3:0] _21333 = {_0, _21331} + {_0, _0, _21332};
  wire _21334 = _12301 < _21333;
  wire _21335 = r1044 ^ _21334;
  wire _21336 = _12298 ? coded_block[1044] : r1044;
  wire _21337 = _12296 ? _21335 : _21336;
  always @ (posedge reset or posedge clock) if (reset) r1044 <= 1'd0; else if (_12300) r1044 <= _21337;
  wire [1:0] _21338 = {_0, _1343} + {_0, _3359};
  wire [1:0] _21339 = {_0, _5470} + {_0, _6303};
  wire [2:0] _21340 = {_0, _21338} + {_0, _21339};
  wire [1:0] _21341 = {_0, _9054} + {_0, _11004};
  wire [3:0] _21342 = {_0, _21340} + {_0, _0, _21341};
  wire _21343 = _12301 < _21342;
  wire _21344 = r1043 ^ _21343;
  wire _21345 = _12298 ? coded_block[1043] : r1043;
  wire _21346 = _12296 ? _21344 : _21345;
  always @ (posedge reset or posedge clock) if (reset) r1043 <= 1'd0; else if (_12300) r1043 <= _21346;
  wire [1:0] _21347 = {_0, _1375} + {_0, _2175};
  wire [1:0] _21348 = {_0, _5438} + {_0, _7548};
  wire [2:0] _21349 = {_0, _21347} + {_0, _21348};
  wire [1:0] _21350 = {_0, _8383} + {_0, _11132};
  wire [3:0] _21351 = {_0, _21349} + {_0, _0, _21350};
  wire _21352 = _12301 < _21351;
  wire _21353 = r1042 ^ _21352;
  wire _21354 = _12298 ? coded_block[1042] : r1042;
  wire _21355 = _12296 ? _21353 : _21354;
  always @ (posedge reset or posedge clock) if (reset) r1042 <= 1'd0; else if (_12300) r1042 <= _21355;
  wire [1:0] _21356 = {_0, _1406} + {_0, _2463};
  wire [1:0] _21357 = {_0, _4256} + {_0, _7517};
  wire [2:0] _21358 = {_0, _21356} + {_0, _21357};
  wire [1:0] _21359 = {_0, _9630} + {_0, _10462};
  wire [3:0] _21360 = {_0, _21358} + {_0, _0, _21359};
  wire _21361 = _12301 < _21360;
  wire _21362 = r1041 ^ _21361;
  wire _21363 = _12298 ? coded_block[1041] : r1041;
  wire _21364 = _12296 ? _21362 : _21363;
  always @ (posedge reset or posedge clock) if (reset) r1041 <= 1'd0; else if (_12300) r1041 <= _21364;
  wire [1:0] _21365 = {_0, _1439} + {_0, _3870};
  wire [1:0] _21366 = {_0, _4542} + {_0, _6334};
  wire [2:0] _21367 = {_0, _21365} + {_0, _21366};
  wire [1:0] _21368 = {_0, _9597} + {_0, _11708};
  wire [3:0] _21369 = {_0, _21367} + {_0, _0, _21368};
  wire _21370 = _12301 < _21369;
  wire _21371 = r1040 ^ _21370;
  wire _21372 = _12298 ? coded_block[1040] : r1040;
  wire _21373 = _12296 ? _21371 : _21372;
  always @ (posedge reset or posedge clock) if (reset) r1040 <= 1'd0; else if (_12300) r1040 <= _21373;
  wire [1:0] _21374 = {_0, _1470} + {_0, _3709};
  wire [1:0] _21375 = {_0, _5949} + {_0, _6621};
  wire [2:0] _21376 = {_0, _21374} + {_0, _21375};
  wire [1:0] _21377 = {_0, _8415} + {_0, _11677};
  wire [3:0] _21378 = {_0, _21376} + {_0, _0, _21377};
  wire _21379 = _12301 < _21378;
  wire _21380 = r1039 ^ _21379;
  wire _21381 = _12298 ? coded_block[1039] : r1039;
  wire _21382 = _12296 ? _21380 : _21381;
  always @ (posedge reset or posedge clock) if (reset) r1039 <= 1'd0; else if (_12300) r1039 <= _21382;
  wire [1:0] _21383 = {_0, _1502} + {_0, _2081};
  wire [1:0] _21384 = {_0, _5790} + {_0, _8028};
  wire [2:0] _21385 = {_0, _21383} + {_0, _21384};
  wire [1:0] _21386 = {_0, _8701} + {_0, _10493};
  wire [3:0] _21387 = {_0, _21385} + {_0, _0, _21386};
  wire _21388 = _12301 < _21387;
  wire _21389 = r1038 ^ _21388;
  wire _21390 = _12298 ? coded_block[1038] : r1038;
  wire _21391 = _12296 ? _21389 : _21390;
  always @ (posedge reset or posedge clock) if (reset) r1038 <= 1'd0; else if (_12300) r1038 <= _21391;
  wire [1:0] _21392 = {_0, _1533} + {_0, _3742};
  wire [1:0] _21393 = {_0, _4129} + {_0, _7868};
  wire [2:0] _21394 = {_0, _21392} + {_0, _21393};
  wire [1:0] _21395 = {_0, _10108} + {_0, _10783};
  wire [3:0] _21396 = {_0, _21394} + {_0, _0, _21395};
  wire _21397 = _12301 < _21396;
  wire _21398 = r1037 ^ _21397;
  wire _21399 = _12298 ? coded_block[1037] : r1037;
  wire _21400 = _12296 ? _21398 : _21399;
  always @ (posedge reset or posedge clock) if (reset) r1037 <= 1'd0; else if (_12300) r1037 <= _21400;
  wire [1:0] _21401 = {_0, _1568} + {_0, _3933};
  wire [1:0] _21402 = {_0, _5821} + {_0, _6176};
  wire [2:0] _21403 = {_0, _21401} + {_0, _21402};
  wire [1:0] _21404 = {_0, _9949} + {_0, _12188};
  wire [3:0] _21405 = {_0, _21403} + {_0, _0, _21404};
  wire _21406 = _12301 < _21405;
  wire _21407 = r1036 ^ _21406;
  wire _21408 = _12298 ? coded_block[1036] : r1036;
  wire _21409 = _12296 ? _21407 : _21408;
  always @ (posedge reset or posedge clock) if (reset) r1036 <= 1'd0; else if (_12300) r1036 <= _21409;
  wire [1:0] _21410 = {_0, _1599} + {_0, _2557};
  wire [1:0] _21411 = {_0, _6012} + {_0, _7900};
  wire [2:0] _21412 = {_0, _21410} + {_0, _21411};
  wire [1:0] _21413 = {_0, _8225} + {_0, _12027};
  wire [3:0] _21414 = {_0, _21412} + {_0, _0, _21413};
  wire _21415 = _12301 < _21414;
  wire _21416 = r1035 ^ _21415;
  wire _21417 = _12298 ? coded_block[1035] : r1035;
  wire _21418 = _12296 ? _21416 : _21417;
  always @ (posedge reset or posedge clock) if (reset) r1035 <= 1'd0; else if (_12300) r1035 <= _21418;
  wire [1:0] _21419 = {_0, _1631} + {_0, _2302};
  wire [1:0] _21420 = {_0, _4640} + {_0, _8092};
  wire [2:0] _21421 = {_0, _21419} + {_0, _21420};
  wire [1:0] _21422 = {_0, _9980} + {_0, _10272};
  wire [3:0] _21423 = {_0, _21421} + {_0, _0, _21422};
  wire _21424 = _12301 < _21423;
  wire _21425 = r1034 ^ _21424;
  wire _21426 = _12298 ? coded_block[1034] : r1034;
  wire _21427 = _12296 ? _21425 : _21426;
  always @ (posedge reset or posedge clock) if (reset) r1034 <= 1'd0; else if (_12300) r1034 <= _21427;
  wire [1:0] _21428 = {_0, _1695} + {_0, _3580};
  wire [1:0] _21429 = {_0, _5597} + {_0, _6462};
  wire [2:0] _21430 = {_0, _21428} + {_0, _21429};
  wire [1:0] _21431 = {_0, _8799} + {_0, _12251};
  wire [3:0] _21432 = {_0, _21430} + {_0, _0, _21431};
  wire _21433 = _12301 < _21432;
  wire _21434 = r1033 ^ _21433;
  wire _21435 = _12298 ? coded_block[1033] : r1033;
  wire _21436 = _12296 ? _21434 : _21435;
  always @ (posedge reset or posedge clock) if (reset) r1033 <= 1'd0; else if (_12300) r1033 <= _21436;
  wire [1:0] _21437 = {_0, _1726} + {_0, _2367};
  wire [1:0] _21438 = {_0, _5663} + {_0, _7675};
  wire [2:0] _21439 = {_0, _21437} + {_0, _21438};
  wire [1:0] _21440 = {_0, _8543} + {_0, _10877};
  wire [3:0] _21441 = {_0, _21439} + {_0, _0, _21440};
  wire _21442 = _12301 < _21441;
  wire _21443 = r1032 ^ _21442;
  wire _21444 = _12298 ? coded_block[1032] : r1032;
  wire _21445 = _12296 ? _21443 : _21444;
  always @ (posedge reset or posedge clock) if (reset) r1032 <= 1'd0; else if (_12300) r1032 <= _21445;
  wire [1:0] _21446 = {_0, _1758} + {_0, _3068};
  wire [1:0] _21447 = {_0, _4447} + {_0, _7741};
  wire [2:0] _21448 = {_0, _21446} + {_0, _21447};
  wire [1:0] _21449 = {_0, _9759} + {_0, _10621};
  wire [3:0] _21450 = {_0, _21448} + {_0, _0, _21449};
  wire _21451 = _12301 < _21450;
  wire _21452 = r1031 ^ _21451;
  wire _21453 = _12298 ? coded_block[1031] : r1031;
  wire _21454 = _12296 ? _21452 : _21453;
  always @ (posedge reset or posedge clock) if (reset) r1031 <= 1'd0; else if (_12300) r1031 <= _21454;
  wire [1:0] _21455 = {_0, _1789} + {_0, _2974};
  wire [1:0] _21456 = {_0, _5152} + {_0, _6525};
  wire [2:0] _21457 = {_0, _21455} + {_0, _21456};
  wire [1:0] _21458 = {_0, _9822} + {_0, _11837};
  wire [3:0] _21459 = {_0, _21457} + {_0, _0, _21458};
  wire _21460 = _12301 < _21459;
  wire _21461 = r1030 ^ _21460;
  wire _21462 = _12298 ? coded_block[1030] : r1030;
  wire _21463 = _12296 ? _21461 : _21462;
  always @ (posedge reset or posedge clock) if (reset) r1030 <= 1'd0; else if (_12300) r1030 <= _21463;
  wire [1:0] _21464 = {_0, _1823} + {_0, _3486};
  wire [1:0] _21465 = {_0, _5053} + {_0, _7230};
  wire [2:0] _21466 = {_0, _21464} + {_0, _21465};
  wire [1:0] _21467 = {_0, _8607} + {_0, _11900};
  wire [3:0] _21468 = {_0, _21466} + {_0, _0, _21467};
  wire _21469 = _12301 < _21468;
  wire _21470 = r1029 ^ _21469;
  wire _21471 = _12298 ? coded_block[1029] : r1029;
  wire _21472 = _12296 ? _21470 : _21471;
  always @ (posedge reset or posedge clock) if (reset) r1029 <= 1'd0; else if (_12300) r1029 <= _21472;
  wire [1:0] _21473 = {_0, _1886} + {_0, _3615};
  wire [1:0] _21474 = {_0, _4415} + {_0, _7644};
  wire [2:0] _21475 = {_0, _21473} + {_0, _21474};
  wire [1:0] _21476 = {_0, _9212} + {_0, _11389};
  wire [3:0] _21477 = {_0, _21475} + {_0, _0, _21476};
  wire _21478 = _12301 < _21477;
  wire _21479 = r1028 ^ _21478;
  wire _21480 = _12298 ? coded_block[1028] : r1028;
  wire _21481 = _12296 ? _21479 : _21480;
  always @ (posedge reset or posedge clock) if (reset) r1028 <= 1'd0; else if (_12300) r1028 <= _21481;
  wire [1:0] _21482 = {_0, _1917} + {_0, _2655};
  wire [1:0] _21483 = {_0, _5694} + {_0, _6494};
  wire [2:0] _21484 = {_0, _21482} + {_0, _21483};
  wire [1:0] _21485 = {_0, _9724} + {_0, _11295};
  wire [3:0] _21486 = {_0, _21484} + {_0, _0, _21485};
  wire _21487 = _12301 < _21486;
  wire _21488 = r1027 ^ _21487;
  wire _21489 = _12298 ? coded_block[1027] : r1027;
  wire _21490 = _12296 ? _21488 : _21489;
  always @ (posedge reset or posedge clock) if (reset) r1027 <= 1'd0; else if (_12300) r1027 <= _21490;
  wire [1:0] _21491 = {_0, _1950} + {_0, _3198};
  wire [1:0] _21492 = {_0, _4734} + {_0, _7773};
  wire [2:0] _21493 = {_0, _21491} + {_0, _21492};
  wire [1:0] _21494 = {_0, _8574} + {_0, _11806};
  wire [3:0] _21495 = {_0, _21493} + {_0, _0, _21494};
  wire _21496 = _12301 < _21495;
  wire _21497 = r1026 ^ _21496;
  wire _21498 = _12298 ? coded_block[1026] : r1026;
  wire _21499 = _12296 ? _21497 : _21498;
  always @ (posedge reset or posedge clock) if (reset) r1026 <= 1'd0; else if (_12300) r1026 <= _21499;
  wire [1:0] _21500 = {_0, _1981} + {_0, _2271};
  wire [1:0] _21501 = {_0, _5279} + {_0, _6814};
  wire [2:0] _21502 = {_0, _21500} + {_0, _21501};
  wire [1:0] _21503 = {_0, _9853} + {_0, _10654};
  wire [3:0] _21504 = {_0, _21502} + {_0, _0, _21503};
  wire _21505 = _12301 < _21504;
  wire _21506 = r1025 ^ _21505;
  wire _21507 = _12298 ? coded_block[1025] : r1025;
  wire _21508 = _12296 ? _21506 : _21507;
  always @ (posedge reset or posedge clock) if (reset) r1025 <= 1'd0; else if (_12300) r1025 <= _21508;
  wire [1:0] _21509 = {_0, _2044} + {_0, _3037};
  wire [1:0] _21510 = {_0, _4671} + {_0, _6431};
  wire [2:0] _21511 = {_0, _21509} + {_0, _21510};
  wire [1:0] _21512 = {_0, _9438} + {_0, _10973};
  wire [3:0] _21513 = {_0, _21511} + {_0, _0, _21512};
  wire _21514 = _12301 < _21513;
  wire _21515 = r1024 ^ _21514;
  wire _21516 = _12298 ? coded_block[1024] : r1024;
  wire _21517 = _12296 ? _21515 : _21516;
  always @ (posedge reset or posedge clock) if (reset) r1024 <= 1'd0; else if (_12300) r1024 <= _21517;
  wire [1:0] _21518 = {_0, _65} + {_0, _2399};
  wire [1:0] _21519 = {_0, _5116} + {_0, _6750};
  wire [2:0] _21520 = {_0, _21518} + {_0, _21519};
  wire [1:0] _21521 = {_0, _8511} + {_0, _11516};
  wire [3:0] _21522 = {_0, _21520} + {_0, _0, _21521};
  wire _21523 = _12301 < _21522;
  wire _21524 = r1023 ^ _21523;
  wire _21525 = _12298 ? coded_block[1023] : r1023;
  wire _21526 = _12296 ? _21524 : _21525;
  always @ (posedge reset or posedge clock) if (reset) r1023 <= 1'd0; else if (_12300) r1023 <= _21526;
  wire [1:0] _21527 = {_0, _97} + {_0, _3325};
  wire [1:0] _21528 = {_0, _4478} + {_0, _7199};
  wire [2:0] _21529 = {_0, _21527} + {_0, _21528};
  wire [1:0] _21530 = {_0, _8830} + {_0, _10590};
  wire [3:0] _21531 = {_0, _21529} + {_0, _0, _21530};
  wire _21532 = _12301 < _21531;
  wire _21533 = r1022 ^ _21532;
  wire _21534 = _12298 ? coded_block[1022] : r1022;
  wire _21535 = _12296 ? _21533 : _21534;
  always @ (posedge reset or posedge clock) if (reset) r1022 <= 1'd0; else if (_12300) r1022 <= _21535;
  wire [1:0] _21536 = {_0, _128} + {_0, _3422};
  wire [1:0] _21537 = {_0, _5407} + {_0, _6558};
  wire [2:0] _21538 = {_0, _21536} + {_0, _21537};
  wire [1:0] _21539 = {_0, _9279} + {_0, _10910};
  wire [3:0] _21540 = {_0, _21538} + {_0, _0, _21539};
  wire _21541 = _12301 < _21540;
  wire _21542 = r1021 ^ _21541;
  wire _21543 = _12298 ? coded_block[1021] : r1021;
  wire _21544 = _12296 ? _21542 : _21543;
  always @ (posedge reset or posedge clock) if (reset) r1021 <= 1'd0; else if (_12300) r1021 <= _21544;
  wire [1:0] _21545 = {_0, _192} + {_0, _3135};
  wire [1:0] _21546 = {_0, _4958} + {_0, _7581};
  wire [2:0] _21547 = {_0, _21545} + {_0, _21546};
  wire [1:0] _21548 = {_0, _9566} + {_0, _10717};
  wire [3:0] _21549 = {_0, _21547} + {_0, _0, _21548};
  wire _21550 = _12301 < _21549;
  wire _21551 = r1020 ^ _21550;
  wire _21552 = _12298 ? coded_block[1020] : r1020;
  wire _21553 = _12296 ? _21551 : _21552;
  always @ (posedge reset or posedge clock) if (reset) r1020 <= 1'd0; else if (_12300) r1020 <= _21553;
  wire [1:0] _21554 = {_0, _224} + {_0, _4028};
  wire [1:0] _21555 = {_0, _5215} + {_0, _7036};
  wire [2:0] _21556 = {_0, _21554} + {_0, _21555};
  wire [1:0] _21557 = {_0, _9661} + {_0, _11644};
  wire [3:0] _21558 = {_0, _21556} + {_0, _0, _21557};
  wire _21559 = _12301 < _21558;
  wire _21560 = r1019 ^ _21559;
  wire _21561 = _12298 ? coded_block[1019] : r1019;
  wire _21562 = _12296 ? _21560 : _21561;
  always @ (posedge reset or posedge clock) if (reset) r1019 <= 1'd0; else if (_12300) r1019 <= _21562;
  wire [1:0] _21563 = {_0, _255} + {_0, _3678};
  wire [1:0] _21564 = {_0, _6108} + {_0, _7293};
  wire [2:0] _21565 = {_0, _21563} + {_0, _21564};
  wire [1:0] _21566 = {_0, _9118} + {_0, _11740};
  wire [3:0] _21567 = {_0, _21565} + {_0, _0, _21566};
  wire _21568 = _12301 < _21567;
  wire _21569 = r1018 ^ _21568;
  wire _21570 = _12298 ? coded_block[1018] : r1018;
  wire _21571 = _12296 ? _21569 : _21570;
  always @ (posedge reset or posedge clock) if (reset) r1018 <= 1'd0; else if (_12300) r1018 <= _21571;
  wire [1:0] _21572 = {_0, _289} + {_0, _3901};
  wire [1:0] _21573 = {_0, _5757} + {_0, _8186};
  wire [2:0] _21574 = {_0, _21572} + {_0, _21573};
  wire [1:0] _21575 = {_0, _9375} + {_0, _11196};
  wire [3:0] _21576 = {_0, _21574} + {_0, _0, _21575};
  wire _21577 = _12301 < _21576;
  wire _21578 = r1017 ^ _21577;
  wire _21579 = _12298 ? coded_block[1017] : r1017;
  wire _21580 = _12296 ? _21578 : _21579;
  always @ (posedge reset or posedge clock) if (reset) r1017 <= 1'd0; else if (_12300) r1017 <= _21580;
  wire [1:0] _21581 = {_0, _320} + {_0, _3773};
  wire [1:0] _21582 = {_0, _5981} + {_0, _7837};
  wire [2:0] _21583 = {_0, _21581} + {_0, _21582};
  wire [1:0] _21584 = {_0, _8256} + {_0, _11453};
  wire [3:0] _21585 = {_0, _21583} + {_0, _0, _21584};
  wire _21586 = _12301 < _21585;
  wire _21587 = r1016 ^ _21586;
  wire _21588 = _12298 ? coded_block[1016] : r1016;
  wire _21589 = _12296 ? _21587 : _21588;
  always @ (posedge reset or posedge clock) if (reset) r1016 <= 1'd0; else if (_12300) r1016 <= _21589;
  wire [1:0] _21590 = {_0, _352} + {_0, _2112};
  wire [1:0] _21591 = {_0, _5853} + {_0, _8059};
  wire [2:0] _21592 = {_0, _21590} + {_0, _21591};
  wire [1:0] _21593 = {_0, _9917} + {_0, _10335};
  wire [3:0] _21594 = {_0, _21592} + {_0, _0, _21593};
  wire _21595 = _12301 < _21594;
  wire _21596 = r1015 ^ _21595;
  wire _21597 = _12298 ? coded_block[1015] : r1015;
  wire _21598 = _12296 ? _21596 : _21597;
  always @ (posedge reset or posedge clock) if (reset) r1015 <= 1'd0; else if (_12300) r1015 <= _21598;
  wire [1:0] _21599 = {_0, _383} + {_0, _2847};
  wire [1:0] _21600 = {_0, _4192} + {_0, _7931};
  wire [2:0] _21601 = {_0, _21599} + {_0, _21600};
  wire [1:0] _21602 = {_0, _10141} + {_0, _11996};
  wire [3:0] _21603 = {_0, _21601} + {_0, _0, _21602};
  wire _21604 = _12301 < _21603;
  wire _21605 = r1014 ^ _21604;
  wire _21606 = _12298 ? coded_block[1014] : r1014;
  wire _21607 = _12296 ? _21605 : _21606;
  always @ (posedge reset or posedge clock) if (reset) r1014 <= 1'd0; else if (_12300) r1014 <= _21607;
  wire [1:0] _21608 = {_0, _447} + {_0, _3005};
  wire [1:0] _21609 = {_0, _5534} + {_0, _7005};
  wire [2:0] _21610 = {_0, _21608} + {_0, _21609};
  wire [1:0] _21611 = {_0, _8352} + {_0, _12092};
  wire [3:0] _21612 = {_0, _21610} + {_0, _0, _21611};
  wire _21613 = _12301 < _21612;
  wire _21614 = r1013 ^ _21613;
  wire _21615 = _12298 ? coded_block[1013] : r1013;
  wire _21616 = _12296 ? _21614 : _21615;
  always @ (posedge reset or posedge clock) if (reset) r1013 <= 1'd0; else if (_12300) r1013 <= _21616;
  wire [1:0] _21617 = {_0, _479} + {_0, _2623};
  wire [1:0] _21618 = {_0, _5085} + {_0, _7612};
  wire [2:0] _21619 = {_0, _21617} + {_0, _21618};
  wire [1:0] _21620 = {_0, _9085} + {_0, _10430};
  wire [3:0] _21621 = {_0, _21619} + {_0, _0, _21620};
  wire _21622 = _12301 < _21621;
  wire _21623 = r1012 ^ _21622;
  wire _21624 = _12298 ? coded_block[1012] : r1012;
  wire _21625 = _12296 ? _21623 : _21624;
  always @ (posedge reset or posedge clock) if (reset) r1012 <= 1'd0; else if (_12300) r1012 <= _21625;
  wire [1:0] _21626 = {_0, _510} + {_0, _3646};
  wire [1:0] _21627 = {_0, _4703} + {_0, _7163};
  wire [2:0] _21628 = {_0, _21626} + {_0, _21627};
  wire [1:0] _21629 = {_0, _9693} + {_0, _11165};
  wire [3:0] _21630 = {_0, _21628} + {_0, _0, _21629};
  wire _21631 = _12301 < _21630;
  wire _21632 = r1011 ^ _21631;
  wire _21633 = _12298 ? coded_block[1011] : r1011;
  wire _21634 = _12296 ? _21632 : _21633;
  always @ (posedge reset or posedge clock) if (reset) r1011 <= 1'd0; else if (_12300) r1011 <= _21634;
  wire [1:0] _21635 = {_0, _545} + {_0, _4060};
  wire [1:0] _21636 = {_0, _5726} + {_0, _6781};
  wire [2:0] _21637 = {_0, _21635} + {_0, _21636};
  wire [1:0] _21638 = {_0, _9248} + {_0, _11771};
  wire [3:0] _21639 = {_0, _21637} + {_0, _0, _21638};
  wire _21640 = _12301 < _21639;
  wire _21641 = r1010 ^ _21640;
  wire _21642 = _12298 ? coded_block[1010] : r1010;
  wire _21643 = _12296 ? _21641 : _21642;
  always @ (posedge reset or posedge clock) if (reset) r1010 <= 1'd0; else if (_12300) r1010 <= _21643;
  wire [1:0] _21644 = {_0, _576} + {_0, _2526};
  wire [1:0] _21645 = {_0, _6139} + {_0, _7804};
  wire [2:0] _21646 = {_0, _21644} + {_0, _21645};
  wire [1:0] _21647 = {_0, _8863} + {_0, _11326};
  wire [3:0] _21648 = {_0, _21646} + {_0, _0, _21647};
  wire _21649 = _12301 < _21648;
  wire _21650 = r1009 ^ _21649;
  wire _21651 = _12298 ? coded_block[1009] : r1009;
  wire _21652 = _12296 ? _21650 : _21651;
  always @ (posedge reset or posedge clock) if (reset) r1009 <= 1'd0; else if (_12300) r1009 <= _21652;
  wire [1:0] _21653 = {_0, _608} + {_0, _3964};
  wire [1:0] _21654 = {_0, _4605} + {_0, _6207};
  wire [2:0] _21655 = {_0, _21653} + {_0, _21654};
  wire [1:0] _21656 = {_0, _9886} + {_0, _10941};
  wire [3:0] _21657 = {_0, _21655} + {_0, _0, _21656};
  wire _21658 = _12301 < _21657;
  wire _21659 = r1008 ^ _21658;
  wire _21660 = _12298 ? coded_block[1008] : r1008;
  wire _21661 = _12296 ? _21659 : _21660;
  always @ (posedge reset or posedge clock) if (reset) r1008 <= 1'd0; else if (_12300) r1008 <= _21661;
  wire [1:0] _21662 = {_0, _672} + {_0, _2941};
  wire [1:0] _21663 = {_0, _5342} + {_0, _8123};
  wire [2:0] _21664 = {_0, _21662} + {_0, _21663};
  wire [1:0] _21665 = {_0, _8767} + {_0, _10366};
  wire [3:0] _21666 = {_0, _21664} + {_0, _0, _21665};
  wire _21667 = _12301 < _21666;
  wire _21668 = r1007 ^ _21667;
  wire _21669 = _12298 ? coded_block[1007] : r1007;
  wire _21670 = _12296 ? _21668 : _21669;
  always @ (posedge reset or posedge clock) if (reset) r1007 <= 1'd0; else if (_12300) r1007 <= _21670;
  wire [1:0] _21671 = {_0, _703} + {_0, _3104};
  wire [1:0] _21672 = {_0, _5022} + {_0, _7420};
  wire [2:0] _21673 = {_0, _21671} + {_0, _21672};
  wire [1:0] _21674 = {_0, _10204} + {_0, _10846};
  wire [3:0] _21675 = {_0, _21673} + {_0, _0, _21674};
  wire _21676 = _12301 < _21675;
  wire _21677 = r1006 ^ _21676;
  wire _21678 = _12298 ? coded_block[1006] : r1006;
  wire _21679 = _12296 ? _21677 : _21678;
  always @ (posedge reset or posedge clock) if (reset) r1006 <= 1'd0; else if (_12300) r1006 <= _21679;
  wire [1:0] _21680 = {_0, _766} + {_0, _3294};
  wire [1:0] _21681 = {_0, _4989} + {_0, _7262};
  wire [2:0] _21682 = {_0, _21680} + {_0, _21681};
  wire [1:0] _21683 = {_0, _9181} + {_0, _11581};
  wire [3:0] _21684 = {_0, _21682} + {_0, _0, _21683};
  wire _21685 = _12301 < _21684;
  wire _21686 = r1005 ^ _21685;
  wire _21687 = _12298 ? coded_block[1005] : r1005;
  wire _21688 = _12296 ? _21686 : _21687;
  always @ (posedge reset or posedge clock) if (reset) r1005 <= 1'd0; else if (_12300) r1005 <= _21688;
  wire [1:0] _21689 = {_0, _800} + {_0, _2430};
  wire [1:0] _21690 = {_0, _5373} + {_0, _7069};
  wire [2:0] _21691 = {_0, _21689} + {_0, _21690};
  wire [1:0] _21692 = {_0, _9342} + {_0, _11259};
  wire [3:0] _21693 = {_0, _21691} + {_0, _0, _21692};
  wire _21694 = _12301 < _21693;
  wire _21695 = r1004 ^ _21694;
  wire _21696 = _12298 ? coded_block[1004] : r1004;
  wire _21697 = _12296 ? _21695 : _21696;
  always @ (posedge reset or posedge clock) if (reset) r1004 <= 1'd0; else if (_12300) r1004 <= _21697;
  wire [1:0] _21698 = {_0, _97} + {_0, _2175};
  wire [1:0] _21699 = {_0, _5022} + {_0, _7773};
  wire [2:0] _21700 = {_0, _21698} + {_0, _21699};
  wire [1:0] _21701 = {_0, _9724} + {_0, _12282};
  wire [3:0] _21702 = {_0, _21700} + {_0, _0, _21701};
  wire _21703 = _12301 < _21702;
  wire _21704 = r1003 ^ _21703;
  wire _21705 = _12298 ? coded_block[1003] : r1003;
  wire _21706 = _12296 ? _21704 : _21705;
  always @ (posedge reset or posedge clock) if (reset) r1003 <= 1'd0; else if (_12300) r1003 <= _21706;
  wire [1:0] _21707 = {_0, _1631} + {_0, _3836};
  wire [1:0] _21708 = {_0, _4129} + {_0, _7965};
  wire [2:0] _21709 = {_0, _21707} + {_0, _21708};
  wire [1:0] _21710 = {_0, _10204} + {_0, _10877};
  wire [3:0] _21711 = {_0, _21709} + {_0, _0, _21710};
  wire _21712 = _12301 < _21711;
  wire _21713 = r1002 ^ _21712;
  wire _21714 = _12298 ? coded_block[1002] : r1002;
  wire _21715 = _12296 ? _21713 : _21714;
  always @ (posedge reset or posedge clock) if (reset) r1002 <= 1'd0; else if (_12300) r1002 <= _21715;
  wire [1:0] _21716 = {_0, _1662} + {_0, _4028};
  wire [1:0] _21717 = {_0, _5918} + {_0, _6176};
  wire [2:0] _21718 = {_0, _21716} + {_0, _21717};
  wire [1:0] _21719 = {_0, _10045} + {_0, _12282};
  wire [3:0] _21720 = {_0, _21718} + {_0, _0, _21719};
  wire _21721 = _12301 < _21720;
  wire _21722 = r1001 ^ _21721;
  wire _21723 = _12298 ? coded_block[1001] : r1001;
  wire _21724 = _12296 ? _21722 : _21723;
  always @ (posedge reset or posedge clock) if (reset) r1001 <= 1'd0; else if (_12300) r1001 <= _21724;
  wire [1:0] _21725 = {_0, _1695} + {_0, _2655};
  wire [1:0] _21726 = {_0, _6108} + {_0, _7996};
  wire [2:0] _21727 = {_0, _21725} + {_0, _21726};
  wire [1:0] _21728 = {_0, _8225} + {_0, _12124};
  wire [3:0] _21729 = {_0, _21727} + {_0, _0, _21728};
  wire _21730 = _12301 < _21729;
  wire _21731 = r1000 ^ _21730;
  wire _21732 = _12298 ? coded_block[1000] : r1000;
  wire _21733 = _12296 ? _21731 : _21732;
  always @ (posedge reset or posedge clock) if (reset) r1000 <= 1'd0; else if (_12300) r1000 <= _21733;
  wire [1:0] _21734 = {_0, _1758} + {_0, _3615};
  wire [1:0] _21735 = {_0, _4478} + {_0, _6814};
  wire [2:0] _21736 = {_0, _21734} + {_0, _21735};
  wire [1:0] _21737 = {_0, _8256} + {_0, _12155};
  wire [3:0] _21738 = {_0, _21736} + {_0, _0, _21737};
  wire _21739 = _12301 < _21738;
  wire _21740 = r999 ^ _21739;
  wire _21741 = _12298 ? coded_block[999] : r999;
  wire _21742 = _12296 ? _21740 : _21741;
  always @ (posedge reset or posedge clock) if (reset) r999 <= 1'd0; else if (_12300) r999 <= _21742;
  wire [1:0] _21743 = {_0, _1789} + {_0, _3678};
  wire [1:0] _21744 = {_0, _5694} + {_0, _6558};
  wire [2:0] _21745 = {_0, _21743} + {_0, _21744};
  wire [1:0] _21746 = {_0, _8894} + {_0, _10335};
  wire [3:0] _21747 = {_0, _21745} + {_0, _0, _21746};
  wire _21748 = _12301 < _21747;
  wire _21749 = r998 ^ _21748;
  wire _21750 = _12298 ? coded_block[998] : r998;
  wire _21751 = _12296 ? _21749 : _21750;
  always @ (posedge reset or posedge clock) if (reset) r998 <= 1'd0; else if (_12300) r998 <= _21751;
  wire [1:0] _21752 = {_0, _1823} + {_0, _2463};
  wire [1:0] _21753 = {_0, _5757} + {_0, _7773};
  wire [2:0] _21754 = {_0, _21752} + {_0, _21753};
  wire [1:0] _21755 = {_0, _8638} + {_0, _10973};
  wire [3:0] _21756 = {_0, _21754} + {_0, _0, _21755};
  wire _21757 = _12301 < _21756;
  wire _21758 = r997 ^ _21757;
  wire _21759 = _12298 ? coded_block[997] : r997;
  wire _21760 = _12296 ? _21758 : _21759;
  always @ (posedge reset or posedge clock) if (reset) r997 <= 1'd0; else if (_12300) r997 <= _21760;
  wire [1:0] _21761 = {_0, _1854} + {_0, _3167};
  wire [1:0] _21762 = {_0, _4542} + {_0, _7837};
  wire [2:0] _21763 = {_0, _21761} + {_0, _21762};
  wire [1:0] _21764 = {_0, _9853} + {_0, _10717};
  wire [3:0] _21765 = {_0, _21763} + {_0, _0, _21764};
  wire _21766 = _12301 < _21765;
  wire _21767 = r996 ^ _21766;
  wire _21768 = _12298 ? coded_block[996] : r996;
  wire _21769 = _12296 ? _21767 : _21768;
  always @ (posedge reset or posedge clock) if (reset) r996 <= 1'd0; else if (_12300) r996 <= _21769;
  wire [1:0] _21770 = {_0, _1886} + {_0, _3068};
  wire [1:0] _21771 = {_0, _5246} + {_0, _6621};
  wire [2:0] _21772 = {_0, _21770} + {_0, _21771};
  wire [1:0] _21773 = {_0, _9917} + {_0, _11933};
  wire [3:0] _21774 = {_0, _21772} + {_0, _0, _21773};
  wire _21775 = _12301 < _21774;
  wire _21776 = r995 ^ _21775;
  wire _21777 = _12298 ? coded_block[995] : r995;
  wire _21778 = _12296 ? _21776 : _21777;
  always @ (posedge reset or posedge clock) if (reset) r995 <= 1'd0; else if (_12300) r995 <= _21778;
  wire [1:0] _21779 = {_0, _1917} + {_0, _3580};
  wire [1:0] _21780 = {_0, _5152} + {_0, _7326};
  wire [2:0] _21781 = {_0, _21779} + {_0, _21780};
  wire [1:0] _21782 = {_0, _8701} + {_0, _11996};
  wire [3:0] _21783 = {_0, _21781} + {_0, _0, _21782};
  wire _21784 = _12301 < _21783;
  wire _21785 = r994 ^ _21784;
  wire _21786 = _12298 ? coded_block[994] : r994;
  wire _21787 = _12296 ? _21785 : _21786;
  always @ (posedge reset or posedge clock) if (reset) r994 <= 1'd0; else if (_12300) r994 <= _21787;
  wire [1:0] _21788 = {_0, _1950} + {_0, _2430};
  wire [1:0] _21789 = {_0, _5663} + {_0, _7230};
  wire [2:0] _21790 = {_0, _21788} + {_0, _21789};
  wire [1:0] _21791 = {_0, _9406} + {_0, _10783};
  wire [3:0] _21792 = {_0, _21790} + {_0, _0, _21791};
  wire _21793 = _12301 < _21792;
  wire _21794 = r993 ^ _21793;
  wire _21795 = _12298 ? coded_block[993] : r993;
  wire _21796 = _12296 ? _21794 : _21795;
  always @ (posedge reset or posedge clock) if (reset) r993 <= 1'd0; else if (_12300) r993 <= _21796;
  wire [1:0] _21797 = {_0, _1981} + {_0, _3709};
  wire [1:0] _21798 = {_0, _4511} + {_0, _7741};
  wire [2:0] _21799 = {_0, _21797} + {_0, _21798};
  wire [1:0] _21800 = {_0, _9311} + {_0, _11485};
  wire [3:0] _21801 = {_0, _21799} + {_0, _0, _21800};
  wire _21802 = _12301 < _21801;
  wire _21803 = r992 ^ _21802;
  wire _21804 = _12298 ? coded_block[992] : r992;
  wire _21805 = _12296 ? _21803 : _21804;
  always @ (posedge reset or posedge clock) if (reset) r992 <= 1'd0; else if (_12300) r992 <= _21805;
  wire [1:0] _21806 = {_0, _2044} + {_0, _3294};
  wire [1:0] _21807 = {_0, _4830} + {_0, _7868};
  wire [2:0] _21808 = {_0, _21806} + {_0, _21807};
  wire [1:0] _21809 = {_0, _8670} + {_0, _11900};
  wire [3:0] _21810 = {_0, _21808} + {_0, _0, _21809};
  wire _21811 = _12301 < _21810;
  wire _21812 = r991 ^ _21811;
  wire _21813 = _12298 ? coded_block[991] : r991;
  wire _21814 = _12296 ? _21812 : _21813;
  always @ (posedge reset or posedge clock) if (reset) r991 <= 1'd0; else if (_12300) r991 <= _21814;
  wire [1:0] _21815 = {_0, _65} + {_0, _2367};
  wire [1:0] _21816 = {_0, _5373} + {_0, _6908};
  wire [2:0] _21817 = {_0, _21815} + {_0, _21816};
  wire [1:0] _21818 = {_0, _9949} + {_0, _10748};
  wire [3:0] _21819 = {_0, _21817} + {_0, _0, _21818};
  wire _21820 = _12301 < _21819;
  wire _21821 = r990 ^ _21820;
  wire _21822 = _12298 ? coded_block[990] : r990;
  wire _21823 = _12296 ? _21821 : _21822;
  always @ (posedge reset or posedge clock) if (reset) r990 <= 1'd0; else if (_12300) r990 <= _21823;
  wire [1:0] _21824 = {_0, _97} + {_0, _2686};
  wire [1:0] _21825 = {_0, _4447} + {_0, _7454};
  wire [2:0] _21826 = {_0, _21824} + {_0, _21825};
  wire [1:0] _21827 = {_0, _8991} + {_0, _12027};
  wire [3:0] _21828 = {_0, _21826} + {_0, _0, _21827};
  wire _21829 = _12301 < _21828;
  wire _21830 = r989 ^ _21829;
  wire _21831 = _12298 ? coded_block[989] : r989;
  wire _21832 = _12296 ? _21830 : _21831;
  always @ (posedge reset or posedge clock) if (reset) r989 <= 1'd0; else if (_12300) r989 <= _21832;
  wire [1:0] _21833 = {_0, _128} + {_0, _3135};
  wire [1:0] _21834 = {_0, _4767} + {_0, _6525};
  wire [2:0] _21835 = {_0, _21833} + {_0, _21834};
  wire [1:0] _21836 = {_0, _9534} + {_0, _11069};
  wire [3:0] _21837 = {_0, _21835} + {_0, _0, _21836};
  wire _21838 = _12301 < _21837;
  wire _21839 = r988 ^ _21838;
  wire _21840 = _12298 ? coded_block[988] : r988;
  wire _21841 = _12296 ? _21839 : _21840;
  always @ (posedge reset or posedge clock) if (reset) r988 <= 1'd0; else if (_12300) r988 <= _21841;
  wire [1:0] _21842 = {_0, _161} + {_0, _2494};
  wire [1:0] _21843 = {_0, _5215} + {_0, _6845};
  wire [2:0] _21844 = {_0, _21842} + {_0, _21843};
  wire [1:0] _21845 = {_0, _8607} + {_0, _11613};
  wire [3:0] _21846 = {_0, _21844} + {_0, _0, _21845};
  wire _21847 = _12301 < _21846;
  wire _21848 = r987 ^ _21847;
  wire _21849 = _12298 ? coded_block[987] : r987;
  wire _21850 = _12296 ? _21848 : _21849;
  always @ (posedge reset or posedge clock) if (reset) r987 <= 1'd0; else if (_12300) r987 <= _21850;
  wire [1:0] _21851 = {_0, _192} + {_0, _3422};
  wire [1:0] _21852 = {_0, _4574} + {_0, _7293};
  wire [2:0] _21853 = {_0, _21851} + {_0, _21852};
  wire [1:0] _21854 = {_0, _8926} + {_0, _10685};
  wire [3:0] _21855 = {_0, _21853} + {_0, _0, _21854};
  wire _21856 = _12301 < _21855;
  wire _21857 = r986 ^ _21856;
  wire _21858 = _12298 ? coded_block[986] : r986;
  wire _21859 = _12296 ? _21857 : _21858;
  always @ (posedge reset or posedge clock) if (reset) r986 <= 1'd0; else if (_12300) r986 <= _21859;
  wire [1:0] _21860 = {_0, _224} + {_0, _3517};
  wire [1:0] _21861 = {_0, _5501} + {_0, _6652};
  wire [2:0] _21862 = {_0, _21860} + {_0, _21861};
  wire [1:0] _21863 = {_0, _9375} + {_0, _11004};
  wire [3:0] _21864 = {_0, _21862} + {_0, _0, _21863};
  wire _21865 = _12301 < _21864;
  wire _21866 = r985 ^ _21865;
  wire _21867 = _12298 ? coded_block[985] : r985;
  wire _21868 = _12296 ? _21866 : _21867;
  always @ (posedge reset or posedge clock) if (reset) r985 <= 1'd0; else if (_12300) r985 <= _21868;
  wire [1:0] _21869 = {_0, _255} + {_0, _2974};
  wire [1:0] _21870 = {_0, _5597} + {_0, _7581};
  wire [2:0] _21871 = {_0, _21869} + {_0, _21870};
  wire [1:0] _21872 = {_0, _8736} + {_0, _11453};
  wire [3:0] _21873 = {_0, _21871} + {_0, _0, _21872};
  wire _21874 = _12301 < _21873;
  wire _21875 = r984 ^ _21874;
  wire _21876 = _12298 ? coded_block[984] : r984;
  wire _21877 = _12296 ? _21875 : _21876;
  always @ (posedge reset or posedge clock) if (reset) r984 <= 1'd0; else if (_12300) r984 <= _21877;
  wire [1:0] _21878 = {_0, _289} + {_0, _3231};
  wire [1:0] _21879 = {_0, _5053} + {_0, _7675};
  wire [2:0] _21880 = {_0, _21878} + {_0, _21879};
  wire [1:0] _21881 = {_0, _9661} + {_0, _10814};
  wire [3:0] _21882 = {_0, _21880} + {_0, _0, _21881};
  wire _21883 = _12301 < _21882;
  wire _21884 = r983 ^ _21883;
  wire _21885 = _12298 ? coded_block[983] : r983;
  wire _21886 = _12296 ? _21884 : _21885;
  always @ (posedge reset or posedge clock) if (reset) r983 <= 1'd0; else if (_12300) r983 <= _21886;
  wire [1:0] _21887 = {_0, _320} + {_0, _2112};
  wire [1:0] _21888 = {_0, _5310} + {_0, _7132};
  wire [2:0] _21889 = {_0, _21887} + {_0, _21888};
  wire [1:0] _21890 = {_0, _9759} + {_0, _11740};
  wire [3:0] _21891 = {_0, _21889} + {_0, _0, _21890};
  wire _21892 = _12301 < _21891;
  wire _21893 = r982 ^ _21892;
  wire _21894 = _12298 ? coded_block[982] : r982;
  wire _21895 = _12296 ? _21893 : _21894;
  always @ (posedge reset or posedge clock) if (reset) r982 <= 1'd0; else if (_12300) r982 <= _21895;
  wire [1:0] _21896 = {_0, _352} + {_0, _3773};
  wire [1:0] _21897 = {_0, _4192} + {_0, _7389};
  wire [2:0] _21898 = {_0, _21896} + {_0, _21897};
  wire [1:0] _21899 = {_0, _9212} + {_0, _11837};
  wire [3:0] _21900 = {_0, _21898} + {_0, _0, _21899};
  wire _21901 = _12301 < _21900;
  wire _21902 = r981 ^ _21901;
  wire _21903 = _12298 ? coded_block[981] : r981;
  wire _21904 = _12296 ? _21902 : _21903;
  always @ (posedge reset or posedge clock) if (reset) r981 <= 1'd0; else if (_12300) r981 <= _21904;
  wire [1:0] _21905 = {_0, _416} + {_0, _3870};
  wire [1:0] _21906 = {_0, _6076} + {_0, _7931};
  wire [2:0] _21907 = {_0, _21905} + {_0, _21906};
  wire [1:0] _21908 = {_0, _8352} + {_0, _11550};
  wire [3:0] _21909 = {_0, _21907} + {_0, _0, _21908};
  wire _21910 = _12301 < _21909;
  wire _21911 = r980 ^ _21910;
  wire _21912 = _12298 ? coded_block[980] : r980;
  wire _21913 = _12296 ? _21911 : _21912;
  always @ (posedge reset or posedge clock) if (reset) r980 <= 1'd0; else if (_12300) r980 <= _21913;
  wire [1:0] _21914 = {_0, _447} + {_0, _2208};
  wire [1:0] _21915 = {_0, _5949} + {_0, _8155};
  wire [2:0] _21916 = {_0, _21914} + {_0, _21915};
  wire [1:0] _21917 = {_0, _10014} + {_0, _10430};
  wire [3:0] _21918 = {_0, _21916} + {_0, _0, _21917};
  wire _21919 = _12301 < _21918;
  wire _21920 = r979 ^ _21919;
  wire _21921 = _12298 ? coded_block[979] : r979;
  wire _21922 = _12296 ? _21920 : _21921;
  always @ (posedge reset or posedge clock) if (reset) r979 <= 1'd0; else if (_12300) r979 <= _21922;
  wire [1:0] _21923 = {_0, _479} + {_0, _2941};
  wire [1:0] _21924 = {_0, _4287} + {_0, _8028};
  wire [2:0] _21925 = {_0, _21923} + {_0, _21924};
  wire [1:0] _21926 = {_0, _10235} + {_0, _12092};
  wire [3:0] _21927 = {_0, _21925} + {_0, _0, _21926};
  wire _21928 = _12301 < _21927;
  wire _21929 = r978 ^ _21928;
  wire _21930 = _12298 ? coded_block[978] : r978;
  wire _21931 = _12296 ? _21929 : _21930;
  always @ (posedge reset or posedge clock) if (reset) r978 <= 1'd0; else if (_12300) r978 <= _21931;
  wire [1:0] _21932 = {_0, _510} + {_0, _3549};
  wire [1:0] _21933 = {_0, _5022} + {_0, _6366};
  wire [2:0] _21934 = {_0, _21932} + {_0, _21933};
  wire [1:0] _21935 = {_0, _10108} + {_0, _10303};
  wire [3:0] _21936 = {_0, _21934} + {_0, _0, _21935};
  wire _21937 = _12301 < _21936;
  wire _21938 = r977 ^ _21937;
  wire _21939 = _12298 ? coded_block[977] : r977;
  wire _21940 = _12296 ? _21938 : _21939;
  always @ (posedge reset or posedge clock) if (reset) r977 <= 1'd0; else if (_12300) r977 <= _21940;
  wire [1:0] _21941 = {_0, _545} + {_0, _3104};
  wire [1:0] _21942 = {_0, _5628} + {_0, _7100};
  wire [2:0] _21943 = {_0, _21941} + {_0, _21942};
  wire [1:0] _21944 = {_0, _8446} + {_0, _12188};
  wire [3:0] _21945 = {_0, _21943} + {_0, _0, _21944};
  wire _21946 = _12301 < _21945;
  wire _21947 = r976 ^ _21946;
  wire _21948 = _12298 ? coded_block[976] : r976;
  wire _21949 = _12296 ? _21947 : _21948;
  always @ (posedge reset or posedge clock) if (reset) r976 <= 1'd0; else if (_12300) r976 <= _21949;
  wire [1:0] _21950 = {_0, _576} + {_0, _2719};
  wire [1:0] _21951 = {_0, _5183} + {_0, _7710};
  wire [2:0] _21952 = {_0, _21950} + {_0, _21951};
  wire [1:0] _21953 = {_0, _9181} + {_0, _10527};
  wire [3:0] _21954 = {_0, _21952} + {_0, _0, _21953};
  wire _21955 = _12301 < _21954;
  wire _21956 = r975 ^ _21955;
  wire _21957 = _12298 ? coded_block[975] : r975;
  wire _21958 = _12296 ? _21956 : _21957;
  always @ (posedge reset or posedge clock) if (reset) r975 <= 1'd0; else if (_12300) r975 <= _21958;
  wire [1:0] _21959 = {_0, _608} + {_0, _3742};
  wire [1:0] _21960 = {_0, _4798} + {_0, _7262};
  wire [2:0] _21961 = {_0, _21959} + {_0, _21960};
  wire [1:0] _21962 = {_0, _9790} + {_0, _11259};
  wire [3:0] _21963 = {_0, _21961} + {_0, _0, _21962};
  wire _21964 = _12301 < _21963;
  wire _21965 = r974 ^ _21964;
  wire _21966 = _12298 ? coded_block[974] : r974;
  wire _21967 = _12296 ? _21965 : _21966;
  always @ (posedge reset or posedge clock) if (reset) r974 <= 1'd0; else if (_12300) r974 <= _21967;
  wire [1:0] _21968 = {_0, _639} + {_0, _2144};
  wire [1:0] _21969 = {_0, _5821} + {_0, _6877};
  wire [2:0] _21970 = {_0, _21968} + {_0, _21969};
  wire [1:0] _21971 = {_0, _9342} + {_0, _11869};
  wire [3:0] _21972 = {_0, _21970} + {_0, _0, _21971};
  wire _21973 = _12301 < _21972;
  wire _21974 = r973 ^ _21973;
  wire _21975 = _12298 ? coded_block[973] : r973;
  wire _21976 = _12296 ? _21974 : _21975;
  always @ (posedge reset or posedge clock) if (reset) r973 <= 1'd0; else if (_12300) r973 <= _21976;
  wire [1:0] _21977 = {_0, _672} + {_0, _2623};
  wire [1:0] _21978 = {_0, _4223} + {_0, _7900};
  wire [2:0] _21979 = {_0, _21977} + {_0, _21978};
  wire [1:0] _21980 = {_0, _8957} + {_0, _11422};
  wire [3:0] _21981 = {_0, _21979} + {_0, _0, _21980};
  wire _21982 = _12301 < _21981;
  wire _21983 = r972 ^ _21982;
  wire _21984 = _12298 ? coded_block[972] : r972;
  wire _21985 = _12296 ? _21983 : _21984;
  always @ (posedge reset or posedge clock) if (reset) r972 <= 1'd0; else if (_12300) r972 <= _21985;
  wire [1:0] _21986 = {_0, _703} + {_0, _4060};
  wire [1:0] _21987 = {_0, _4703} + {_0, _6303};
  wire [2:0] _21988 = {_0, _21986} + {_0, _21987};
  wire [1:0] _21989 = {_0, _9980} + {_0, _11038};
  wire [3:0] _21990 = {_0, _21988} + {_0, _0, _21989};
  wire _21991 = _12301 < _21990;
  wire _21992 = r971 ^ _21991;
  wire _21993 = _12298 ? coded_block[971] : r971;
  wire _21994 = _12296 ? _21992 : _21993;
  always @ (posedge reset or posedge clock) if (reset) r971 <= 1'd0; else if (_12300) r971 <= _21994;
  wire [1:0] _21995 = {_0, _735} + {_0, _3359};
  wire [1:0] _21996 = {_0, _6139} + {_0, _6781};
  wire [2:0] _21997 = {_0, _21995} + {_0, _21996};
  wire [1:0] _21998 = {_0, _8383} + {_0, _12061};
  wire [3:0] _21999 = {_0, _21997} + {_0, _0, _21998};
  wire _22000 = _12301 < _21999;
  wire _22001 = r970 ^ _22000;
  wire _22002 = _12298 ? coded_block[970] : r970;
  wire _22003 = _12296 ? _22001 : _22002;
  always @ (posedge reset or posedge clock) if (reset) r970 <= 1'd0; else if (_12300) r970 <= _22003;
  wire [1:0] _22004 = {_0, _766} + {_0, _3037};
  wire [1:0] _22005 = {_0, _5438} + {_0, _6207};
  wire [2:0] _22006 = {_0, _22004} + {_0, _22005};
  wire [1:0] _22007 = {_0, _8863} + {_0, _10462};
  wire [3:0] _22008 = {_0, _22006} + {_0, _0, _22007};
  wire _22009 = _12301 < _22008;
  wire _22010 = r969 ^ _22009;
  wire _22011 = _12298 ? coded_block[969] : r969;
  wire _22012 = _12296 ? _22010 : _22011;
  always @ (posedge reset or posedge clock) if (reset) r969 <= 1'd0; else if (_12300) r969 <= _22012;
  wire [1:0] _22013 = {_0, _800} + {_0, _3198};
  wire [1:0] _22014 = {_0, _5116} + {_0, _7517};
  wire [2:0] _22015 = {_0, _22013} + {_0, _22014};
  wire [1:0] _22016 = {_0, _8288} + {_0, _10941};
  wire [3:0] _22017 = {_0, _22015} + {_0, _0, _22016};
  wire _22018 = _12301 < _22017;
  wire _22019 = r968 ^ _22018;
  wire _22020 = _12298 ? coded_block[968] : r968;
  wire _22021 = _12296 ? _22019 : _22020;
  always @ (posedge reset or posedge clock) if (reset) r968 <= 1'd0; else if (_12300) r968 <= _22021;
  wire [1:0] _22022 = {_0, _831} + {_0, _3005};
  wire [1:0] _22023 = {_0, _5279} + {_0, _7199};
  wire [2:0] _22024 = {_0, _22022} + {_0, _22023};
  wire [1:0] _22025 = {_0, _9597} + {_0, _10366};
  wire [3:0] _22026 = {_0, _22024} + {_0, _0, _22025};
  wire _22027 = _12301 < _22026;
  wire _22028 = r967 ^ _22027;
  wire _22029 = _12298 ? coded_block[967] : r967;
  wire _22030 = _12296 ? _22028 : _22029;
  always @ (posedge reset or posedge clock) if (reset) r967 <= 1'd0; else if (_12300) r967 <= _22030;
  wire [1:0] _22031 = {_0, _863} + {_0, _3390};
  wire [1:0] _22032 = {_0, _5085} + {_0, _7357};
  wire [2:0] _22033 = {_0, _22031} + {_0, _22032};
  wire [1:0] _22034 = {_0, _9279} + {_0, _11677};
  wire [3:0] _22035 = {_0, _22033} + {_0, _0, _22034};
  wire _22036 = _12301 < _22035;
  wire _22037 = r966 ^ _22036;
  wire _22038 = _12298 ? coded_block[966] : r966;
  wire _22039 = _12296 ? _22037 : _22038;
  always @ (posedge reset or posedge clock) if (reset) r966 <= 1'd0; else if (_12300) r966 <= _22039;
  wire [1:0] _22040 = {_0, _894} + {_0, _2526};
  wire [1:0] _22041 = {_0, _5470} + {_0, _7163};
  wire [2:0] _22042 = {_0, _22040} + {_0, _22041};
  wire [1:0] _22043 = {_0, _9438} + {_0, _11358};
  wire [3:0] _22044 = {_0, _22042} + {_0, _0, _22043};
  wire _22045 = _12301 < _22044;
  wire _22046 = r965 ^ _22045;
  wire _22047 = _12298 ? coded_block[965] : r965;
  wire _22048 = _12296 ? _22046 : _22047;
  always @ (posedge reset or posedge clock) if (reset) r965 <= 1'd0; else if (_12300) r965 <= _22048;
  wire [1:0] _22049 = {_0, _927} + {_0, _2302};
  wire [1:0] _22050 = {_0, _4605} + {_0, _7548};
  wire [2:0] _22051 = {_0, _22049} + {_0, _22050};
  wire [1:0] _22052 = {_0, _9248} + {_0, _11516};
  wire [3:0] _22053 = {_0, _22051} + {_0, _0, _22052};
  wire _22054 = _12301 < _22053;
  wire _22055 = r964 ^ _22054;
  wire _22056 = _12298 ? coded_block[964] : r964;
  wire _22057 = _12296 ? _22055 : _22056;
  always @ (posedge reset or posedge clock) if (reset) r964 <= 1'd0; else if (_12300) r964 <= _22057;
  wire [1:0] _22058 = {_0, _990} + {_0, _2813};
  wire [1:0] _22059 = {_0, _4958} + {_0, _6462};
  wire [2:0] _22060 = {_0, _22058} + {_0, _22059};
  wire [1:0] _22061 = {_0, _8767} + {_0, _11708};
  wire [3:0] _22062 = {_0, _22060} + {_0, _0, _22061};
  wire _22063 = _12301 < _22062;
  wire _22064 = r963 ^ _22063;
  wire _22065 = _12298 ? coded_block[963] : r963;
  wire _22066 = _12296 ? _22064 : _22065;
  always @ (posedge reset or posedge clock) if (reset) r963 <= 1'd0; else if (_12300) r963 <= _22066;
  wire [1:0] _22067 = {_0, _1021} + {_0, _3933};
  wire [1:0] _22068 = {_0, _4895} + {_0, _7036};
  wire [2:0] _22069 = {_0, _22067} + {_0, _22068};
  wire [1:0] _22070 = {_0, _8543} + {_0, _10846};
  wire [3:0] _22071 = {_0, _22069} + {_0, _0, _22070};
  wire _22072 = _12301 < _22071;
  wire _22073 = r962 ^ _22072;
  wire _22074 = _12298 ? coded_block[962] : r962;
  wire _22075 = _12296 ? _22073 : _22074;
  always @ (posedge reset or posedge clock) if (reset) r962 <= 1'd0; else if (_12300) r962 <= _22075;
  wire [1:0] _22076 = {_0, _1057} + {_0, _2592};
  wire [1:0] _22077 = {_0, _6012} + {_0, _6973};
  wire [2:0] _22078 = {_0, _22076} + {_0, _22077};
  wire [1:0] _22079 = {_0, _9118} + {_0, _10621};
  wire [3:0] _22080 = {_0, _22078} + {_0, _0, _22079};
  wire _22081 = _12301 < _22080;
  wire _22082 = r961 ^ _22081;
  wire _22083 = _12298 ? coded_block[961] : r961;
  wire _22084 = _12296 ? _22082 : _22083;
  always @ (posedge reset or posedge clock) if (reset) r961 <= 1'd0; else if (_12300) r961 <= _22084;
  wire [1:0] _22085 = {_0, _1088} + {_0, _2175};
  wire [1:0] _22086 = {_0, _4671} + {_0, _8092};
  wire [2:0] _22087 = {_0, _22085} + {_0, _22086};
  wire [1:0] _22088 = {_0, _9054} + {_0, _11196};
  wire [3:0] _22089 = {_0, _22087} + {_0, _0, _22088};
  wire _22090 = _12301 < _22089;
  wire _22091 = r960 ^ _22090;
  wire _22092 = _12298 ? coded_block[960] : r960;
  wire _22093 = _12296 ? _22091 : _22092;
  always @ (posedge reset or posedge clock) if (reset) r960 <= 1'd0; else if (_12300) r960 <= _22093;
  wire [1:0] _22094 = {_0, _1120} + {_0, _3901};
  wire [1:0] _22095 = {_0, _4256} + {_0, _6750};
  wire [2:0] _22096 = {_0, _22094} + {_0, _22095};
  wire [1:0] _22097 = {_0, _10172} + {_0, _11132};
  wire [3:0] _22098 = {_0, _22096} + {_0, _0, _22097};
  wire _22099 = _12301 < _22098;
  wire _22100 = r959 ^ _22099;
  wire _22101 = _12298 ? coded_block[959] : r959;
  wire _22102 = _12296 ? _22100 : _22101;
  always @ (posedge reset or posedge clock) if (reset) r959 <= 1'd0; else if (_12300) r959 <= _22102;
  wire [1:0] _22103 = {_0, _1151} + {_0, _2847};
  wire [1:0] _22104 = {_0, _5981} + {_0, _6334};
  wire [2:0] _22105 = {_0, _22103} + {_0, _22104};
  wire [1:0] _22106 = {_0, _8830} + {_0, _12251};
  wire [3:0] _22107 = {_0, _22105} + {_0, _0, _22106};
  wire _22108 = _12301 < _22107;
  wire _22109 = r958 ^ _22108;
  wire _22110 = _12298 ? coded_block[958] : r958;
  wire _22111 = _12296 ? _22109 : _22110;
  always @ (posedge reset or posedge clock) if (reset) r958 <= 1'd0; else if (_12300) r958 <= _22111;
  wire [1:0] _22112 = {_0, _1184} + {_0, _2336};
  wire [1:0] _22113 = {_0, _4926} + {_0, _8059};
  wire [2:0] _22114 = {_0, _22112} + {_0, _22113};
  wire [1:0] _22115 = {_0, _8415} + {_0, _10910};
  wire [3:0] _22116 = {_0, _22114} + {_0, _0, _22115};
  wire _22117 = _12301 < _22116;
  wire _22118 = r957 ^ _22117;
  wire _22119 = _12298 ? coded_block[957] : r957;
  wire _22120 = _12296 ? _22118 : _22119;
  always @ (posedge reset or posedge clock) if (reset) r957 <= 1'd0; else if (_12300) r957 <= _22120;
  wire [1:0] _22121 = {_0, _1215} + {_0, _3325};
  wire [1:0] _22122 = {_0, _4415} + {_0, _7005};
  wire [2:0] _22123 = {_0, _22121} + {_0, _22122};
  wire [1:0] _22124 = {_0, _10141} + {_0, _10493};
  wire [3:0] _22125 = {_0, _22123} + {_0, _0, _22124};
  wire _22126 = _12301 < _22125;
  wire _22127 = r956 ^ _22126;
  wire _22128 = _12298 ? coded_block[956] : r956;
  wire _22129 = _12296 ? _22127 : _22128;
  always @ (posedge reset or posedge clock) if (reset) r956 <= 1'd0; else if (_12300) r956 <= _22129;
  wire [1:0] _22130 = {_0, _1247} + {_0, _4091};
  wire [1:0] _22131 = {_0, _5407} + {_0, _6494};
  wire [2:0] _22132 = {_0, _22130} + {_0, _22131};
  wire [1:0] _22133 = {_0, _9085} + {_0, _12219};
  wire [3:0] _22134 = {_0, _22132} + {_0, _0, _22133};
  wire _22135 = _12301 < _22134;
  wire _22136 = r955 ^ _22135;
  wire _22137 = _12298 ? coded_block[955] : r955;
  wire _22138 = _12296 ? _22136 : _22137;
  always @ (posedge reset or posedge clock) if (reset) r955 <= 1'd0; else if (_12300) r955 <= _22138;
  wire [1:0] _22139 = {_0, _1278} + {_0, _3262};
  wire [1:0] _22140 = {_0, _4160} + {_0, _7485};
  wire [2:0] _22141 = {_0, _22139} + {_0, _22140};
  wire [1:0] _22142 = {_0, _8574} + {_0, _11165};
  wire [3:0] _22143 = {_0, _22141} + {_0, _0, _22142};
  wire _22144 = _12301 < _22143;
  wire _22145 = r954 ^ _22144;
  wire _22146 = _12298 ? coded_block[954] : r954;
  wire _22147 = _12296 ? _22145 : _22146;
  always @ (posedge reset or posedge clock) if (reset) r954 <= 1'd0; else if (_12300) r954 <= _22147;
  wire [1:0] _22148 = {_0, _1312} + {_0, _2782};
  wire [1:0] _22149 = {_0, _5342} + {_0, _6239};
  wire [2:0] _22150 = {_0, _22148} + {_0, _22149};
  wire [1:0] _22151 = {_0, _9566} + {_0, _10654};
  wire [3:0] _22152 = {_0, _22150} + {_0, _0, _22151};
  wire _22153 = _12301 < _22152;
  wire _22154 = r953 ^ _22153;
  wire _22155 = _12298 ? coded_block[953] : r953;
  wire _22156 = _12296 ? _22154 : _22155;
  always @ (posedge reset or posedge clock) if (reset) r953 <= 1'd0; else if (_12300) r953 <= _22156;
  wire [1:0] _22157 = {_0, _1343} + {_0, _2910};
  wire [1:0] _22158 = {_0, _4861} + {_0, _7420};
  wire [2:0] _22159 = {_0, _22157} + {_0, _22158};
  wire [1:0] _22160 = {_0, _8319} + {_0, _11644};
  wire [3:0] _22161 = {_0, _22159} + {_0, _0, _22160};
  wire _22162 = _12301 < _22161;
  wire _22163 = r952 ^ _22162;
  wire _22164 = _12298 ? coded_block[952] : r952;
  wire _22165 = _12296 ? _22163 : _22164;
  always @ (posedge reset or posedge clock) if (reset) r952 <= 1'd0; else if (_12300) r952 <= _22165;
  wire [1:0] _22166 = {_0, _1375} + {_0, _2239};
  wire [1:0] _22167 = {_0, _4989} + {_0, _6942};
  wire [2:0] _22168 = {_0, _22166} + {_0, _22167};
  wire [1:0] _22169 = {_0, _9503} + {_0, _10399};
  wire [3:0] _22170 = {_0, _22168} + {_0, _0, _22169};
  wire _22171 = _12301 < _22170;
  wire _22172 = r951 ^ _22171;
  wire _22173 = _12298 ? coded_block[951] : r951;
  wire _22174 = _12296 ? _22172 : _22173;
  always @ (posedge reset or posedge clock) if (reset) r951 <= 1'd0; else if (_12300) r951 <= _22174;
  wire [1:0] _22175 = {_0, _1406} + {_0, _3486};
  wire [1:0] _22176 = {_0, _4319} + {_0, _7069};
  wire [2:0] _22177 = {_0, _22175} + {_0, _22176};
  wire [1:0] _22178 = {_0, _9022} + {_0, _11581};
  wire [3:0] _22179 = {_0, _22177} + {_0, _0, _22178};
  wire _22180 = _12301 < _22179;
  wire _22181 = r950 ^ _22180;
  wire _22182 = _12298 ? coded_block[950] : r950;
  wire _22183 = _12296 ? _22181 : _22182;
  always @ (posedge reset or posedge clock) if (reset) r950 <= 1'd0; else if (_12300) r950 <= _22183;
  wire [1:0] _22184 = {_0, _1439} + {_0, _3453};
  wire [1:0] _22185 = {_0, _5565} + {_0, _6397};
  wire [2:0] _22186 = {_0, _22184} + {_0, _22185};
  wire [1:0] _22187 = {_0, _9149} + {_0, _11101};
  wire [3:0] _22188 = {_0, _22186} + {_0, _0, _22187};
  wire _22189 = _12301 < _22188;
  wire _22190 = r949 ^ _22189;
  wire _22191 = _12298 ? coded_block[949] : r949;
  wire _22192 = _12296 ? _22190 : _22191;
  always @ (posedge reset or posedge clock) if (reset) r949 <= 1'd0; else if (_12300) r949 <= _22192;
  wire [1:0] _22193 = {_0, _1470} + {_0, _2271};
  wire [1:0] _22194 = {_0, _5534} + {_0, _7644};
  wire [2:0] _22195 = {_0, _22193} + {_0, _22194};
  wire [1:0] _22196 = {_0, _8480} + {_0, _11228};
  wire [3:0] _22197 = {_0, _22195} + {_0, _0, _22196};
  wire _22198 = _12301 < _22197;
  wire _22199 = r948 ^ _22198;
  wire _22200 = _12298 ? coded_block[948] : r948;
  wire _22201 = _12296 ? _22199 : _22200;
  always @ (posedge reset or posedge clock) if (reset) r948 <= 1'd0; else if (_12300) r948 <= _22201;
  wire [1:0] _22202 = {_0, _1502} + {_0, _2557};
  wire [1:0] _22203 = {_0, _4350} + {_0, _7612};
  wire [2:0] _22204 = {_0, _22202} + {_0, _22203};
  wire [1:0] _22205 = {_0, _9724} + {_0, _10558};
  wire [3:0] _22206 = {_0, _22204} + {_0, _0, _22205};
  wire _22207 = _12301 < _22206;
  wire _22208 = r947 ^ _22207;
  wire _22209 = _12298 ? coded_block[947] : r947;
  wire _22210 = _12296 ? _22208 : _22209;
  always @ (posedge reset or posedge clock) if (reset) r947 <= 1'd0; else if (_12300) r947 <= _22210;
  wire [1:0] _22211 = {_0, _1533} + {_0, _3964};
  wire [1:0] _22212 = {_0, _4640} + {_0, _6431};
  wire [2:0] _22213 = {_0, _22211} + {_0, _22212};
  wire [1:0] _22214 = {_0, _9693} + {_0, _11806};
  wire [3:0] _22215 = {_0, _22213} + {_0, _0, _22214};
  wire _22216 = _12301 < _22215;
  wire _22217 = r946 ^ _22216;
  wire _22218 = _12298 ? coded_block[946] : r946;
  wire _22219 = _12296 ? _22217 : _22218;
  always @ (posedge reset or posedge clock) if (reset) r946 <= 1'd0; else if (_12300) r946 <= _22219;
  wire [1:0] _22220 = {_0, _1568} + {_0, _3805};
  wire [1:0] _22221 = {_0, _6045} + {_0, _6718};
  wire [2:0] _22222 = {_0, _22220} + {_0, _22221};
  wire [1:0] _22223 = {_0, _8511} + {_0, _11771};
  wire [3:0] _22224 = {_0, _22222} + {_0, _0, _22223};
  wire _22225 = _12301 < _22224;
  wire _22226 = r945 ^ _22225;
  wire _22227 = _12298 ? coded_block[945] : r945;
  wire _22228 = _12296 ? _22226 : _22227;
  always @ (posedge reset or posedge clock) if (reset) r945 <= 1'd0; else if (_12300) r945 <= _22228;
  wire [1:0] _22229 = {_0, _1599} + {_0, _2081};
  wire [1:0] _22230 = {_0, _5884} + {_0, _8123};
  wire [2:0] _22231 = {_0, _22229} + {_0, _22230};
  wire [1:0] _22232 = {_0, _8799} + {_0, _10590};
  wire [3:0] _22233 = {_0, _22231} + {_0, _0, _22232};
  wire _22234 = _12301 < _22233;
  wire _22235 = r944 ^ _22234;
  wire _22236 = _12298 ? coded_block[944] : r944;
  wire _22237 = _12296 ? _22235 : _22236;
  always @ (posedge reset or posedge clock) if (reset) r944 <= 1'd0; else if (_12300) r944 <= _22237;
  wire [1:0] _22238 = {_0, _1470} + {_0, _2112};
  wire [1:0] _22239 = {_0, _5407} + {_0, _7420};
  wire [2:0] _22240 = {_0, _22238} + {_0, _22239};
  wire [1:0] _22241 = {_0, _8288} + {_0, _10621};
  wire [3:0] _22242 = {_0, _22240} + {_0, _0, _22241};
  wire _22243 = _12301 < _22242;
  wire _22244 = r943 ^ _22243;
  wire _22245 = _12298 ? coded_block[943] : r943;
  wire _22246 = _12296 ? _22244 : _22245;
  always @ (posedge reset or posedge clock) if (reset) r943 <= 1'd0; else if (_12300) r943 <= _22246;
  wire [1:0] _22247 = {_0, _1533} + {_0, _2719};
  wire [1:0] _22248 = {_0, _4895} + {_0, _6270};
  wire [2:0] _22249 = {_0, _22247} + {_0, _22248};
  wire [1:0] _22250 = {_0, _9566} + {_0, _11581};
  wire [3:0] _22251 = {_0, _22249} + {_0, _0, _22250};
  wire _22252 = _12301 < _22251;
  wire _22253 = r942 ^ _22252;
  wire _22254 = _12298 ? coded_block[942] : r942;
  wire _22255 = _12296 ? _22253 : _22254;
  always @ (posedge reset or posedge clock) if (reset) r942 <= 1'd0; else if (_12300) r942 <= _22255;
  wire [1:0] _22256 = {_0, _1568} + {_0, _3231};
  wire [1:0] _22257 = {_0, _4798} + {_0, _6973};
  wire [2:0] _22258 = {_0, _22256} + {_0, _22257};
  wire [1:0] _22259 = {_0, _8352} + {_0, _11644};
  wire [3:0] _22260 = {_0, _22258} + {_0, _0, _22259};
  wire _22261 = _12301 < _22260;
  wire _22262 = r941 ^ _22261;
  wire _22263 = _12298 ? coded_block[941] : r941;
  wire _22264 = _12296 ? _22262 : _22263;
  always @ (posedge reset or posedge clock) if (reset) r941 <= 1'd0; else if (_12300) r941 <= _22264;
  wire [1:0] _22265 = {_0, _1599} + {_0, _4091};
  wire [1:0] _22266 = {_0, _5310} + {_0, _6877};
  wire [2:0] _22267 = {_0, _22265} + {_0, _22266};
  wire [1:0] _22268 = {_0, _9054} + {_0, _10430};
  wire [3:0] _22269 = {_0, _22267} + {_0, _0, _22268};
  wire _22270 = _12301 < _22269;
  wire _22271 = r940 ^ _22270;
  wire _22272 = _12298 ? coded_block[940] : r940;
  wire _22273 = _12296 ? _22271 : _22272;
  always @ (posedge reset or posedge clock) if (reset) r940 <= 1'd0; else if (_12300) r940 <= _22273;
  wire [1:0] _22274 = {_0, _1631} + {_0, _3359};
  wire [1:0] _22275 = {_0, _4160} + {_0, _7389};
  wire [2:0] _22276 = {_0, _22274} + {_0, _22275};
  wire [1:0] _22277 = {_0, _8957} + {_0, _11132};
  wire [3:0] _22278 = {_0, _22276} + {_0, _0, _22277};
  wire _22279 = _12301 < _22278;
  wire _22280 = r939 ^ _22279;
  wire _22281 = _12298 ? coded_block[939] : r939;
  wire _22282 = _12296 ? _22280 : _22281;
  always @ (posedge reset or posedge clock) if (reset) r939 <= 1'd0; else if (_12300) r939 <= _22282;
  wire [1:0] _22283 = {_0, _1662} + {_0, _2399};
  wire [1:0] _22284 = {_0, _5438} + {_0, _6239};
  wire [2:0] _22285 = {_0, _22283} + {_0, _22284};
  wire [1:0] _22286 = {_0, _9469} + {_0, _11038};
  wire [3:0] _22287 = {_0, _22285} + {_0, _0, _22286};
  wire _22288 = _12301 < _22287;
  wire _22289 = r938 ^ _22288;
  wire _22290 = _12298 ? coded_block[938] : r938;
  wire _22291 = _12296 ? _22289 : _22290;
  always @ (posedge reset or posedge clock) if (reset) r938 <= 1'd0; else if (_12300) r938 <= _22291;
  wire [1:0] _22292 = {_0, _1695} + {_0, _2941};
  wire [1:0] _22293 = {_0, _4478} + {_0, _7517};
  wire [2:0] _22294 = {_0, _22292} + {_0, _22293};
  wire [1:0] _22295 = {_0, _8319} + {_0, _11550};
  wire [3:0] _22296 = {_0, _22294} + {_0, _0, _22295};
  wire _22297 = _12301 < _22296;
  wire _22298 = r937 ^ _22297;
  wire _22299 = _12298 ? coded_block[937] : r937;
  wire _22300 = _12296 ? _22298 : _22299;
  always @ (posedge reset or posedge clock) if (reset) r937 <= 1'd0; else if (_12300) r937 <= _22300;
  wire [1:0] _22301 = {_0, _1726} + {_0, _4028};
  wire [1:0] _22302 = {_0, _5022} + {_0, _6558};
  wire [2:0] _22303 = {_0, _22301} + {_0, _22302};
  wire [1:0] _22304 = {_0, _9597} + {_0, _10399};
  wire [3:0] _22305 = {_0, _22303} + {_0, _0, _22304};
  wire _22306 = _12301 < _22305;
  wire _22307 = r936 ^ _22306;
  wire _22308 = _12298 ? coded_block[936] : r936;
  wire _22309 = _12296 ? _22307 : _22308;
  always @ (posedge reset or posedge clock) if (reset) r936 <= 1'd0; else if (_12300) r936 <= _22309;
  wire [1:0] _22310 = {_0, _1758} + {_0, _2336};
  wire [1:0] _22311 = {_0, _6108} + {_0, _7100};
  wire [2:0] _22312 = {_0, _22310} + {_0, _22311};
  wire [1:0] _22313 = {_0, _8638} + {_0, _11677};
  wire [3:0] _22314 = {_0, _22312} + {_0, _0, _22313};
  wire _22315 = _12301 < _22314;
  wire _22316 = r935 ^ _22315;
  wire _22317 = _12298 ? coded_block[935] : r935;
  wire _22318 = _12296 ? _22316 : _22317;
  always @ (posedge reset or posedge clock) if (reset) r935 <= 1'd0; else if (_12300) r935 <= _22318;
  wire [1:0] _22319 = {_0, _1789} + {_0, _2782};
  wire [1:0] _22320 = {_0, _4415} + {_0, _8186};
  wire [2:0] _22321 = {_0, _22319} + {_0, _22320};
  wire [1:0] _22322 = {_0, _9181} + {_0, _10717};
  wire [3:0] _22323 = {_0, _22321} + {_0, _0, _22322};
  wire _22324 = _12301 < _22323;
  wire _22325 = r934 ^ _22324;
  wire _22326 = _12298 ? coded_block[934] : r934;
  wire _22327 = _12296 ? _22325 : _22326;
  always @ (posedge reset or posedge clock) if (reset) r934 <= 1'd0; else if (_12300) r934 <= _22327;
  wire [1:0] _22328 = {_0, _1823} + {_0, _2144};
  wire [1:0] _22329 = {_0, _4861} + {_0, _6494};
  wire [2:0] _22330 = {_0, _22328} + {_0, _22329};
  wire [1:0] _22331 = {_0, _8256} + {_0, _11259};
  wire [3:0] _22332 = {_0, _22330} + {_0, _0, _22331};
  wire _22333 = _12301 < _22332;
  wire _22334 = r933 ^ _22333;
  wire _22335 = _12298 ? coded_block[933] : r933;
  wire _22336 = _12296 ? _22334 : _22335;
  always @ (posedge reset or posedge clock) if (reset) r933 <= 1'd0; else if (_12300) r933 <= _22336;
  wire [1:0] _22337 = {_0, _1854} + {_0, _3068};
  wire [1:0] _22338 = {_0, _4223} + {_0, _6942};
  wire [2:0] _22339 = {_0, _22337} + {_0, _22338};
  wire [1:0] _22340 = {_0, _8574} + {_0, _10335};
  wire [3:0] _22341 = {_0, _22339} + {_0, _0, _22340};
  wire _22342 = _12301 < _22341;
  wire _22343 = r932 ^ _22342;
  wire _22344 = _12298 ? coded_block[932] : r932;
  wire _22345 = _12296 ? _22343 : _22344;
  always @ (posedge reset or posedge clock) if (reset) r932 <= 1'd0; else if (_12300) r932 <= _22345;
  wire [1:0] _22346 = {_0, _1886} + {_0, _3167};
  wire [1:0] _22347 = {_0, _5152} + {_0, _6303};
  wire [2:0] _22348 = {_0, _22346} + {_0, _22347};
  wire [1:0] _22349 = {_0, _9022} + {_0, _10654};
  wire [3:0] _22350 = {_0, _22348} + {_0, _0, _22349};
  wire _22351 = _12301 < _22350;
  wire _22352 = r931 ^ _22351;
  wire _22353 = _12298 ? coded_block[931] : r931;
  wire _22354 = _12296 ? _22352 : _22353;
  always @ (posedge reset or posedge clock) if (reset) r931 <= 1'd0; else if (_12300) r931 <= _22354;
  wire [1:0] _22355 = {_0, _1981} + {_0, _3773};
  wire [1:0] _22356 = {_0, _4958} + {_0, _6781};
  wire [2:0] _22357 = {_0, _22355} + {_0, _22356};
  wire [1:0] _22358 = {_0, _9406} + {_0, _11389};
  wire [3:0] _22359 = {_0, _22357} + {_0, _0, _22358};
  wire _22360 = _12301 < _22359;
  wire _22361 = r930 ^ _22360;
  wire _22362 = _12298 ? coded_block[930] : r930;
  wire _22363 = _12296 ? _22361 : _22362;
  always @ (posedge reset or posedge clock) if (reset) r930 <= 1'd0; else if (_12300) r930 <= _22363;
  wire [1:0] _22364 = {_0, _2013} + {_0, _3422};
  wire [1:0] _22365 = {_0, _5853} + {_0, _7036};
  wire [2:0] _22366 = {_0, _22364} + {_0, _22365};
  wire [1:0] _22367 = {_0, _8863} + {_0, _11485};
  wire [3:0] _22368 = {_0, _22366} + {_0, _0, _22367};
  wire _22369 = _12301 < _22368;
  wire _22370 = r929 ^ _22369;
  wire _22371 = _12298 ? coded_block[929] : r929;
  wire _22372 = _12296 ? _22370 : _22371;
  always @ (posedge reset or posedge clock) if (reset) r929 <= 1'd0; else if (_12300) r929 <= _22372;
  wire [1:0] _22373 = {_0, _2044} + {_0, _3646};
  wire [1:0] _22374 = {_0, _5501} + {_0, _7931};
  wire [2:0] _22375 = {_0, _22373} + {_0, _22374};
  wire [1:0] _22376 = {_0, _9118} + {_0, _10941};
  wire [3:0] _22377 = {_0, _22375} + {_0, _0, _22376};
  wire _22378 = _12301 < _22377;
  wire _22379 = r928 ^ _22378;
  wire _22380 = _12298 ? coded_block[928] : r928;
  wire _22381 = _12296 ? _22379 : _22380;
  always @ (posedge reset or posedge clock) if (reset) r928 <= 1'd0; else if (_12300) r928 <= _22381;
  wire [1:0] _22382 = {_0, _65} + {_0, _3517};
  wire [1:0] _22383 = {_0, _5726} + {_0, _7581};
  wire [2:0] _22384 = {_0, _22382} + {_0, _22383};
  wire [1:0] _22385 = {_0, _10014} + {_0, _11196};
  wire [3:0] _22386 = {_0, _22384} + {_0, _0, _22385};
  wire _22387 = _12301 < _22386;
  wire _22388 = r927 ^ _22387;
  wire _22389 = _12298 ? coded_block[927] : r927;
  wire _22390 = _12296 ? _22388 : _22389;
  always @ (posedge reset or posedge clock) if (reset) r927 <= 1'd0; else if (_12300) r927 <= _22390;
  wire [1:0] _22391 = {_0, _128} + {_0, _2592};
  wire [1:0] _22392 = {_0, _5949} + {_0, _7675};
  wire [2:0] _22393 = {_0, _22391} + {_0, _22392};
  wire [1:0] _22394 = {_0, _9886} + {_0, _11740};
  wire [3:0] _22395 = {_0, _22393} + {_0, _0, _22394};
  wire _22396 = _12301 < _22395;
  wire _22397 = r926 ^ _22396;
  wire _22398 = _12298 ? coded_block[926] : r926;
  wire _22399 = _12296 ? _22397 : _22398;
  always @ (posedge reset or posedge clock) if (reset) r926 <= 1'd0; else if (_12300) r926 <= _22399;
  wire [1:0] _22400 = {_0, _161} + {_0, _3198};
  wire [1:0] _22401 = {_0, _4671} + {_0, _8028};
  wire [2:0] _22402 = {_0, _22400} + {_0, _22401};
  wire [1:0] _22403 = {_0, _9759} + {_0, _11964};
  wire [3:0] _22404 = {_0, _22402} + {_0, _0, _22403};
  wire _22405 = _12301 < _22404;
  wire _22406 = r925 ^ _22405;
  wire _22407 = _12298 ? coded_block[925] : r925;
  wire _22408 = _12296 ? _22406 : _22407;
  always @ (posedge reset or posedge clock) if (reset) r925 <= 1'd0; else if (_12300) r925 <= _22408;
  wire [1:0] _22409 = {_0, _192} + {_0, _2750};
  wire [1:0] _22410 = {_0, _5279} + {_0, _6750};
  wire [2:0] _22411 = {_0, _22409} + {_0, _22410};
  wire [1:0] _22412 = {_0, _10108} + {_0, _11837};
  wire [3:0] _22413 = {_0, _22411} + {_0, _0, _22412};
  wire _22414 = _12301 < _22413;
  wire _22415 = r924 ^ _22414;
  wire _22416 = _12298 ? coded_block[924] : r924;
  wire _22417 = _12296 ? _22415 : _22416;
  always @ (posedge reset or posedge clock) if (reset) r924 <= 1'd0; else if (_12300) r924 <= _22417;
  wire [1:0] _22418 = {_0, _224} + {_0, _2367};
  wire [1:0] _22419 = {_0, _4830} + {_0, _7357};
  wire [2:0] _22420 = {_0, _22418} + {_0, _22419};
  wire [1:0] _22421 = {_0, _8830} + {_0, _12188};
  wire [3:0] _22422 = {_0, _22420} + {_0, _0, _22421};
  wire _22423 = _12301 < _22422;
  wire _22424 = r923 ^ _22423;
  wire _22425 = _12298 ? coded_block[923] : r923;
  wire _22426 = _12296 ? _22424 : _22425;
  always @ (posedge reset or posedge clock) if (reset) r923 <= 1'd0; else if (_12300) r923 <= _22426;
  wire [1:0] _22427 = {_0, _255} + {_0, _3390};
  wire [1:0] _22428 = {_0, _4447} + {_0, _6908};
  wire [2:0] _22429 = {_0, _22427} + {_0, _22428};
  wire [1:0] _22430 = {_0, _9438} + {_0, _10910};
  wire [3:0] _22431 = {_0, _22429} + {_0, _0, _22430};
  wire _22432 = _12301 < _22431;
  wire _22433 = r922 ^ _22432;
  wire _22434 = _12298 ? coded_block[922] : r922;
  wire _22435 = _12296 ? _22433 : _22434;
  always @ (posedge reset or posedge clock) if (reset) r922 <= 1'd0; else if (_12300) r922 <= _22435;
  wire [1:0] _22436 = {_0, _320} + {_0, _2271};
  wire [1:0] _22437 = {_0, _5884} + {_0, _7548};
  wire [2:0] _22438 = {_0, _22436} + {_0, _22437};
  wire [1:0] _22439 = {_0, _8607} + {_0, _11069};
  wire [3:0] _22440 = {_0, _22438} + {_0, _0, _22439};
  wire _22441 = _12301 < _22440;
  wire _22442 = r921 ^ _22441;
  wire _22443 = _12298 ? coded_block[921] : r921;
  wire _22444 = _12296 ? _22442 : _22443;
  always @ (posedge reset or posedge clock) if (reset) r921 <= 1'd0; else if (_12300) r921 <= _22444;
  wire [1:0] _22445 = {_0, _352} + {_0, _3709};
  wire [1:0] _22446 = {_0, _4350} + {_0, _7965};
  wire [2:0] _22447 = {_0, _22445} + {_0, _22446};
  wire [1:0] _22448 = {_0, _9630} + {_0, _10685};
  wire [3:0] _22449 = {_0, _22447} + {_0, _0, _22448};
  wire _22450 = _12301 < _22449;
  wire _22451 = r920 ^ _22450;
  wire _22452 = _12298 ? coded_block[920] : r920;
  wire _22453 = _12296 ? _22451 : _22452;
  always @ (posedge reset or posedge clock) if (reset) r920 <= 1'd0; else if (_12300) r920 <= _22453;
  wire [1:0] _22454 = {_0, _383} + {_0, _3005};
  wire [1:0] _22455 = {_0, _5790} + {_0, _6431};
  wire [2:0] _22456 = {_0, _22454} + {_0, _22455};
  wire [1:0] _22457 = {_0, _10045} + {_0, _11708};
  wire [3:0] _22458 = {_0, _22456} + {_0, _0, _22457};
  wire _22459 = _12301 < _22458;
  wire _22460 = r919 ^ _22459;
  wire _22461 = _12298 ? coded_block[919] : r919;
  wire _22462 = _12296 ? _22460 : _22461;
  always @ (posedge reset or posedge clock) if (reset) r919 <= 1'd0; else if (_12300) r919 <= _22462;
  wire [1:0] _22463 = {_0, _416} + {_0, _2686};
  wire [1:0] _22464 = {_0, _5085} + {_0, _7868};
  wire [2:0] _22465 = {_0, _22463} + {_0, _22464};
  wire [1:0] _22466 = {_0, _8511} + {_0, _12124};
  wire [3:0] _22467 = {_0, _22465} + {_0, _0, _22466};
  wire _22468 = _12301 < _22467;
  wire _22469 = r918 ^ _22468;
  wire _22470 = _12298 ? coded_block[918] : r918;
  wire _22471 = _12296 ? _22469 : _22470;
  always @ (posedge reset or posedge clock) if (reset) r918 <= 1'd0; else if (_12300) r918 <= _22471;
  wire [1:0] _22472 = {_0, _447} + {_0, _2847};
  wire [1:0] _22473 = {_0, _4767} + {_0, _7163};
  wire [2:0] _22474 = {_0, _22472} + {_0, _22473};
  wire [1:0] _22475 = {_0, _9949} + {_0, _10590};
  wire [3:0] _22476 = {_0, _22474} + {_0, _0, _22475};
  wire _22477 = _12301 < _22476;
  wire _22478 = r917 ^ _22477;
  wire _22479 = _12298 ? coded_block[917] : r917;
  wire _22480 = _12296 ? _22478 : _22479;
  always @ (posedge reset or posedge clock) if (reset) r917 <= 1'd0; else if (_12300) r917 <= _22480;
  wire [1:0] _22481 = {_0, _479} + {_0, _2655};
  wire [1:0] _22482 = {_0, _4926} + {_0, _6845};
  wire [2:0] _22483 = {_0, _22481} + {_0, _22482};
  wire [1:0] _22484 = {_0, _9248} + {_0, _12027};
  wire [3:0] _22485 = {_0, _22483} + {_0, _0, _22484};
  wire _22486 = _12301 < _22485;
  wire _22487 = r916 ^ _22486;
  wire _22488 = _12298 ? coded_block[916] : r916;
  wire _22489 = _12296 ? _22487 : _22488;
  always @ (posedge reset or posedge clock) if (reset) r916 <= 1'd0; else if (_12300) r916 <= _22489;
  wire [1:0] _22490 = {_0, _510} + {_0, _3037};
  wire [1:0] _22491 = {_0, _4734} + {_0, _7005};
  wire [2:0] _22492 = {_0, _22490} + {_0, _22491};
  wire [1:0] _22493 = {_0, _8926} + {_0, _11326};
  wire [3:0] _22494 = {_0, _22492} + {_0, _0, _22493};
  wire _22495 = _12301 < _22494;
  wire _22496 = r915 ^ _22495;
  wire _22497 = _12298 ? coded_block[915] : r915;
  wire _22498 = _12296 ? _22496 : _22497;
  always @ (posedge reset or posedge clock) if (reset) r915 <= 1'd0; else if (_12300) r915 <= _22498;
  wire [1:0] _22499 = {_0, _576} + {_0, _3964};
  wire [1:0] _22500 = {_0, _4256} + {_0, _7199};
  wire [2:0] _22501 = {_0, _22499} + {_0, _22500};
  wire [1:0] _22502 = {_0, _8894} + {_0, _11165};
  wire [3:0] _22503 = {_0, _22501} + {_0, _0, _22502};
  wire _22504 = _12301 < _22503;
  wire _22505 = r914 ^ _22504;
  wire _22506 = _12298 ? coded_block[914] : r914;
  wire _22507 = _12296 ? _22505 : _22506;
  always @ (posedge reset or posedge clock) if (reset) r914 <= 1'd0; else if (_12300) r914 <= _22507;
  wire [1:0] _22508 = {_0, _608} + {_0, _2526};
  wire [1:0] _22509 = {_0, _6045} + {_0, _6334};
  wire [2:0] _22510 = {_0, _22508} + {_0, _22509};
  wire [1:0] _22511 = {_0, _9279} + {_0, _10973};
  wire [3:0] _22512 = {_0, _22510} + {_0, _0, _22511};
  wire _22513 = _12301 < _22512;
  wire _22514 = r913 ^ _22513;
  wire _22515 = _12298 ? coded_block[913] : r913;
  wire _22516 = _12296 ? _22514 : _22515;
  always @ (posedge reset or posedge clock) if (reset) r913 <= 1'd0; else if (_12300) r913 <= _22516;
  wire [1:0] _22517 = {_0, _639} + {_0, _2463};
  wire [1:0] _22518 = {_0, _4605} + {_0, _8123};
  wire [2:0] _22519 = {_0, _22517} + {_0, _22518};
  wire [1:0] _22520 = {_0, _8415} + {_0, _11358};
  wire [3:0] _22521 = {_0, _22519} + {_0, _0, _22520};
  wire _22522 = _12301 < _22521;
  wire _22523 = r912 ^ _22522;
  wire _22524 = _12298 ? coded_block[912] : r912;
  wire _22525 = _12296 ? _22523 : _22524;
  always @ (posedge reset or posedge clock) if (reset) r912 <= 1'd0; else if (_12300) r912 <= _22525;
  wire [1:0] _22526 = {_0, _672} + {_0, _3580};
  wire [1:0] _22527 = {_0, _4542} + {_0, _6687};
  wire [2:0] _22528 = {_0, _22526} + {_0, _22527};
  wire [1:0] _22529 = {_0, _10204} + {_0, _10493};
  wire [3:0] _22530 = {_0, _22528} + {_0, _0, _22529};
  wire _22531 = _12301 < _22530;
  wire _22532 = r911 ^ _22531;
  wire _22533 = _12298 ? coded_block[911] : r911;
  wire _22534 = _12296 ? _22532 : _22533;
  always @ (posedge reset or posedge clock) if (reset) r911 <= 1'd0; else if (_12300) r911 <= _22534;
  wire [1:0] _22535 = {_0, _703} + {_0, _2239};
  wire [1:0] _22536 = {_0, _5663} + {_0, _6621};
  wire [2:0] _22537 = {_0, _22535} + {_0, _22536};
  wire [1:0] _22538 = {_0, _8767} + {_0, _12282};
  wire [3:0] _22539 = {_0, _22537} + {_0, _0, _22538};
  wire _22540 = _12301 < _22539;
  wire _22541 = r910 ^ _22540;
  wire _22542 = _12298 ? coded_block[910] : r910;
  wire _22543 = _12296 ? _22541 : _22542;
  always @ (posedge reset or posedge clock) if (reset) r910 <= 1'd0; else if (_12300) r910 <= _22543;
  wire [1:0] _22544 = {_0, _766} + {_0, _3549};
  wire [1:0] _22545 = {_0, _5918} + {_0, _6397};
  wire [2:0] _22546 = {_0, _22544} + {_0, _22545};
  wire [1:0] _22547 = {_0, _9822} + {_0, _10783};
  wire [3:0] _22548 = {_0, _22546} + {_0, _0, _22547};
  wire _22549 = _12301 < _22548;
  wire _22550 = r909 ^ _22549;
  wire _22551 = _12298 ? coded_block[909] : r909;
  wire _22552 = _12296 ? _22550 : _22551;
  always @ (posedge reset or posedge clock) if (reset) r909 <= 1'd0; else if (_12300) r909 <= _22552;
  wire [1:0] _22553 = {_0, _800} + {_0, _2494};
  wire [1:0] _22554 = {_0, _5628} + {_0, _7996};
  wire [2:0] _22555 = {_0, _22553} + {_0, _22554};
  wire [1:0] _22556 = {_0, _8480} + {_0, _11900};
  wire [3:0] _22557 = {_0, _22555} + {_0, _0, _22556};
  wire _22558 = _12301 < _22557;
  wire _22559 = r908 ^ _22558;
  wire _22560 = _12298 ? coded_block[908] : r908;
  wire _22561 = _12296 ? _22559 : _22560;
  always @ (posedge reset or posedge clock) if (reset) r908 <= 1'd0; else if (_12300) r908 <= _22561;
  wire [1:0] _22562 = {_0, _831} + {_0, _3997};
  wire [1:0] _22563 = {_0, _4574} + {_0, _7710};
  wire [2:0] _22564 = {_0, _22562} + {_0, _22563};
  wire [1:0] _22565 = {_0, _10077} + {_0, _10558};
  wire [3:0] _22566 = {_0, _22564} + {_0, _0, _22565};
  wire _22567 = _12301 < _22566;
  wire _22568 = r907 ^ _22567;
  wire _22569 = _12298 ? coded_block[907] : r907;
  wire _22570 = _12296 ? _22568 : _22569;
  always @ (posedge reset or posedge clock) if (reset) r907 <= 1'd0; else if (_12300) r907 <= _22570;
  wire [1:0] _22571 = {_0, _863} + {_0, _2974};
  wire [1:0] _22572 = {_0, _6076} + {_0, _6652};
  wire [2:0] _22573 = {_0, _22571} + {_0, _22572};
  wire [1:0] _22574 = {_0, _9790} + {_0, _12155};
  wire [3:0] _22575 = {_0, _22573} + {_0, _0, _22574};
  wire _22576 = _12301 < _22575;
  wire _22577 = r906 ^ _22576;
  wire _22578 = _12298 ? coded_block[906] : r906;
  wire _22579 = _12296 ? _22577 : _22578;
  always @ (posedge reset or posedge clock) if (reset) r906 <= 1'd0; else if (_12300) r906 <= _22579;
  wire [1:0] _22580 = {_0, _894} + {_0, _3742};
  wire [1:0] _22581 = {_0, _5053} + {_0, _8155};
  wire [2:0] _22582 = {_0, _22580} + {_0, _22581};
  wire [1:0] _22583 = {_0, _8736} + {_0, _11869};
  wire [3:0] _22584 = {_0, _22582} + {_0, _0, _22583};
  wire _22585 = _12301 < _22584;
  wire _22586 = r905 ^ _22585;
  wire _22587 = _12298 ? coded_block[905] : r905;
  wire _22588 = _12296 ? _22586 : _22587;
  always @ (posedge reset or posedge clock) if (reset) r905 <= 1'd0; else if (_12300) r905 <= _22588;
  wire [1:0] _22589 = {_0, _927} + {_0, _2910};
  wire [1:0] _22590 = {_0, _5821} + {_0, _7132};
  wire [2:0] _22591 = {_0, _22589} + {_0, _22590};
  wire [1:0] _22592 = {_0, _10235} + {_0, _10814};
  wire [3:0] _22593 = {_0, _22591} + {_0, _0, _22592};
  wire _22594 = _12301 < _22593;
  wire _22595 = r904 ^ _22594;
  wire _22596 = _12298 ? coded_block[904] : r904;
  wire _22597 = _12296 ? _22595 : _22596;
  always @ (posedge reset or posedge clock) if (reset) r904 <= 1'd0; else if (_12300) r904 <= _22597;
  wire [1:0] _22598 = {_0, _958} + {_0, _2430};
  wire [1:0] _22599 = {_0, _4989} + {_0, _7900};
  wire [2:0] _22600 = {_0, _22598} + {_0, _22599};
  wire [1:0] _22601 = {_0, _9212} + {_0, _10303};
  wire [3:0] _22602 = {_0, _22600} + {_0, _0, _22601};
  wire _22603 = _12301 < _22602;
  wire _22604 = r903 ^ _22603;
  wire _22605 = _12298 ? coded_block[903] : r903;
  wire _22606 = _12296 ? _22604 : _22605;
  always @ (posedge reset or posedge clock) if (reset) r903 <= 1'd0; else if (_12300) r903 <= _22606;
  wire [1:0] _22607 = {_0, _990} + {_0, _2557};
  wire [1:0] _22608 = {_0, _4511} + {_0, _7069};
  wire [2:0] _22609 = {_0, _22607} + {_0, _22608};
  wire [1:0] _22610 = {_0, _9980} + {_0, _11295};
  wire [3:0] _22611 = {_0, _22609} + {_0, _0, _22610};
  wire _22612 = _12301 < _22611;
  wire _22613 = r902 ^ _22612;
  wire _22614 = _12298 ? coded_block[902] : r902;
  wire _22615 = _12296 ? _22613 : _22614;
  always @ (posedge reset or posedge clock) if (reset) r902 <= 1'd0; else if (_12300) r902 <= _22615;
  wire [1:0] _22616 = {_0, _1021} + {_0, _3901};
  wire [1:0] _22617 = {_0, _4640} + {_0, _6589};
  wire [2:0] _22618 = {_0, _22616} + {_0, _22617};
  wire [1:0] _22619 = {_0, _9149} + {_0, _12061};
  wire [3:0] _22620 = {_0, _22618} + {_0, _0, _22619};
  wire _22621 = _12301 < _22620;
  wire _22622 = r901 ^ _22621;
  wire _22623 = _12298 ? coded_block[901] : r901;
  wire _22624 = _12296 ? _22622 : _22623;
  always @ (posedge reset or posedge clock) if (reset) r901 <= 1'd0; else if (_12300) r901 <= _22624;
  wire [1:0] _22625 = {_0, _1057} + {_0, _3135};
  wire [1:0] _22626 = {_0, _5981} + {_0, _6718};
  wire [2:0] _22627 = {_0, _22625} + {_0, _22626};
  wire [1:0] _22628 = {_0, _8670} + {_0, _11228};
  wire [3:0] _22629 = {_0, _22627} + {_0, _0, _22628};
  wire _22630 = _12301 < _22629;
  wire _22631 = r900 ^ _22630;
  wire _22632 = _12298 ? coded_block[900] : r900;
  wire _22633 = _12296 ? _22631 : _22632;
  always @ (posedge reset or posedge clock) if (reset) r900 <= 1'd0; else if (_12300) r900 <= _22633;
  wire [1:0] _22634 = {_0, _1088} + {_0, _3104};
  wire [1:0] _22635 = {_0, _5215} + {_0, _8059};
  wire [2:0] _22636 = {_0, _22634} + {_0, _22635};
  wire [1:0] _22637 = {_0, _8799} + {_0, _10748};
  wire [3:0] _22638 = {_0, _22636} + {_0, _0, _22637};
  wire _22639 = _12301 < _22638;
  wire _22640 = r899 ^ _22639;
  wire _22641 = _12298 ? coded_block[899] : r899;
  wire _22642 = _12296 ? _22640 : _22641;
  always @ (posedge reset or posedge clock) if (reset) r899 <= 1'd0; else if (_12300) r899 <= _22642;
  wire [1:0] _22643 = {_0, _1120} + {_0, _3933};
  wire [1:0] _22644 = {_0, _5183} + {_0, _7293};
  wire [2:0] _22645 = {_0, _22643} + {_0, _22644};
  wire [1:0] _22646 = {_0, _10141} + {_0, _10877};
  wire [3:0] _22647 = {_0, _22645} + {_0, _0, _22646};
  wire _22648 = _12301 < _22647;
  wire _22649 = r898 ^ _22648;
  wire _22650 = _12298 ? coded_block[898] : r898;
  wire _22651 = _12296 ? _22649 : _22650;
  always @ (posedge reset or posedge clock) if (reset) r898 <= 1'd0; else if (_12300) r898 <= _22651;
  wire [1:0] _22652 = {_0, _1151} + {_0, _2208};
  wire [1:0] _22653 = {_0, _6012} + {_0, _7262};
  wire [2:0] _22654 = {_0, _22652} + {_0, _22653};
  wire [1:0] _22655 = {_0, _9375} + {_0, _12219};
  wire [3:0] _22656 = {_0, _22654} + {_0, _0, _22655};
  wire _22657 = _12301 < _22656;
  wire _22658 = r897 ^ _22657;
  wire _22659 = _12298 ? coded_block[897] : r897;
  wire _22660 = _12296 ? _22658 : _22659;
  always @ (posedge reset or posedge clock) if (reset) r897 <= 1'd0; else if (_12300) r897 <= _22660;
  wire [1:0] _22661 = {_0, _1184} + {_0, _3615};
  wire [1:0] _22662 = {_0, _4287} + {_0, _8092};
  wire [2:0] _22663 = {_0, _22661} + {_0, _22662};
  wire [1:0] _22664 = {_0, _9342} + {_0, _11453};
  wire [3:0] _22665 = {_0, _22663} + {_0, _0, _22664};
  wire _22666 = _12301 < _22665;
  wire _22667 = r896 ^ _22666;
  wire _22668 = _12298 ? coded_block[896] : r896;
  wire _22669 = _12296 ? _22667 : _22668;
  always @ (posedge reset or posedge clock) if (reset) r896 <= 1'd0; else if (_12300) r896 <= _22669;
  wire [1:0] _22670 = {_0, _1215} + {_0, _3453};
  wire [1:0] _22671 = {_0, _5694} + {_0, _6366};
  wire [2:0] _22672 = {_0, _22670} + {_0, _22671};
  wire [1:0] _22673 = {_0, _10172} + {_0, _11422};
  wire [3:0] _22674 = {_0, _22672} + {_0, _0, _22673};
  wire _22675 = _12301 < _22674;
  wire _22676 = r895 ^ _22675;
  wire _22677 = _12298 ? coded_block[895] : r895;
  wire _22678 = _12296 ? _22676 : _22677;
  always @ (posedge reset or posedge clock) if (reset) r895 <= 1'd0; else if (_12300) r895 <= _22678;
  wire [1:0] _22679 = {_0, _1247} + {_0, _2081};
  wire [1:0] _22680 = {_0, _5534} + {_0, _7773};
  wire [2:0] _22681 = {_0, _22679} + {_0, _22680};
  wire [1:0] _22682 = {_0, _8446} + {_0, _12251};
  wire [3:0] _22683 = {_0, _22681} + {_0, _0, _22682};
  wire _22684 = _12301 < _22683;
  wire _22685 = r894 ^ _22684;
  wire _22686 = _12298 ? coded_block[894] : r894;
  wire _22687 = _12296 ? _22685 : _22686;
  always @ (posedge reset or posedge clock) if (reset) r894 <= 1'd0; else if (_12300) r894 <= _22687;
  wire [1:0] _22688 = {_0, _1278} + {_0, _3486};
  wire [1:0] _22689 = {_0, _4129} + {_0, _7612};
  wire [2:0] _22690 = {_0, _22688} + {_0, _22689};
  wire [1:0] _22691 = {_0, _9853} + {_0, _10527};
  wire [3:0] _22692 = {_0, _22690} + {_0, _0, _22691};
  wire _22693 = _12301 < _22692;
  wire _22694 = r893 ^ _22693;
  wire _22695 = _12298 ? coded_block[893] : r893;
  wire _22696 = _12296 ? _22694 : _22695;
  always @ (posedge reset or posedge clock) if (reset) r893 <= 1'd0; else if (_12300) r893 <= _22696;
  wire [1:0] _22697 = {_0, _1312} + {_0, _3678};
  wire [1:0] _22698 = {_0, _5565} + {_0, _6176};
  wire [2:0] _22699 = {_0, _22697} + {_0, _22698};
  wire [1:0] _22700 = {_0, _9693} + {_0, _11933};
  wire [3:0] _22701 = {_0, _22699} + {_0, _0, _22700};
  wire _22702 = _12301 < _22701;
  wire _22703 = r892 ^ _22702;
  wire _22704 = _12298 ? coded_block[892] : r892;
  wire _22705 = _12296 ? _22703 : _22704;
  always @ (posedge reset or posedge clock) if (reset) r892 <= 1'd0; else if (_12300) r892 <= _22705;
  wire [1:0] _22706 = {_0, _1343} + {_0, _2302};
  wire [1:0] _22707 = {_0, _5757} + {_0, _7644};
  wire [2:0] _22708 = {_0, _22706} + {_0, _22707};
  wire [1:0] _22709 = {_0, _8225} + {_0, _11771};
  wire [3:0] _22710 = {_0, _22708} + {_0, _0, _22709};
  wire _22711 = _12301 < _22710;
  wire _22712 = r891 ^ _22711;
  wire _22713 = _12298 ? coded_block[891] : r891;
  wire _22714 = _12296 ? _22712 : _22713;
  always @ (posedge reset or posedge clock) if (reset) r891 <= 1'd0; else if (_12300) r891 <= _22714;
  wire [1:0] _22715 = {_0, _1375} + {_0, _4060};
  wire [1:0] _22716 = {_0, _4384} + {_0, _7837};
  wire [2:0] _22717 = {_0, _22715} + {_0, _22716};
  wire [1:0] _22718 = {_0, _9724} + {_0, _10272};
  wire [3:0] _22719 = {_0, _22717} + {_0, _0, _22718};
  wire _22720 = _12301 < _22719;
  wire _22721 = r890 ^ _22720;
  wire _22722 = _12298 ? coded_block[890] : r890;
  wire _22723 = _12296 ? _22721 : _22722;
  always @ (posedge reset or posedge clock) if (reset) r890 <= 1'd0; else if (_12300) r890 <= _22723;
  wire [1:0] _22724 = {_0, _1406} + {_0, _3262};
  wire [1:0] _22725 = {_0, _6139} + {_0, _6462};
  wire [2:0] _22726 = {_0, _22724} + {_0, _22725};
  wire [1:0] _22727 = {_0, _9917} + {_0, _11806};
  wire [3:0] _22728 = {_0, _22726} + {_0, _0, _22727};
  wire _22729 = _12301 < _22728;
  wire _22730 = r889 ^ _22729;
  wire _22731 = _12298 ? coded_block[889] : r889;
  wire _22732 = _12296 ? _22730 : _22731;
  always @ (posedge reset or posedge clock) if (reset) r889 <= 1'd0; else if (_12300) r889 <= _22732;
  wire [1:0] _22733 = {_0, _1439} + {_0, _3325};
  wire [1:0] _22734 = {_0, _5342} + {_0, _6207};
  wire [2:0] _22735 = {_0, _22733} + {_0, _22734};
  wire [1:0] _22736 = {_0, _8543} + {_0, _11996};
  wire [3:0] _22737 = {_0, _22735} + {_0, _0, _22736};
  wire _22738 = _12301 < _22737;
  wire _22739 = r888 ^ _22738;
  wire _22740 = _12298 ? coded_block[888] : r888;
  wire _22741 = _12296 ? _22739 : _22740;
  always @ (posedge reset or posedge clock) if (reset) r888 <= 1'd0; else if (_12300) r888 <= _22741;
  wire [1:0] _22742 = {_0, _161} + {_0, _2974};
  wire [1:0] _22743 = {_0, _4223} + {_0, _6334};
  wire [2:0] _22744 = {_0, _22742} + {_0, _22743};
  wire [1:0] _22745 = {_0, _9181} + {_0, _11933};
  wire [3:0] _22746 = {_0, _22744} + {_0, _0, _22745};
  wire _22747 = _12301 < _22746;
  wire _22748 = r887 ^ _22747;
  wire _22749 = _12298 ? coded_block[887] : r887;
  wire _22750 = _12296 ? _22748 : _22749;
  always @ (posedge reset or posedge clock) if (reset) r887 <= 1'd0; else if (_12300) r887 <= _22750;
  wire [1:0] _22751 = {_0, _863} + {_0, _3997};
  wire [1:0] _22752 = {_0, _5053} + {_0, _7517};
  wire [2:0] _22753 = {_0, _22751} + {_0, _22752};
  wire [1:0] _22754 = {_0, _10045} + {_0, _11516};
  wire [3:0] _22755 = {_0, _22753} + {_0, _0, _22754};
  wire _22756 = _12301 < _22755;
  wire _22757 = r886 ^ _22756;
  wire _22758 = _12298 ? coded_block[886] : r886;
  wire _22759 = _12296 ? _22757 : _22758;
  always @ (posedge reset or posedge clock) if (reset) r886 <= 1'd0; else if (_12300) r886 <= _22759;
  wire [1:0] _22760 = {_0, _894} + {_0, _2399};
  wire [1:0] _22761 = {_0, _6076} + {_0, _7132};
  wire [2:0] _22762 = {_0, _22760} + {_0, _22761};
  wire [1:0] _22763 = {_0, _9597} + {_0, _12124};
  wire [3:0] _22764 = {_0, _22762} + {_0, _0, _22763};
  wire _22765 = _12301 < _22764;
  wire _22766 = r885 ^ _22765;
  wire _22767 = _12298 ? coded_block[885] : r885;
  wire _22768 = _12296 ? _22766 : _22767;
  always @ (posedge reset or posedge clock) if (reset) r885 <= 1'd0; else if (_12300) r885 <= _22768;
  wire [1:0] _22769 = {_0, _927} + {_0, _2878};
  wire [1:0] _22770 = {_0, _4478} + {_0, _8155};
  wire [2:0] _22771 = {_0, _22769} + {_0, _22770};
  wire [1:0] _22772 = {_0, _9212} + {_0, _11677};
  wire [3:0] _22773 = {_0, _22771} + {_0, _0, _22772};
  wire _22774 = _12301 < _22773;
  wire _22775 = r884 ^ _22774;
  wire _22776 = _12298 ? coded_block[884] : r884;
  wire _22777 = _12296 ? _22775 : _22776;
  always @ (posedge reset or posedge clock) if (reset) r884 <= 1'd0; else if (_12300) r884 <= _22777;
  wire [1:0] _22778 = {_0, _958} + {_0, _2302};
  wire [1:0] _22779 = {_0, _4958} + {_0, _6558};
  wire [2:0] _22780 = {_0, _22778} + {_0, _22779};
  wire [1:0] _22781 = {_0, _10235} + {_0, _11295};
  wire [3:0] _22782 = {_0, _22780} + {_0, _0, _22781};
  wire _22783 = _12301 < _22782;
  wire _22784 = r883 ^ _22783;
  wire _22785 = _12298 ? coded_block[883] : r883;
  wire _22786 = _12296 ? _22784 : _22785;
  always @ (posedge reset or posedge clock) if (reset) r883 <= 1'd0; else if (_12300) r883 <= _22786;
  wire [1:0] _22787 = {_0, _990} + {_0, _3615};
  wire [1:0] _22788 = {_0, _4384} + {_0, _7036};
  wire [2:0] _22789 = {_0, _22787} + {_0, _22788};
  wire [1:0] _22790 = {_0, _8638} + {_0, _10303};
  wire [3:0] _22791 = {_0, _22789} + {_0, _0, _22790};
  wire _22792 = _12301 < _22791;
  wire _22793 = r882 ^ _22792;
  wire _22794 = _12298 ? coded_block[882] : r882;
  wire _22795 = _12296 ? _22793 : _22794;
  always @ (posedge reset or posedge clock) if (reset) r882 <= 1'd0; else if (_12300) r882 <= _22795;
  wire [1:0] _22796 = {_0, _1021} + {_0, _3294};
  wire [1:0] _22797 = {_0, _5694} + {_0, _6462};
  wire [2:0] _22798 = {_0, _22796} + {_0, _22797};
  wire [1:0] _22799 = {_0, _9118} + {_0, _10717};
  wire [3:0] _22800 = {_0, _22798} + {_0, _0, _22799};
  wire _22801 = _12301 < _22800;
  wire _22802 = r881 ^ _22801;
  wire _22803 = _12298 ? coded_block[881] : r881;
  wire _22804 = _12296 ? _22802 : _22803;
  always @ (posedge reset or posedge clock) if (reset) r881 <= 1'd0; else if (_12300) r881 <= _22804;
  wire [1:0] _22805 = {_0, _1057} + {_0, _3453};
  wire [1:0] _22806 = {_0, _5373} + {_0, _7773};
  wire [2:0] _22807 = {_0, _22805} + {_0, _22806};
  wire [1:0] _22808 = {_0, _8543} + {_0, _11196};
  wire [3:0] _22809 = {_0, _22807} + {_0, _0, _22808};
  wire _22810 = _12301 < _22809;
  wire _22811 = r880 ^ _22810;
  wire _22812 = _12298 ? coded_block[880] : r880;
  wire _22813 = _12296 ? _22811 : _22812;
  always @ (posedge reset or posedge clock) if (reset) r880 <= 1'd0; else if (_12300) r880 <= _22813;
  wire [1:0] _22814 = {_0, _1088} + {_0, _3262};
  wire [1:0] _22815 = {_0, _5534} + {_0, _7454};
  wire [2:0] _22816 = {_0, _22814} + {_0, _22815};
  wire [1:0] _22817 = {_0, _9853} + {_0, _10621};
  wire [3:0] _22818 = {_0, _22816} + {_0, _0, _22817};
  wire _22819 = _12301 < _22818;
  wire _22820 = r879 ^ _22819;
  wire _22821 = _12298 ? coded_block[879] : r879;
  wire _22822 = _12296 ? _22820 : _22821;
  always @ (posedge reset or posedge clock) if (reset) r879 <= 1'd0; else if (_12300) r879 <= _22822;
  wire [1:0] _22823 = {_0, _1120} + {_0, _3646};
  wire [1:0] _22824 = {_0, _5342} + {_0, _7612};
  wire [2:0] _22825 = {_0, _22823} + {_0, _22824};
  wire [1:0] _22826 = {_0, _9534} + {_0, _11933};
  wire [3:0] _22827 = {_0, _22825} + {_0, _0, _22826};
  wire _22828 = _12301 < _22827;
  wire _22829 = r878 ^ _22828;
  wire _22830 = _12298 ? coded_block[878] : r878;
  wire _22831 = _12296 ? _22829 : _22830;
  always @ (posedge reset or posedge clock) if (reset) r878 <= 1'd0; else if (_12300) r878 <= _22831;
  wire [1:0] _22832 = {_0, _1151} + {_0, _2782};
  wire [1:0] _22833 = {_0, _5726} + {_0, _7420};
  wire [2:0] _22834 = {_0, _22832} + {_0, _22833};
  wire [1:0] _22835 = {_0, _9693} + {_0, _11613};
  wire [3:0] _22836 = {_0, _22834} + {_0, _0, _22835};
  wire _22837 = _12301 < _22836;
  wire _22838 = r877 ^ _22837;
  wire _22839 = _12298 ? coded_block[877] : r877;
  wire _22840 = _12296 ? _22838 : _22839;
  always @ (posedge reset or posedge clock) if (reset) r877 <= 1'd0; else if (_12300) r877 <= _22840;
  wire [1:0] _22841 = {_0, _1215} + {_0, _3135};
  wire [1:0] _22842 = {_0, _4640} + {_0, _6942};
  wire [2:0] _22843 = {_0, _22841} + {_0, _22842};
  wire [1:0] _22844 = {_0, _9886} + {_0, _11581};
  wire [3:0] _22845 = {_0, _22843} + {_0, _0, _22844};
  wire _22846 = _12301 < _22845;
  wire _22847 = r876 ^ _22846;
  wire _22848 = _12298 ? coded_block[876] : r876;
  wire _22849 = _12296 ? _22847 : _22848;
  always @ (posedge reset or posedge clock) if (reset) r876 <= 1'd0; else if (_12300) r876 <= _22849;
  wire [1:0] _22850 = {_0, _1247} + {_0, _3068};
  wire [1:0] _22851 = {_0, _5215} + {_0, _6718};
  wire [2:0] _22852 = {_0, _22850} + {_0, _22851};
  wire [1:0] _22853 = {_0, _9022} + {_0, _11964};
  wire [3:0] _22854 = {_0, _22852} + {_0, _0, _22853};
  wire _22855 = _12301 < _22854;
  wire _22856 = r875 ^ _22855;
  wire _22857 = _12298 ? coded_block[875] : r875;
  wire _22858 = _12296 ? _22856 : _22857;
  always @ (posedge reset or posedge clock) if (reset) r875 <= 1'd0; else if (_12300) r875 <= _22858;
  wire [1:0] _22859 = {_0, _1278} + {_0, _2175};
  wire [1:0] _22860 = {_0, _5152} + {_0, _7293};
  wire [2:0] _22861 = {_0, _22859} + {_0, _22860};
  wire [1:0] _22862 = {_0, _8799} + {_0, _11101};
  wire [3:0] _22863 = {_0, _22861} + {_0, _0, _22862};
  wire _22864 = _12301 < _22863;
  wire _22865 = r874 ^ _22864;
  wire _22866 = _12298 ? coded_block[874] : r874;
  wire _22867 = _12296 ? _22865 : _22866;
  always @ (posedge reset or posedge clock) if (reset) r874 <= 1'd0; else if (_12300) r874 <= _22867;
  wire [1:0] _22868 = {_0, _1312} + {_0, _2847};
  wire [1:0] _22869 = {_0, _4256} + {_0, _7230};
  wire [2:0] _22870 = {_0, _22868} + {_0, _22869};
  wire [1:0] _22871 = {_0, _9375} + {_0, _10877};
  wire [3:0] _22872 = {_0, _22870} + {_0, _0, _22871};
  wire _22873 = _12301 < _22872;
  wire _22874 = r873 ^ _22873;
  wire _22875 = _12298 ? coded_block[873] : r873;
  wire _22876 = _12296 ? _22874 : _22875;
  always @ (posedge reset or posedge clock) if (reset) r873 <= 1'd0; else if (_12300) r873 <= _22876;
  wire [1:0] _22877 = {_0, _1343} + {_0, _2430};
  wire [1:0] _22878 = {_0, _4926} + {_0, _6334};
  wire [2:0] _22879 = {_0, _22877} + {_0, _22878};
  wire [1:0] _22880 = {_0, _9311} + {_0, _11453};
  wire [3:0] _22881 = {_0, _22879} + {_0, _0, _22880};
  wire _22882 = _12301 < _22881;
  wire _22883 = r872 ^ _22882;
  wire _22884 = _12298 ? coded_block[872] : r872;
  wire _22885 = _12296 ? _22883 : _22884;
  always @ (posedge reset or posedge clock) if (reset) r872 <= 1'd0; else if (_12300) r872 <= _22885;
  wire [1:0] _22886 = {_0, _1375} + {_0, _2144};
  wire [1:0] _22887 = {_0, _4511} + {_0, _7005};
  wire [2:0] _22888 = {_0, _22886} + {_0, _22887};
  wire [1:0] _22889 = {_0, _8415} + {_0, _11389};
  wire [3:0] _22890 = {_0, _22888} + {_0, _0, _22889};
  wire _22891 = _12301 < _22890;
  wire _22892 = r871 ^ _22891;
  wire _22893 = _12298 ? coded_block[871] : r871;
  wire _22894 = _12296 ? _22892 : _22893;
  always @ (posedge reset or posedge clock) if (reset) r871 <= 1'd0; else if (_12300) r871 <= _22894;
  wire [1:0] _22895 = {_0, _1406} + {_0, _3104};
  wire [1:0] _22896 = {_0, _4223} + {_0, _6589};
  wire [2:0] _22897 = {_0, _22895} + {_0, _22896};
  wire [1:0] _22898 = {_0, _9085} + {_0, _10493};
  wire [3:0] _22899 = {_0, _22897} + {_0, _0, _22898};
  wire _22900 = _12301 < _22899;
  wire _22901 = r870 ^ _22900;
  wire _22902 = _12298 ? coded_block[870] : r870;
  wire _22903 = _12296 ? _22901 : _22902;
  always @ (posedge reset or posedge clock) if (reset) r870 <= 1'd0; else if (_12300) r870 <= _22903;
  wire [1:0] _22904 = {_0, _1439} + {_0, _2592};
  wire [1:0] _22905 = {_0, _5183} + {_0, _6303};
  wire [2:0] _22906 = {_0, _22904} + {_0, _22905};
  wire [1:0] _22907 = {_0, _8670} + {_0, _11165};
  wire [3:0] _22908 = {_0, _22906} + {_0, _0, _22907};
  wire _22909 = _12301 < _22908;
  wire _22910 = r869 ^ _22909;
  wire _22911 = _12298 ? coded_block[869] : r869;
  wire _22912 = _12296 ? _22910 : _22911;
  always @ (posedge reset or posedge clock) if (reset) r869 <= 1'd0; else if (_12300) r869 <= _22912;
  wire [1:0] _22913 = {_0, _1470} + {_0, _3580};
  wire [1:0] _22914 = {_0, _4671} + {_0, _7262};
  wire [2:0] _22915 = {_0, _22913} + {_0, _22914};
  wire [1:0] _22916 = {_0, _8383} + {_0, _10748};
  wire [3:0] _22917 = {_0, _22915} + {_0, _0, _22916};
  wire _22918 = _12301 < _22917;
  wire _22919 = r868 ^ _22918;
  wire _22920 = _12298 ? coded_block[868] : r868;
  wire _22921 = _12296 ? _22919 : _22920;
  always @ (posedge reset or posedge clock) if (reset) r868 <= 1'd0; else if (_12300) r868 <= _22921;
  wire [1:0] _22922 = {_0, _1502} + {_0, _2336};
  wire [1:0] _22923 = {_0, _5663} + {_0, _6750};
  wire [2:0] _22924 = {_0, _22922} + {_0, _22923};
  wire [1:0] _22925 = {_0, _9342} + {_0, _10462};
  wire [3:0] _22926 = {_0, _22924} + {_0, _0, _22925};
  wire _22927 = _12301 < _22926;
  wire _22928 = r867 ^ _22927;
  wire _22929 = _12298 ? coded_block[867] : r867;
  wire _22930 = _12296 ? _22928 : _22929;
  always @ (posedge reset or posedge clock) if (reset) r867 <= 1'd0; else if (_12300) r867 <= _22930;
  wire [1:0] _22931 = {_0, _1599} + {_0, _3167};
  wire [1:0] _22932 = {_0, _5116} + {_0, _7675};
  wire [2:0] _22933 = {_0, _22931} + {_0, _22932};
  wire [1:0] _22934 = {_0, _8574} + {_0, _11900};
  wire [3:0] _22935 = {_0, _22933} + {_0, _0, _22934};
  wire _22936 = _12301 < _22935;
  wire _22937 = r866 ^ _22936;
  wire _22938 = _12298 ? coded_block[866] : r866;
  wire _22939 = _12296 ? _22937 : _22938;
  always @ (posedge reset or posedge clock) if (reset) r866 <= 1'd0; else if (_12300) r866 <= _22939;
  wire [1:0] _22940 = {_0, _1631} + {_0, _2494};
  wire [1:0] _22941 = {_0, _5246} + {_0, _7199};
  wire [2:0] _22942 = {_0, _22940} + {_0, _22941};
  wire [1:0] _22943 = {_0, _9759} + {_0, _10654};
  wire [3:0] _22944 = {_0, _22942} + {_0, _0, _22943};
  wire _22945 = _12301 < _22944;
  wire _22946 = r865 ^ _22945;
  wire _22947 = _12298 ? coded_block[865] : r865;
  wire _22948 = _12296 ? _22946 : _22947;
  always @ (posedge reset or posedge clock) if (reset) r865 <= 1'd0; else if (_12300) r865 <= _22948;
  wire [1:0] _22949 = {_0, _1695} + {_0, _3709};
  wire [1:0] _22950 = {_0, _5821} + {_0, _6652};
  wire [2:0] _22951 = {_0, _22949} + {_0, _22950};
  wire [1:0] _22952 = {_0, _9406} + {_0, _11358};
  wire [3:0] _22953 = {_0, _22951} + {_0, _0, _22952};
  wire _22954 = _12301 < _22953;
  wire _22955 = r864 ^ _22954;
  wire _22956 = _12298 ? coded_block[864] : r864;
  wire _22957 = _12296 ? _22955 : _22956;
  always @ (posedge reset or posedge clock) if (reset) r864 <= 1'd0; else if (_12300) r864 <= _22957;
  wire [1:0] _22958 = {_0, _1726} + {_0, _2526};
  wire [1:0] _22959 = {_0, _5790} + {_0, _7900};
  wire [2:0] _22960 = {_0, _22958} + {_0, _22959};
  wire [1:0] _22961 = {_0, _8736} + {_0, _11485};
  wire [3:0] _22962 = {_0, _22960} + {_0, _0, _22961};
  wire _22963 = _12301 < _22962;
  wire _22964 = r863 ^ _22963;
  wire _22965 = _12298 ? coded_block[863] : r863;
  wire _22966 = _12296 ? _22964 : _22965;
  always @ (posedge reset or posedge clock) if (reset) r863 <= 1'd0; else if (_12300) r863 <= _22966;
  wire [1:0] _22967 = {_0, _1758} + {_0, _2813};
  wire [1:0] _22968 = {_0, _4605} + {_0, _7868};
  wire [2:0] _22969 = {_0, _22967} + {_0, _22968};
  wire [1:0] _22970 = {_0, _9980} + {_0, _10814};
  wire [3:0] _22971 = {_0, _22969} + {_0, _0, _22970};
  wire _22972 = _12301 < _22971;
  wire _22973 = r862 ^ _22972;
  wire _22974 = _12298 ? coded_block[862] : r862;
  wire _22975 = _12296 ? _22973 : _22974;
  always @ (posedge reset or posedge clock) if (reset) r862 <= 1'd0; else if (_12300) r862 <= _22975;
  wire [1:0] _22976 = {_0, _1789} + {_0, _2208};
  wire [1:0] _22977 = {_0, _4895} + {_0, _6687};
  wire [2:0] _22978 = {_0, _22976} + {_0, _22977};
  wire [1:0] _22979 = {_0, _9949} + {_0, _12061};
  wire [3:0] _22980 = {_0, _22978} + {_0, _0, _22979};
  wire _22981 = _12301 < _22980;
  wire _22982 = r861 ^ _22981;
  wire _22983 = _12298 ? coded_block[861] : r861;
  wire _22984 = _12296 ? _22982 : _22983;
  always @ (posedge reset or posedge clock) if (reset) r861 <= 1'd0; else if (_12300) r861 <= _22984;
  wire [1:0] _22985 = {_0, _1823} + {_0, _4060};
  wire [1:0] _22986 = {_0, _4287} + {_0, _6973};
  wire [2:0] _22987 = {_0, _22985} + {_0, _22986};
  wire [1:0] _22988 = {_0, _8767} + {_0, _12027};
  wire [3:0] _22989 = {_0, _22987} + {_0, _0, _22988};
  wire _22990 = _12301 < _22989;
  wire _22991 = r860 ^ _22990;
  wire _22992 = _12298 ? coded_block[860] : r860;
  wire _22993 = _12296 ? _22991 : _22992;
  always @ (posedge reset or posedge clock) if (reset) r860 <= 1'd0; else if (_12300) r860 <= _22993;
  wire [1:0] _22994 = {_0, _1854} + {_0, _2081};
  wire [1:0] _22995 = {_0, _6139} + {_0, _6366};
  wire [2:0] _22996 = {_0, _22994} + {_0, _22995};
  wire [1:0] _22997 = {_0, _9054} + {_0, _10846};
  wire [3:0] _22998 = {_0, _22996} + {_0, _0, _22997};
  wire _22999 = _12301 < _22998;
  wire _23000 = r859 ^ _22999;
  wire _23001 = _12298 ? coded_block[859] : r859;
  wire _23002 = _12296 ? _23000 : _23001;
  always @ (posedge reset or posedge clock) if (reset) r859 <= 1'd0; else if (_12300) r859 <= _23002;
  wire [1:0] _23003 = {_0, _1886} + {_0, _4091};
  wire [1:0] _23004 = {_0, _4129} + {_0, _6207};
  wire [2:0] _23005 = {_0, _23003} + {_0, _23004};
  wire [1:0] _23006 = {_0, _8446} + {_0, _11132};
  wire [3:0] _23007 = {_0, _23005} + {_0, _0, _23006};
  wire _23008 = _12301 < _23007;
  wire _23009 = r858 ^ _23008;
  wire _23010 = _12298 ? coded_block[858] : r858;
  wire _23011 = _12296 ? _23009 : _23010;
  always @ (posedge reset or posedge clock) if (reset) r858 <= 1'd0; else if (_12300) r858 <= _23011;
  wire [1:0] _23012 = {_0, _1917} + {_0, _2271};
  wire [1:0] _23013 = {_0, _4160} + {_0, _6176};
  wire [2:0] _23014 = {_0, _23012} + {_0, _23013};
  wire [1:0] _23015 = {_0, _8288} + {_0, _10527};
  wire [3:0] _23016 = {_0, _23014} + {_0, _0, _23015};
  wire _23017 = _12301 < _23016;
  wire _23018 = r857 ^ _23017;
  wire _23019 = _12298 ? coded_block[857] : r857;
  wire _23020 = _12296 ? _23018 : _23019;
  always @ (posedge reset or posedge clock) if (reset) r857 <= 1'd0; else if (_12300) r857 <= _23020;
  wire [1:0] _23021 = {_0, _1981} + {_0, _2655};
  wire [1:0] _23022 = {_0, _4989} + {_0, _6431};
  wire [2:0] _23023 = {_0, _23021} + {_0, _23022};
  wire [1:0] _23024 = {_0, _8319} + {_0, _10272};
  wire [3:0] _23025 = {_0, _23023} + {_0, _0, _23024};
  wire _23026 = _12301 < _23025;
  wire _23027 = r856 ^ _23026;
  wire _23028 = _12298 ? coded_block[856] : r856;
  wire _23029 = _12296 ? _23027 : _23028;
  always @ (posedge reset or posedge clock) if (reset) r856 <= 1'd0; else if (_12300) r856 <= _23029;
  wire [1:0] _23030 = {_0, _2013} + {_0, _3870};
  wire [1:0] _23031 = {_0, _4734} + {_0, _7069};
  wire [2:0] _23032 = {_0, _23030} + {_0, _23031};
  wire [1:0] _23033 = {_0, _8511} + {_0, _10399};
  wire [3:0] _23034 = {_0, _23032} + {_0, _0, _23033};
  wire _23035 = _12301 < _23034;
  wire _23036 = r855 ^ _23035;
  wire _23037 = _12298 ? coded_block[855] : r855;
  wire _23038 = _12296 ? _23036 : _23037;
  always @ (posedge reset or posedge clock) if (reset) r855 <= 1'd0; else if (_12300) r855 <= _23038;
  wire [1:0] _23039 = {_0, _65} + {_0, _2719};
  wire [1:0] _23040 = {_0, _6012} + {_0, _8028};
  wire [2:0] _23041 = {_0, _23039} + {_0, _23040};
  wire [1:0] _23042 = {_0, _8894} + {_0, _11228};
  wire [3:0] _23043 = {_0, _23041} + {_0, _0, _23042};
  wire _23044 = _12301 < _23043;
  wire _23045 = r854 ^ _23044;
  wire _23046 = _12298 ? coded_block[854] : r854;
  wire _23047 = _12296 ? _23045 : _23046;
  always @ (posedge reset or posedge clock) if (reset) r854 <= 1'd0; else if (_12300) r854 <= _23047;
  wire [1:0] _23048 = {_0, _97} + {_0, _3422};
  wire [1:0] _23049 = {_0, _4798} + {_0, _8092};
  wire [2:0] _23050 = {_0, _23048} + {_0, _23049};
  wire [1:0] _23051 = {_0, _10108} + {_0, _10973};
  wire [3:0] _23052 = {_0, _23050} + {_0, _0, _23051};
  wire _23053 = _12301 < _23052;
  wire _23054 = r853 ^ _23053;
  wire _23055 = _12298 ? coded_block[853] : r853;
  wire _23056 = _12296 ? _23054 : _23055;
  always @ (posedge reset or posedge clock) if (reset) r853 <= 1'd0; else if (_12300) r853 <= _23056;
  wire [1:0] _23057 = {_0, _128} + {_0, _3325};
  wire [1:0] _23058 = {_0, _5501} + {_0, _6877};
  wire [2:0] _23059 = {_0, _23057} + {_0, _23058};
  wire [1:0] _23060 = {_0, _10172} + {_0, _12188};
  wire [3:0] _23061 = {_0, _23059} + {_0, _0, _23060};
  wire _23062 = _12301 < _23061;
  wire _23063 = r852 ^ _23062;
  wire _23064 = _12298 ? coded_block[852] : r852;
  wire _23065 = _12296 ? _23063 : _23064;
  always @ (posedge reset or posedge clock) if (reset) r852 <= 1'd0; else if (_12300) r852 <= _23065;
  wire [1:0] _23066 = {_0, _161} + {_0, _3836};
  wire [1:0] _23067 = {_0, _5407} + {_0, _7581};
  wire [2:0] _23068 = {_0, _23066} + {_0, _23067};
  wire [1:0] _23069 = {_0, _8957} + {_0, _12251};
  wire [3:0] _23070 = {_0, _23068} + {_0, _0, _23069};
  wire _23071 = _12301 < _23070;
  wire _23072 = r851 ^ _23071;
  wire _23073 = _12298 ? coded_block[851] : r851;
  wire _23074 = _12296 ? _23072 : _23073;
  always @ (posedge reset or posedge clock) if (reset) r851 <= 1'd0; else if (_12300) r851 <= _23074;
  wire [1:0] _23075 = {_0, _192} + {_0, _2686};
  wire [1:0] _23076 = {_0, _5918} + {_0, _7485};
  wire [2:0] _23077 = {_0, _23075} + {_0, _23076};
  wire [1:0] _23078 = {_0, _9661} + {_0, _11038};
  wire [3:0] _23079 = {_0, _23077} + {_0, _0, _23078};
  wire _23080 = _12301 < _23079;
  wire _23081 = r850 ^ _23080;
  wire _23082 = _12298 ? coded_block[850] : r850;
  wire _23083 = _12296 ? _23081 : _23082;
  always @ (posedge reset or posedge clock) if (reset) r850 <= 1'd0; else if (_12300) r850 <= _23083;
  wire [1:0] _23084 = {_0, _224} + {_0, _3964};
  wire [1:0] _23085 = {_0, _4767} + {_0, _7996};
  wire [2:0] _23086 = {_0, _23084} + {_0, _23085};
  wire [1:0] _23087 = {_0, _9566} + {_0, _11740};
  wire [3:0] _23088 = {_0, _23086} + {_0, _0, _23087};
  wire _23089 = _12301 < _23088;
  wire _23090 = r849 ^ _23089;
  wire _23091 = _12298 ? coded_block[849] : r849;
  wire _23092 = _12296 ? _23090 : _23091;
  always @ (posedge reset or posedge clock) if (reset) r849 <= 1'd0; else if (_12300) r849 <= _23092;
  wire [1:0] _23093 = {_0, _255} + {_0, _3005};
  wire [1:0] _23094 = {_0, _6045} + {_0, _6845};
  wire [2:0] _23095 = {_0, _23093} + {_0, _23094};
  wire [1:0] _23096 = {_0, _10077} + {_0, _11644};
  wire [3:0] _23097 = {_0, _23095} + {_0, _0, _23096};
  wire _23098 = _12301 < _23097;
  wire _23099 = r848 ^ _23098;
  wire _23100 = _12298 ? coded_block[848] : r848;
  wire _23101 = _12296 ? _23099 : _23100;
  always @ (posedge reset or posedge clock) if (reset) r848 <= 1'd0; else if (_12300) r848 <= _23101;
  wire [1:0] _23102 = {_0, _289} + {_0, _3549};
  wire [1:0] _23103 = {_0, _5085} + {_0, _8123};
  wire [2:0] _23104 = {_0, _23102} + {_0, _23103};
  wire [1:0] _23105 = {_0, _8926} + {_0, _12155};
  wire [3:0] _23106 = {_0, _23104} + {_0, _0, _23105};
  wire _23107 = _12301 < _23106;
  wire _23108 = r847 ^ _23107;
  wire _23109 = _12298 ? coded_block[847] : r847;
  wire _23110 = _12296 ? _23108 : _23109;
  always @ (posedge reset or posedge clock) if (reset) r847 <= 1'd0; else if (_12300) r847 <= _23110;
  wire [1:0] _23111 = {_0, _320} + {_0, _2623};
  wire [1:0] _23112 = {_0, _5628} + {_0, _7163};
  wire [2:0] _23113 = {_0, _23111} + {_0, _23112};
  wire [1:0] _23114 = {_0, _10204} + {_0, _11004};
  wire [3:0] _23115 = {_0, _23113} + {_0, _0, _23114};
  wire _23116 = _12301 < _23115;
  wire _23117 = r846 ^ _23116;
  wire _23118 = _12298 ? coded_block[846] : r846;
  wire _23119 = _12296 ? _23117 : _23118;
  always @ (posedge reset or posedge clock) if (reset) r846 <= 1'd0; else if (_12300) r846 <= _23119;
  wire [1:0] _23120 = {_0, _352} + {_0, _2941};
  wire [1:0] _23121 = {_0, _4703} + {_0, _7710};
  wire [2:0] _23122 = {_0, _23120} + {_0, _23121};
  wire [1:0] _23123 = {_0, _9248} + {_0, _12282};
  wire [3:0] _23124 = {_0, _23122} + {_0, _0, _23123};
  wire _23125 = _12301 < _23124;
  wire _23126 = r845 ^ _23125;
  wire _23127 = _12298 ? coded_block[845] : r845;
  wire _23128 = _12296 ? _23126 : _23127;
  always @ (posedge reset or posedge clock) if (reset) r845 <= 1'd0; else if (_12300) r845 <= _23128;
  wire [1:0] _23129 = {_0, _383} + {_0, _3390};
  wire [1:0] _23130 = {_0, _5022} + {_0, _6781};
  wire [2:0] _23131 = {_0, _23129} + {_0, _23130};
  wire [1:0] _23132 = {_0, _9790} + {_0, _11326};
  wire [3:0] _23133 = {_0, _23131} + {_0, _0, _23132};
  wire _23134 = _12301 < _23133;
  wire _23135 = r844 ^ _23134;
  wire _23136 = _12298 ? coded_block[844] : r844;
  wire _23137 = _12296 ? _23135 : _23136;
  always @ (posedge reset or posedge clock) if (reset) r844 <= 1'd0; else if (_12300) r844 <= _23137;
  wire [1:0] _23138 = {_0, _416} + {_0, _2750};
  wire [1:0] _23139 = {_0, _5470} + {_0, _7100};
  wire [2:0] _23140 = {_0, _23138} + {_0, _23139};
  wire [1:0] _23141 = {_0, _8863} + {_0, _11869};
  wire [3:0] _23142 = {_0, _23140} + {_0, _0, _23141};
  wire _23143 = _12301 < _23142;
  wire _23144 = r843 ^ _23143;
  wire _23145 = _12298 ? coded_block[843] : r843;
  wire _23146 = _12296 ? _23144 : _23145;
  always @ (posedge reset or posedge clock) if (reset) r843 <= 1'd0; else if (_12300) r843 <= _23146;
  wire [1:0] _23147 = {_0, _447} + {_0, _3678};
  wire [1:0] _23148 = {_0, _4830} + {_0, _7548};
  wire [2:0] _23149 = {_0, _23147} + {_0, _23148};
  wire [1:0] _23150 = {_0, _9181} + {_0, _10941};
  wire [3:0] _23151 = {_0, _23149} + {_0, _0, _23150};
  wire _23152 = _12301 < _23151;
  wire _23153 = r842 ^ _23152;
  wire _23154 = _12298 ? coded_block[842] : r842;
  wire _23155 = _12296 ? _23153 : _23154;
  always @ (posedge reset or posedge clock) if (reset) r842 <= 1'd0; else if (_12300) r842 <= _23155;
  wire [1:0] _23156 = {_0, _479} + {_0, _3773};
  wire [1:0] _23157 = {_0, _5757} + {_0, _6908};
  wire [2:0] _23158 = {_0, _23156} + {_0, _23157};
  wire [1:0] _23159 = {_0, _9630} + {_0, _11259};
  wire [3:0] _23160 = {_0, _23158} + {_0, _0, _23159};
  wire _23161 = _12301 < _23160;
  wire _23162 = r841 ^ _23161;
  wire _23163 = _12298 ? coded_block[841] : r841;
  wire _23164 = _12296 ? _23162 : _23163;
  always @ (posedge reset or posedge clock) if (reset) r841 <= 1'd0; else if (_12300) r841 <= _23164;
  wire [1:0] _23165 = {_0, _510} + {_0, _3231};
  wire [1:0] _23166 = {_0, _5853} + {_0, _7837};
  wire [2:0] _23167 = {_0, _23165} + {_0, _23166};
  wire [1:0] _23168 = {_0, _8991} + {_0, _11708};
  wire [3:0] _23169 = {_0, _23167} + {_0, _0, _23168};
  wire _23170 = _12301 < _23169;
  wire _23171 = r840 ^ _23170;
  wire _23172 = _12298 ? coded_block[840] : r840;
  wire _23173 = _12296 ? _23171 : _23172;
  always @ (posedge reset or posedge clock) if (reset) r840 <= 1'd0; else if (_12300) r840 <= _23173;
  wire [1:0] _23174 = {_0, _545} + {_0, _3486};
  wire [1:0] _23175 = {_0, _5310} + {_0, _7931};
  wire [2:0] _23176 = {_0, _23174} + {_0, _23175};
  wire [1:0] _23177 = {_0, _9917} + {_0, _11069};
  wire [3:0] _23178 = {_0, _23176} + {_0, _0, _23177};
  wire _23179 = _12301 < _23178;
  wire _23180 = r839 ^ _23179;
  wire _23181 = _12298 ? coded_block[839] : r839;
  wire _23182 = _12296 ? _23180 : _23181;
  always @ (posedge reset or posedge clock) if (reset) r839 <= 1'd0; else if (_12300) r839 <= _23182;
  wire [1:0] _23183 = {_0, _576} + {_0, _2367};
  wire [1:0] _23184 = {_0, _5565} + {_0, _7389};
  wire [2:0] _23185 = {_0, _23183} + {_0, _23184};
  wire [1:0] _23186 = {_0, _10014} + {_0, _11996};
  wire [3:0] _23187 = {_0, _23185} + {_0, _0, _23186};
  wire _23188 = _12301 < _23187;
  wire _23189 = r838 ^ _23188;
  wire _23190 = _12298 ? coded_block[838] : r838;
  wire _23191 = _12296 ? _23189 : _23190;
  always @ (posedge reset or posedge clock) if (reset) r838 <= 1'd0; else if (_12300) r838 <= _23191;
  wire [1:0] _23192 = {_0, _608} + {_0, _4028};
  wire [1:0] _23193 = {_0, _4447} + {_0, _7644};
  wire [2:0] _23194 = {_0, _23192} + {_0, _23193};
  wire [1:0] _23195 = {_0, _9469} + {_0, _12092};
  wire [3:0] _23196 = {_0, _23194} + {_0, _0, _23195};
  wire _23197 = _12301 < _23196;
  wire _23198 = r837 ^ _23197;
  wire _23199 = _12298 ? coded_block[837] : r837;
  wire _23200 = _12296 ? _23198 : _23199;
  always @ (posedge reset or posedge clock) if (reset) r837 <= 1'd0; else if (_12300) r837 <= _23200;
  wire [1:0] _23201 = {_0, _639} + {_0, _2239};
  wire [1:0] _23202 = {_0, _6108} + {_0, _6525};
  wire [2:0] _23203 = {_0, _23201} + {_0, _23202};
  wire [1:0] _23204 = {_0, _9724} + {_0, _11550};
  wire [3:0] _23205 = {_0, _23203} + {_0, _0, _23204};
  wire _23206 = _12301 < _23205;
  wire _23207 = r836 ^ _23206;
  wire _23208 = _12298 ? coded_block[836] : r836;
  wire _23209 = _12296 ? _23207 : _23208;
  always @ (posedge reset or posedge clock) if (reset) r836 <= 1'd0; else if (_12300) r836 <= _23209;
  wire [1:0] _23210 = {_0, _703} + {_0, _2463};
  wire [1:0] _23211 = {_0, _4192} + {_0, _6397};
  wire [2:0] _23212 = {_0, _23210} + {_0, _23211};
  wire [1:0] _23213 = {_0, _8256} + {_0, _10685};
  wire [3:0] _23214 = {_0, _23212} + {_0, _0, _23213};
  wire _23215 = _12301 < _23214;
  wire _23216 = r835 ^ _23215;
  wire _23217 = _12298 ? coded_block[835] : r835;
  wire _23218 = _12296 ? _23216 : _23217;
  always @ (posedge reset or posedge clock) if (reset) r835 <= 1'd0; else if (_12300) r835 <= _23218;
  wire [1:0] _23219 = {_0, _735} + {_0, _3198};
  wire [1:0] _23220 = {_0, _4542} + {_0, _6270};
  wire [2:0] _23221 = {_0, _23219} + {_0, _23220};
  wire [1:0] _23222 = {_0, _8480} + {_0, _10335};
  wire [3:0] _23223 = {_0, _23221} + {_0, _0, _23222};
  wire _23224 = _12301 < _23223;
  wire _23225 = r834 ^ _23224;
  wire _23226 = _12298 ? coded_block[834] : r834;
  wire _23227 = _12296 ? _23225 : _23226;
  always @ (posedge reset or posedge clock) if (reset) r834 <= 1'd0; else if (_12300) r834 <= _23227;
  wire [1:0] _23228 = {_0, _766} + {_0, _3805};
  wire [1:0] _23229 = {_0, _5279} + {_0, _6621};
  wire [2:0] _23230 = {_0, _23228} + {_0, _23229};
  wire [1:0] _23231 = {_0, _8352} + {_0, _10558};
  wire [3:0] _23232 = {_0, _23230} + {_0, _0, _23231};
  wire _23233 = _12301 < _23232;
  wire _23234 = r833 ^ _23233;
  wire _23235 = _12298 ? coded_block[833] : r833;
  wire _23236 = _12296 ? _23234 : _23235;
  always @ (posedge reset or posedge clock) if (reset) r833 <= 1'd0; else if (_12300) r833 <= _23236;
  wire [1:0] _23237 = {_0, _800} + {_0, _3359};
  wire [1:0] _23238 = {_0, _5884} + {_0, _7357};
  wire [2:0] _23239 = {_0, _23237} + {_0, _23238};
  wire [1:0] _23240 = {_0, _8701} + {_0, _10430};
  wire [3:0] _23241 = {_0, _23239} + {_0, _0, _23240};
  wire _23242 = _12301 < _23241;
  wire _23243 = r832 ^ _23242;
  wire _23244 = _12298 ? coded_block[832] : r832;
  wire _23245 = _12296 ? _23243 : _23244;
  always @ (posedge reset or posedge clock) if (reset) r832 <= 1'd0; else if (_12300) r832 <= _23245;
  wire [1:0] _23246 = {_0, _831} + {_0, _2974};
  wire [1:0] _23247 = {_0, _5438} + {_0, _7965};
  wire [2:0] _23248 = {_0, _23246} + {_0, _23247};
  wire [1:0] _23249 = {_0, _9438} + {_0, _10783};
  wire [3:0] _23250 = {_0, _23248} + {_0, _0, _23249};
  wire _23251 = _12301 < _23250;
  wire _23252 = r831 ^ _23251;
  wire _23253 = _12298 ? coded_block[831] : r831;
  wire _23254 = _12296 ? _23252 : _23253;
  always @ (posedge reset or posedge clock) if (reset) r831 <= 1'd0; else if (_12300) r831 <= _23254;
  wire [1:0] _23255 = {_0, _192} + {_0, _3262};
  wire [1:0] _23256 = {_0, _5053} + {_0, _6303};
  wire [2:0] _23257 = {_0, _23255} + {_0, _23256};
  wire [1:0] _23258 = {_0, _8415} + {_0, _11259};
  wire [3:0] _23259 = {_0, _23257} + {_0, _0, _23258};
  wire _23260 = _12301 < _23259;
  wire _23261 = r830 ^ _23260;
  wire _23262 = _12298 ? coded_block[830] : r830;
  wire _23263 = _12296 ? _23261 : _23262;
  always @ (posedge reset or posedge clock) if (reset) r830 <= 1'd0; else if (_12300) r830 <= _23263;
  wire [1:0] _23264 = {_0, _863} + {_0, _2655};
  wire [1:0] _23265 = {_0, _5853} + {_0, _7675};
  wire [2:0] _23266 = {_0, _23264} + {_0, _23265};
  wire [1:0] _23267 = {_0, _8288} + {_0, _12282};
  wire [3:0] _23268 = {_0, _23266} + {_0, _0, _23267};
  wire _23269 = _12301 < _23268;
  wire _23270 = r829 ^ _23269;
  wire _23271 = _12298 ? coded_block[829] : r829;
  wire _23272 = _12296 ? _23270 : _23271;
  always @ (posedge reset or posedge clock) if (reset) r829 <= 1'd0; else if (_12300) r829 <= _23272;
  wire [1:0] _23273 = {_0, _894} + {_0, _2302};
  wire [1:0] _23274 = {_0, _4734} + {_0, _7931};
  wire [2:0] _23275 = {_0, _23273} + {_0, _23274};
  wire [1:0] _23276 = {_0, _9759} + {_0, _10366};
  wire [3:0] _23277 = {_0, _23275} + {_0, _0, _23276};
  wire _23278 = _12301 < _23277;
  wire _23279 = r828 ^ _23278;
  wire _23280 = _12298 ? coded_block[828] : r828;
  wire _23281 = _12296 ? _23279 : _23280;
  always @ (posedge reset or posedge clock) if (reset) r828 <= 1'd0; else if (_12300) r828 <= _23281;
  wire [1:0] _23282 = {_0, _927} + {_0, _2526};
  wire [1:0] _23283 = {_0, _4384} + {_0, _6814};
  wire [2:0] _23284 = {_0, _23282} + {_0, _23283};
  wire [1:0] _23285 = {_0, _10014} + {_0, _11837};
  wire [3:0] _23286 = {_0, _23284} + {_0, _0, _23285};
  wire _23287 = _12301 < _23286;
  wire _23288 = r827 ^ _23287;
  wire _23289 = _12298 ? coded_block[827] : r827;
  wire _23290 = _12296 ? _23288 : _23289;
  always @ (posedge reset or posedge clock) if (reset) r827 <= 1'd0; else if (_12300) r827 <= _23290;
  wire [1:0] _23291 = {_0, _1021} + {_0, _3486};
  wire [1:0] _23292 = {_0, _4830} + {_0, _6558};
  wire [2:0] _23293 = {_0, _23291} + {_0, _23292};
  wire [1:0] _23294 = {_0, _8767} + {_0, _10621};
  wire [3:0] _23295 = {_0, _23293} + {_0, _0, _23294};
  wire _23296 = _12301 < _23295;
  wire _23297 = r826 ^ _23296;
  wire _23298 = _12298 ? coded_block[826] : r826;
  wire _23299 = _12296 ? _23297 : _23298;
  always @ (posedge reset or posedge clock) if (reset) r826 <= 1'd0; else if (_12300) r826 <= _23299;
  wire [1:0] _23300 = {_0, _1057} + {_0, _4091};
  wire [1:0] _23301 = {_0, _5565} + {_0, _6908};
  wire [2:0] _23302 = {_0, _23300} + {_0, _23301};
  wire [1:0] _23303 = {_0, _8638} + {_0, _10846};
  wire [3:0] _23304 = {_0, _23302} + {_0, _0, _23303};
  wire _23305 = _12301 < _23304;
  wire _23306 = r825 ^ _23305;
  wire _23307 = _12298 ? coded_block[825] : r825;
  wire _23308 = _12296 ? _23306 : _23307;
  always @ (posedge reset or posedge clock) if (reset) r825 <= 1'd0; else if (_12300) r825 <= _23308;
  wire [1:0] _23309 = {_0, _1088} + {_0, _3646};
  wire [1:0] _23310 = {_0, _4160} + {_0, _7644};
  wire [2:0] _23311 = {_0, _23309} + {_0, _23310};
  wire [1:0] _23312 = {_0, _8991} + {_0, _10717};
  wire [3:0] _23313 = {_0, _23311} + {_0, _0, _23312};
  wire _23314 = _12301 < _23313;
  wire _23315 = r824 ^ _23314;
  wire _23316 = _12298 ? coded_block[824] : r824;
  wire _23317 = _12296 ? _23315 : _23316;
  always @ (posedge reset or posedge clock) if (reset) r824 <= 1'd0; else if (_12300) r824 <= _23317;
  wire [1:0] _23318 = {_0, _1120} + {_0, _3262};
  wire [1:0] _23319 = {_0, _5726} + {_0, _6239};
  wire [2:0] _23320 = {_0, _23318} + {_0, _23319};
  wire [1:0] _23321 = {_0, _9724} + {_0, _11069};
  wire [3:0] _23322 = {_0, _23320} + {_0, _0, _23321};
  wire _23323 = _12301 < _23322;
  wire _23324 = r823 ^ _23323;
  wire _23325 = _12298 ? coded_block[823] : r823;
  wire _23326 = _12296 ? _23324 : _23325;
  always @ (posedge reset or posedge clock) if (reset) r823 <= 1'd0; else if (_12300) r823 <= _23326;
  wire [1:0] _23327 = {_0, _1151} + {_0, _2271};
  wire [1:0] _23328 = {_0, _5342} + {_0, _7804};
  wire [2:0] _23329 = {_0, _23327} + {_0, _23328};
  wire [1:0] _23330 = {_0, _8319} + {_0, _11806};
  wire [3:0] _23331 = {_0, _23329} + {_0, _0, _23330};
  wire _23332 = _12301 < _23331;
  wire _23333 = r822 ^ _23332;
  wire _23334 = _12298 ? coded_block[822] : r822;
  wire _23335 = _12296 ? _23333 : _23334;
  always @ (posedge reset or posedge clock) if (reset) r822 <= 1'd0; else if (_12300) r822 <= _23335;
  wire [1:0] _23336 = {_0, _1184} + {_0, _2686};
  wire [1:0] _23337 = {_0, _4350} + {_0, _7420};
  wire [2:0] _23338 = {_0, _23336} + {_0, _23337};
  wire [1:0] _23339 = {_0, _9886} + {_0, _10399};
  wire [3:0] _23340 = {_0, _23338} + {_0, _0, _23339};
  wire _23341 = _12301 < _23340;
  wire _23342 = r821 ^ _23341;
  wire _23343 = _12298 ? coded_block[821] : r821;
  wire _23344 = _12296 ? _23342 : _23343;
  always @ (posedge reset or posedge clock) if (reset) r821 <= 1'd0; else if (_12300) r821 <= _23344;
  wire [1:0] _23345 = {_0, _1215} + {_0, _3167};
  wire [1:0] _23346 = {_0, _4767} + {_0, _6431};
  wire [2:0] _23347 = {_0, _23345} + {_0, _23346};
  wire [1:0] _23348 = {_0, _9503} + {_0, _11964};
  wire [3:0] _23349 = {_0, _23347} + {_0, _0, _23348};
  wire _23350 = _12301 < _23349;
  wire _23351 = r820 ^ _23350;
  wire _23352 = _12298 ? coded_block[820] : r820;
  wire _23353 = _12296 ? _23351 : _23352;
  always @ (posedge reset or posedge clock) if (reset) r820 <= 1'd0; else if (_12300) r820 <= _23353;
  wire [1:0] _23354 = {_0, _1278} + {_0, _3901};
  wire [1:0] _23355 = {_0, _4671} + {_0, _7326};
  wire [2:0] _23356 = {_0, _23354} + {_0, _23355};
  wire [1:0] _23357 = {_0, _8926} + {_0, _10590};
  wire [3:0] _23358 = {_0, _23356} + {_0, _0, _23357};
  wire _23359 = _12301 < _23358;
  wire _23360 = r819 ^ _23359;
  wire _23361 = _12298 ? coded_block[819] : r819;
  wire _23362 = _12296 ? _23360 : _23361;
  always @ (posedge reset or posedge clock) if (reset) r819 <= 1'd0; else if (_12300) r819 <= _23362;
  wire [1:0] _23363 = {_0, _1312} + {_0, _3580};
  wire [1:0] _23364 = {_0, _5981} + {_0, _6750};
  wire [2:0] _23365 = {_0, _23363} + {_0, _23364};
  wire [1:0] _23366 = {_0, _9406} + {_0, _11004};
  wire [3:0] _23367 = {_0, _23365} + {_0, _0, _23366};
  wire _23368 = _12301 < _23367;
  wire _23369 = r818 ^ _23368;
  wire _23370 = _12298 ? coded_block[818] : r818;
  wire _23371 = _12296 ? _23369 : _23370;
  always @ (posedge reset or posedge clock) if (reset) r818 <= 1'd0; else if (_12300) r818 <= _23371;
  wire [1:0] _23372 = {_0, _1343} + {_0, _3742};
  wire [1:0] _23373 = {_0, _5663} + {_0, _8059};
  wire [2:0] _23374 = {_0, _23372} + {_0, _23373};
  wire [1:0] _23375 = {_0, _8830} + {_0, _11485};
  wire [3:0] _23376 = {_0, _23374} + {_0, _0, _23375};
  wire _23377 = _12301 < _23376;
  wire _23378 = r817 ^ _23377;
  wire _23379 = _12298 ? coded_block[817] : r817;
  wire _23380 = _12296 ? _23378 : _23379;
  always @ (posedge reset or posedge clock) if (reset) r817 <= 1'd0; else if (_12300) r817 <= _23380;
  wire [1:0] _23381 = {_0, _1375} + {_0, _3549};
  wire [1:0] _23382 = {_0, _5821} + {_0, _7741};
  wire [2:0] _23383 = {_0, _23381} + {_0, _23382};
  wire [1:0] _23384 = {_0, _10141} + {_0, _10910};
  wire [3:0] _23385 = {_0, _23383} + {_0, _0, _23384};
  wire _23386 = _12301 < _23385;
  wire _23387 = r816 ^ _23386;
  wire _23388 = _12298 ? coded_block[816] : r816;
  wire _23389 = _12296 ? _23387 : _23388;
  always @ (posedge reset or posedge clock) if (reset) r816 <= 1'd0; else if (_12300) r816 <= _23389;
  wire [1:0] _23390 = {_0, _1406} + {_0, _3933};
  wire [1:0] _23391 = {_0, _5628} + {_0, _7900};
  wire [2:0] _23392 = {_0, _23390} + {_0, _23391};
  wire [1:0] _23393 = {_0, _9822} + {_0, _12219};
  wire [3:0] _23394 = {_0, _23392} + {_0, _0, _23393};
  wire _23395 = _12301 < _23394;
  wire _23396 = r815 ^ _23395;
  wire _23397 = _12298 ? coded_block[815] : r815;
  wire _23398 = _12296 ? _23396 : _23397;
  always @ (posedge reset or posedge clock) if (reset) r815 <= 1'd0; else if (_12300) r815 <= _23398;
  wire [1:0] _23399 = {_0, _1439} + {_0, _3068};
  wire [1:0] _23400 = {_0, _6012} + {_0, _7710};
  wire [2:0] _23401 = {_0, _23399} + {_0, _23400};
  wire [1:0] _23402 = {_0, _9980} + {_0, _11900};
  wire [3:0] _23403 = {_0, _23401} + {_0, _0, _23402};
  wire _23404 = _12301 < _23403;
  wire _23405 = r814 ^ _23404;
  wire _23406 = _12298 ? coded_block[814] : r814;
  wire _23407 = _12296 ? _23405 : _23406;
  always @ (posedge reset or posedge clock) if (reset) r814 <= 1'd0; else if (_12300) r814 <= _23407;
  wire [1:0] _23408 = {_0, _1470} + {_0, _2847};
  wire [1:0] _23409 = {_0, _5152} + {_0, _8092};
  wire [2:0] _23410 = {_0, _23408} + {_0, _23409};
  wire [1:0] _23411 = {_0, _9790} + {_0, _12061};
  wire [3:0] _23412 = {_0, _23410} + {_0, _0, _23411};
  wire _23413 = _12301 < _23412;
  wire _23414 = r813 ^ _23413;
  wire _23415 = _12298 ? coded_block[813] : r813;
  wire _23416 = _12296 ? _23414 : _23415;
  always @ (posedge reset or posedge clock) if (reset) r813 <= 1'd0; else if (_12300) r813 <= _23416;
  wire [1:0] _23417 = {_0, _1502} + {_0, _3422};
  wire [1:0] _23418 = {_0, _4926} + {_0, _7230};
  wire [2:0] _23419 = {_0, _23417} + {_0, _23418};
  wire [1:0] _23420 = {_0, _10172} + {_0, _11869};
  wire [3:0] _23421 = {_0, _23419} + {_0, _0, _23420};
  wire _23422 = _12301 < _23421;
  wire _23423 = r812 ^ _23422;
  wire _23424 = _12298 ? coded_block[812] : r812;
  wire _23425 = _12296 ? _23423 : _23424;
  always @ (posedge reset or posedge clock) if (reset) r812 <= 1'd0; else if (_12300) r812 <= _23425;
  wire [1:0] _23426 = {_0, _1533} + {_0, _3359};
  wire [1:0] _23427 = {_0, _5501} + {_0, _7005};
  wire [2:0] _23428 = {_0, _23426} + {_0, _23427};
  wire [1:0] _23429 = {_0, _9311} + {_0, _12251};
  wire [3:0] _23430 = {_0, _23428} + {_0, _0, _23429};
  wire _23431 = _12301 < _23430;
  wire _23432 = r811 ^ _23431;
  wire _23433 = _12298 ? coded_block[811] : r811;
  wire _23434 = _12296 ? _23432 : _23433;
  always @ (posedge reset or posedge clock) if (reset) r811 <= 1'd0; else if (_12300) r811 <= _23434;
  wire [1:0] _23435 = {_0, _1568} + {_0, _2463};
  wire [1:0] _23436 = {_0, _5438} + {_0, _7581};
  wire [2:0] _23437 = {_0, _23435} + {_0, _23436};
  wire [1:0] _23438 = {_0, _9085} + {_0, _11389};
  wire [3:0] _23439 = {_0, _23437} + {_0, _0, _23438};
  wire _23440 = _12301 < _23439;
  wire _23441 = r810 ^ _23440;
  wire _23442 = _12298 ? coded_block[810] : r810;
  wire _23443 = _12296 ? _23441 : _23442;
  always @ (posedge reset or posedge clock) if (reset) r810 <= 1'd0; else if (_12300) r810 <= _23443;
  wire [1:0] _23444 = {_0, _1599} + {_0, _3135};
  wire [1:0] _23445 = {_0, _4542} + {_0, _7517};
  wire [2:0] _23446 = {_0, _23444} + {_0, _23445};
  wire [1:0] _23447 = {_0, _9661} + {_0, _11165};
  wire [3:0] _23448 = {_0, _23446} + {_0, _0, _23447};
  wire _23449 = _12301 < _23448;
  wire _23450 = r809 ^ _23449;
  wire _23451 = _12298 ? coded_block[809] : r809;
  wire _23452 = _12296 ? _23450 : _23451;
  always @ (posedge reset or posedge clock) if (reset) r809 <= 1'd0; else if (_12300) r809 <= _23452;
  wire [1:0] _23453 = {_0, _1631} + {_0, _2719};
  wire [1:0] _23454 = {_0, _5215} + {_0, _6621};
  wire [2:0] _23455 = {_0, _23453} + {_0, _23454};
  wire [1:0] _23456 = {_0, _9597} + {_0, _11740};
  wire [3:0] _23457 = {_0, _23455} + {_0, _0, _23456};
  wire _23458 = _12301 < _23457;
  wire _23459 = r808 ^ _23458;
  wire _23460 = _12298 ? coded_block[808] : r808;
  wire _23461 = _12296 ? _23459 : _23460;
  always @ (posedge reset or posedge clock) if (reset) r808 <= 1'd0; else if (_12300) r808 <= _23461;
  wire [1:0] _23462 = {_0, _1662} + {_0, _2430};
  wire [1:0] _23463 = {_0, _4798} + {_0, _7293};
  wire [2:0] _23464 = {_0, _23462} + {_0, _23463};
  wire [1:0] _23465 = {_0, _8701} + {_0, _11677};
  wire [3:0] _23466 = {_0, _23464} + {_0, _0, _23465};
  wire _23467 = _12301 < _23466;
  wire _23468 = r807 ^ _23467;
  wire _23469 = _12298 ? coded_block[807] : r807;
  wire _23470 = _12296 ? _23468 : _23469;
  always @ (posedge reset or posedge clock) if (reset) r807 <= 1'd0; else if (_12300) r807 <= _23470;
  wire [1:0] _23471 = {_0, _1695} + {_0, _3390};
  wire [1:0] _23472 = {_0, _4511} + {_0, _6877};
  wire [2:0] _23473 = {_0, _23471} + {_0, _23472};
  wire [1:0] _23474 = {_0, _9375} + {_0, _10783};
  wire [3:0] _23475 = {_0, _23473} + {_0, _0, _23474};
  wire _23476 = _12301 < _23475;
  wire _23477 = r806 ^ _23476;
  wire _23478 = _12298 ? coded_block[806] : r806;
  wire _23479 = _12296 ? _23477 : _23478;
  always @ (posedge reset or posedge clock) if (reset) r806 <= 1'd0; else if (_12300) r806 <= _23479;
  wire [1:0] _23480 = {_0, _1758} + {_0, _3870};
  wire [1:0] _23481 = {_0, _4958} + {_0, _7548};
  wire [2:0] _23482 = {_0, _23480} + {_0, _23481};
  wire [1:0] _23483 = {_0, _8670} + {_0, _11038};
  wire [3:0] _23484 = {_0, _23482} + {_0, _0, _23483};
  wire _23485 = _12301 < _23484;
  wire _23486 = r805 ^ _23485;
  wire _23487 = _12298 ? coded_block[805] : r805;
  wire _23488 = _12296 ? _23486 : _23487;
  always @ (posedge reset or posedge clock) if (reset) r805 <= 1'd0; else if (_12300) r805 <= _23488;
  wire [1:0] _23489 = {_0, _1789} + {_0, _2623};
  wire [1:0] _23490 = {_0, _5949} + {_0, _7036};
  wire [2:0] _23491 = {_0, _23489} + {_0, _23490};
  wire [1:0] _23492 = {_0, _9630} + {_0, _10748};
  wire [3:0] _23493 = {_0, _23491} + {_0, _0, _23492};
  wire _23494 = _12301 < _23493;
  wire _23495 = r804 ^ _23494;
  wire _23496 = _12298 ? coded_block[804] : r804;
  wire _23497 = _12296 ? _23495 : _23496;
  always @ (posedge reset or posedge clock) if (reset) r804 <= 1'd0; else if (_12300) r804 <= _23497;
  wire [1:0] _23498 = {_0, _1823} + {_0, _3805};
  wire [1:0] _23499 = {_0, _4703} + {_0, _8028};
  wire [2:0] _23500 = {_0, _23498} + {_0, _23499};
  wire [1:0] _23501 = {_0, _9118} + {_0, _11708};
  wire [3:0] _23502 = {_0, _23500} + {_0, _0, _23501};
  wire _23503 = _12301 < _23502;
  wire _23504 = r803 ^ _23503;
  wire _23505 = _12298 ? coded_block[803] : r803;
  wire _23506 = _12296 ? _23504 : _23505;
  always @ (posedge reset or posedge clock) if (reset) r803 <= 1'd0; else if (_12300) r803 <= _23506;
  wire [1:0] _23507 = {_0, _1854} + {_0, _3325};
  wire [1:0] _23508 = {_0, _5884} + {_0, _6781};
  wire [2:0] _23509 = {_0, _23507} + {_0, _23508};
  wire [1:0] _23510 = {_0, _10108} + {_0, _11196};
  wire [3:0] _23511 = {_0, _23509} + {_0, _0, _23510};
  wire _23512 = _12301 < _23511;
  wire _23513 = r802 ^ _23512;
  wire _23514 = _12298 ? coded_block[802] : r802;
  wire _23515 = _12296 ? _23513 : _23514;
  always @ (posedge reset or posedge clock) if (reset) r802 <= 1'd0; else if (_12300) r802 <= _23515;
  wire [1:0] _23516 = {_0, _1886} + {_0, _3453};
  wire [1:0] _23517 = {_0, _5407} + {_0, _7965};
  wire [2:0] _23518 = {_0, _23516} + {_0, _23517};
  wire [1:0] _23519 = {_0, _8863} + {_0, _12188};
  wire [3:0] _23520 = {_0, _23518} + {_0, _0, _23519};
  wire _23521 = _12301 < _23520;
  wire _23522 = r801 ^ _23521;
  wire _23523 = _12298 ? coded_block[801] : r801;
  wire _23524 = _12296 ? _23522 : _23523;
  always @ (posedge reset or posedge clock) if (reset) r801 <= 1'd0; else if (_12300) r801 <= _23524;
  wire [1:0] _23525 = {_0, _1950} + {_0, _4028};
  wire [1:0] _23526 = {_0, _4861} + {_0, _7612};
  wire [2:0] _23527 = {_0, _23525} + {_0, _23526};
  wire [1:0] _23528 = {_0, _9566} + {_0, _12124};
  wire [3:0] _23529 = {_0, _23527} + {_0, _0, _23528};
  wire _23530 = _12301 < _23529;
  wire _23531 = r800 ^ _23530;
  wire _23532 = _12298 ? coded_block[800] : r800;
  wire _23533 = _12296 ? _23531 : _23532;
  always @ (posedge reset or posedge clock) if (reset) r800 <= 1'd0; else if (_12300) r800 <= _23533;
  wire [1:0] _23534 = {_0, _2013} + {_0, _2813};
  wire [1:0] _23535 = {_0, _6076} + {_0, _8186};
  wire [2:0] _23536 = {_0, _23534} + {_0, _23535};
  wire [1:0] _23537 = {_0, _9022} + {_0, _11771};
  wire [3:0] _23538 = {_0, _23536} + {_0, _0, _23537};
  wire _23539 = _12301 < _23538;
  wire _23540 = r799 ^ _23539;
  wire _23541 = _12298 ? coded_block[799] : r799;
  wire _23542 = _12296 ? _23540 : _23541;
  always @ (posedge reset or posedge clock) if (reset) r799 <= 1'd0; else if (_12300) r799 <= _23542;
  wire [1:0] _23543 = {_0, _2044} + {_0, _3104};
  wire [1:0] _23544 = {_0, _4895} + {_0, _8155};
  wire [2:0] _23545 = {_0, _23543} + {_0, _23544};
  wire [1:0] _23546 = {_0, _8256} + {_0, _11101};
  wire [3:0] _23547 = {_0, _23545} + {_0, _0, _23546};
  wire _23548 = _12301 < _23547;
  wire _23549 = r798 ^ _23548;
  wire _23550 = _12298 ? coded_block[798] : r798;
  wire _23551 = _12296 ? _23549 : _23550;
  always @ (posedge reset or posedge clock) if (reset) r798 <= 1'd0; else if (_12300) r798 <= _23551;
  wire [1:0] _23552 = {_0, _65} + {_0, _2494};
  wire [1:0] _23553 = {_0, _5183} + {_0, _6973};
  wire [2:0] _23554 = {_0, _23552} + {_0, _23553};
  wire [1:0] _23555 = {_0, _10235} + {_0, _10335};
  wire [3:0] _23556 = {_0, _23554} + {_0, _0, _23555};
  wire _23557 = _12301 < _23556;
  wire _23558 = r797 ^ _23557;
  wire _23559 = _12298 ? coded_block[797] : r797;
  wire _23560 = _12296 ? _23558 : _23559;
  always @ (posedge reset or posedge clock) if (reset) r797 <= 1'd0; else if (_12300) r797 <= _23560;
  wire [1:0] _23561 = {_0, _128} + {_0, _2081};
  wire [1:0] _23562 = {_0, _4415} + {_0, _6652};
  wire [2:0] _23563 = {_0, _23561} + {_0, _23562};
  wire [1:0] _23564 = {_0, _9342} + {_0, _11132};
  wire [3:0] _23565 = {_0, _23563} + {_0, _0, _23564};
  wire _23566 = _12301 < _23565;
  wire _23567 = r796 ^ _23566;
  wire _23568 = _12298 ? coded_block[796] : r796;
  wire _23569 = _12296 ? _23567 : _23568;
  always @ (posedge reset or posedge clock) if (reset) r796 <= 1'd0; else if (_12300) r796 <= _23569;
  wire [1:0] _23570 = {_0, _161} + {_0, _2367};
  wire [1:0] _23571 = {_0, _4129} + {_0, _6494};
  wire [2:0] _23572 = {_0, _23570} + {_0, _23571};
  wire [1:0] _23573 = {_0, _8736} + {_0, _11422};
  wire [3:0] _23574 = {_0, _23572} + {_0, _0, _23573};
  wire _23575 = _12301 < _23574;
  wire _23576 = r795 ^ _23575;
  wire _23577 = _12298 ? coded_block[795] : r795;
  wire _23578 = _12296 ? _23576 : _23577;
  always @ (posedge reset or posedge clock) if (reset) r795 <= 1'd0; else if (_12300) r795 <= _23578;
  wire [1:0] _23579 = {_0, _192} + {_0, _2557};
  wire [1:0] _23580 = {_0, _4447} + {_0, _6176};
  wire [2:0] _23581 = {_0, _23579} + {_0, _23580};
  wire [1:0] _23582 = {_0, _8574} + {_0, _10814};
  wire [3:0] _23583 = {_0, _23581} + {_0, _0, _23582};
  wire _23584 = _12301 < _23583;
  wire _23585 = r794 ^ _23584;
  wire _23586 = _12298 ? coded_block[794] : r794;
  wire _23587 = _12296 ? _23585 : _23586;
  always @ (posedge reset or posedge clock) if (reset) r794 <= 1'd0; else if (_12300) r794 <= _23587;
  wire [1:0] _23588 = {_0, _224} + {_0, _3198};
  wire [1:0] _23589 = {_0, _4640} + {_0, _6525};
  wire [2:0] _23590 = {_0, _23588} + {_0, _23589};
  wire [1:0] _23591 = {_0, _8225} + {_0, _10654};
  wire [3:0] _23592 = {_0, _23590} + {_0, _0, _23591};
  wire _23593 = _12301 < _23592;
  wire _23594 = r793 ^ _23593;
  wire _23595 = _12298 ? coded_block[793] : r793;
  wire _23596 = _12296 ? _23594 : _23595;
  always @ (posedge reset or posedge clock) if (reset) r793 <= 1'd0; else if (_12300) r793 <= _23596;
  wire [1:0] _23597 = {_0, _255} + {_0, _2941};
  wire [1:0] _23598 = {_0, _5279} + {_0, _6718};
  wire [2:0] _23599 = {_0, _23597} + {_0, _23598};
  wire [1:0] _23600 = {_0, _8607} + {_0, _10272};
  wire [3:0] _23601 = {_0, _23599} + {_0, _0, _23600};
  wire _23602 = _12301 < _23601;
  wire _23603 = r792 ^ _23602;
  wire _23604 = _12298 ? coded_block[792] : r792;
  wire _23605 = _12296 ? _23603 : _23604;
  always @ (posedge reset or posedge clock) if (reset) r792 <= 1'd0; else if (_12300) r792 <= _23605;
  wire [1:0] _23606 = {_0, _320} + {_0, _2208};
  wire [1:0] _23607 = {_0, _4223} + {_0, _7100};
  wire [2:0] _23608 = {_0, _23606} + {_0, _23607};
  wire [1:0] _23609 = {_0, _9438} + {_0, _10877};
  wire [3:0] _23610 = {_0, _23608} + {_0, _0, _23609};
  wire _23611 = _12301 < _23610;
  wire _23612 = r791 ^ _23611;
  wire _23613 = _12298 ? coded_block[791] : r791;
  wire _23614 = _12296 ? _23612 : _23613;
  always @ (posedge reset or posedge clock) if (reset) r791 <= 1'd0; else if (_12300) r791 <= _23614;
  wire [1:0] _23615 = {_0, _352} + {_0, _3005};
  wire [1:0] _23616 = {_0, _4287} + {_0, _6303};
  wire [2:0] _23617 = {_0, _23615} + {_0, _23616};
  wire [1:0] _23618 = {_0, _9181} + {_0, _11516};
  wire [3:0] _23619 = {_0, _23617} + {_0, _0, _23618};
  wire _23620 = _12301 < _23619;
  wire _23621 = r790 ^ _23620;
  wire _23622 = _12298 ? coded_block[790] : r790;
  wire _23623 = _12296 ? _23621 : _23622;
  always @ (posedge reset or posedge clock) if (reset) r790 <= 1'd0; else if (_12300) r790 <= _23623;
  wire [1:0] _23624 = {_0, _383} + {_0, _3709};
  wire [1:0] _23625 = {_0, _5085} + {_0, _6366};
  wire [2:0] _23626 = {_0, _23624} + {_0, _23625};
  wire [1:0] _23627 = {_0, _8383} + {_0, _11259};
  wire [3:0] _23628 = {_0, _23626} + {_0, _0, _23627};
  wire _23629 = _12301 < _23628;
  wire _23630 = r789 ^ _23629;
  wire _23631 = _12298 ? coded_block[789] : r789;
  wire _23632 = _12296 ? _23630 : _23631;
  always @ (posedge reset or posedge clock) if (reset) r789 <= 1'd0; else if (_12300) r789 <= _23632;
  wire [1:0] _23633 = {_0, _416} + {_0, _3615};
  wire [1:0] _23634 = {_0, _5790} + {_0, _7163};
  wire [2:0] _23635 = {_0, _23633} + {_0, _23634};
  wire [1:0] _23636 = {_0, _8446} + {_0, _10462};
  wire [3:0] _23637 = {_0, _23635} + {_0, _0, _23636};
  wire _23638 = _12301 < _23637;
  wire _23639 = r788 ^ _23638;
  wire _23640 = _12298 ? coded_block[788] : r788;
  wire _23641 = _12296 ? _23639 : _23640;
  always @ (posedge reset or posedge clock) if (reset) r788 <= 1'd0; else if (_12300) r788 <= _23641;
  wire [1:0] _23642 = {_0, _447} + {_0, _2112};
  wire [1:0] _23643 = {_0, _5694} + {_0, _7868};
  wire [2:0] _23644 = {_0, _23642} + {_0, _23643};
  wire [1:0] _23645 = {_0, _9248} + {_0, _10527};
  wire [3:0] _23646 = {_0, _23644} + {_0, _0, _23645};
  wire _23647 = _12301 < _23646;
  wire _23648 = r787 ^ _23647;
  wire _23649 = _12298 ? coded_block[787] : r787;
  wire _23650 = _12296 ? _23648 : _23649;
  always @ (posedge reset or posedge clock) if (reset) r787 <= 1'd0; else if (_12300) r787 <= _23650;
  wire [1:0] _23651 = {_0, _479} + {_0, _2974};
  wire [1:0] _23652 = {_0, _4192} + {_0, _7773};
  wire [2:0] _23653 = {_0, _23651} + {_0, _23652};
  wire [1:0] _23654 = {_0, _9949} + {_0, _11326};
  wire [3:0] _23655 = {_0, _23653} + {_0, _0, _23654};
  wire _23656 = _12301 < _23655;
  wire _23657 = r786 ^ _23656;
  wire _23658 = _12298 ? coded_block[786] : r786;
  wire _23659 = _12296 ? _23657 : _23658;
  always @ (posedge reset or posedge clock) if (reset) r786 <= 1'd0; else if (_12300) r786 <= _23659;
  wire [1:0] _23660 = {_0, _510} + {_0, _2239};
  wire [1:0] _23661 = {_0, _5053} + {_0, _6270};
  wire [2:0] _23662 = {_0, _23660} + {_0, _23661};
  wire [1:0] _23663 = {_0, _9853} + {_0, _12027};
  wire [3:0] _23664 = {_0, _23662} + {_0, _0, _23663};
  wire _23665 = _12301 < _23664;
  wire _23666 = r785 ^ _23665;
  wire _23667 = _12298 ? coded_block[785] : r785;
  wire _23668 = _12296 ? _23666 : _23667;
  always @ (posedge reset or posedge clock) if (reset) r785 <= 1'd0; else if (_12300) r785 <= _23668;
  wire [1:0] _23669 = {_0, _576} + {_0, _3836};
  wire [1:0] _23670 = {_0, _5373} + {_0, _6397};
  wire [2:0] _23671 = {_0, _23669} + {_0, _23670};
  wire [1:0] _23672 = {_0, _9212} + {_0, _10430};
  wire [3:0] _23673 = {_0, _23671} + {_0, _0, _23672};
  wire _23674 = _12301 < _23673;
  wire _23675 = r784 ^ _23674;
  wire _23676 = _12298 ? coded_block[784] : r784;
  wire _23677 = _12296 ? _23675 : _23676;
  always @ (posedge reset or posedge clock) if (reset) r784 <= 1'd0; else if (_12300) r784 <= _23677;
  wire [1:0] _23678 = {_0, _608} + {_0, _2910};
  wire [1:0] _23679 = {_0, _5918} + {_0, _7454};
  wire [2:0] _23680 = {_0, _23678} + {_0, _23679};
  wire [1:0] _23681 = {_0, _8480} + {_0, _11295};
  wire [3:0] _23682 = {_0, _23680} + {_0, _0, _23681};
  wire _23683 = _12301 < _23682;
  wire _23684 = r783 ^ _23683;
  wire _23685 = _12298 ? coded_block[783] : r783;
  wire _23686 = _12296 ? _23684 : _23685;
  always @ (posedge reset or posedge clock) if (reset) r783 <= 1'd0; else if (_12300) r783 <= _23686;
  wire [1:0] _23687 = {_0, _639} + {_0, _3231};
  wire [1:0] _23688 = {_0, _4989} + {_0, _7996};
  wire [2:0] _23689 = {_0, _23687} + {_0, _23688};
  wire [1:0] _23690 = {_0, _9534} + {_0, _10558};
  wire [3:0] _23691 = {_0, _23689} + {_0, _0, _23690};
  wire _23692 = _12301 < _23691;
  wire _23693 = r782 ^ _23692;
  wire _23694 = _12298 ? coded_block[782] : r782;
  wire _23695 = _12296 ? _23693 : _23694;
  always @ (posedge reset or posedge clock) if (reset) r782 <= 1'd0; else if (_12300) r782 <= _23695;
  wire [1:0] _23696 = {_0, _672} + {_0, _3678};
  wire [1:0] _23697 = {_0, _5310} + {_0, _7069};
  wire [2:0] _23698 = {_0, _23696} + {_0, _23697};
  wire [1:0] _23699 = {_0, _10077} + {_0, _11613};
  wire [3:0] _23700 = {_0, _23698} + {_0, _0, _23699};
  wire _23701 = _12301 < _23700;
  wire _23702 = r781 ^ _23701;
  wire _23703 = _12298 ? coded_block[781] : r781;
  wire _23704 = _12296 ? _23702 : _23703;
  always @ (posedge reset or posedge clock) if (reset) r781 <= 1'd0; else if (_12300) r781 <= _23704;
  wire [1:0] _23705 = {_0, _703} + {_0, _3037};
  wire [1:0] _23706 = {_0, _5757} + {_0, _7389};
  wire [2:0] _23707 = {_0, _23705} + {_0, _23706};
  wire [1:0] _23708 = {_0, _9149} + {_0, _12155};
  wire [3:0] _23709 = {_0, _23707} + {_0, _0, _23708};
  wire _23710 = _12301 < _23709;
  wire _23711 = r780 ^ _23710;
  wire _23712 = _12298 ? coded_block[780] : r780;
  wire _23713 = _12296 ? _23711 : _23712;
  always @ (posedge reset or posedge clock) if (reset) r780 <= 1'd0; else if (_12300) r780 <= _23713;
  wire [1:0] _23714 = {_0, _766} + {_0, _4060};
  wire [1:0] _23715 = {_0, _6045} + {_0, _7199};
  wire [2:0] _23716 = {_0, _23714} + {_0, _23715};
  wire [1:0] _23717 = {_0, _9917} + {_0, _11550};
  wire [3:0] _23718 = {_0, _23716} + {_0, _0, _23717};
  wire _23719 = _12301 < _23718;
  wire _23720 = r779 ^ _23719;
  wire _23721 = _12298 ? coded_block[779] : r779;
  wire _23722 = _12296 ? _23720 : _23721;
  always @ (posedge reset or posedge clock) if (reset) r779 <= 1'd0; else if (_12300) r779 <= _23722;
  wire [1:0] _23723 = {_0, _800} + {_0, _3517};
  wire [1:0] _23724 = {_0, _6139} + {_0, _8123};
  wire [2:0] _23725 = {_0, _23723} + {_0, _23724};
  wire [1:0] _23726 = {_0, _9279} + {_0, _11996};
  wire [3:0] _23727 = {_0, _23725} + {_0, _0, _23726};
  wire _23728 = _12301 < _23727;
  wire _23729 = r778 ^ _23728;
  wire _23730 = _12298 ? coded_block[778] : r778;
  wire _23731 = _12296 ? _23729 : _23730;
  always @ (posedge reset or posedge clock) if (reset) r778 <= 1'd0; else if (_12300) r778 <= _23731;
  wire [1:0] _23732 = {_0, _224} + {_0, _2655};
  wire [1:0] _23733 = {_0, _5342} + {_0, _7132};
  wire [2:0] _23734 = {_0, _23732} + {_0, _23733};
  wire [1:0] _23735 = {_0, _8383} + {_0, _10493};
  wire [3:0] _23736 = {_0, _23734} + {_0, _0, _23735};
  wire _23737 = _12301 < _23736;
  wire _23738 = r777 ^ _23737;
  wire _23739 = _12298 ? coded_block[777] : r777;
  wire _23740 = _12296 ? _23738 : _23739;
  always @ (posedge reset or posedge clock) if (reset) r777 <= 1'd0; else if (_12300) r777 <= _23740;
  wire [1:0] _23741 = {_0, _1502} + {_0, _3037};
  wire [1:0] _23742 = {_0, _4447} + {_0, _7420};
  wire [2:0] _23743 = {_0, _23741} + {_0, _23742};
  wire [1:0] _23744 = {_0, _9566} + {_0, _11069};
  wire [3:0] _23745 = {_0, _23743} + {_0, _0, _23744};
  wire _23746 = _12301 < _23745;
  wire _23747 = r776 ^ _23746;
  wire _23748 = _12298 ? coded_block[776] : r776;
  wire _23749 = _12296 ? _23747 : _23748;
  always @ (posedge reset or posedge clock) if (reset) r776 <= 1'd0; else if (_12300) r776 <= _23749;
  wire [1:0] _23750 = {_0, _1568} + {_0, _2336};
  wire [1:0] _23751 = {_0, _4703} + {_0, _7199};
  wire [2:0] _23752 = {_0, _23750} + {_0, _23751};
  wire [1:0] _23753 = {_0, _8607} + {_0, _11581};
  wire [3:0] _23754 = {_0, _23752} + {_0, _0, _23753};
  wire _23755 = _12301 < _23754;
  wire _23756 = r775 ^ _23755;
  wire _23757 = _12298 ? coded_block[775] : r775;
  wire _23758 = _12296 ? _23756 : _23757;
  always @ (posedge reset or posedge clock) if (reset) r775 <= 1'd0; else if (_12300) r775 <= _23758;
  wire [1:0] _23759 = {_0, _1599} + {_0, _3294};
  wire [1:0] _23760 = {_0, _4415} + {_0, _6781};
  wire [2:0] _23761 = {_0, _23759} + {_0, _23760};
  wire [1:0] _23762 = {_0, _9279} + {_0, _10685};
  wire [3:0] _23763 = {_0, _23761} + {_0, _0, _23762};
  wire _23764 = _12301 < _23763;
  wire _23765 = r774 ^ _23764;
  wire _23766 = _12298 ? coded_block[774] : r774;
  wire _23767 = _12296 ? _23765 : _23766;
  always @ (posedge reset or posedge clock) if (reset) r774 <= 1'd0; else if (_12300) r774 <= _23767;
  wire [1:0] _23768 = {_0, _1631} + {_0, _2782};
  wire [1:0] _23769 = {_0, _5373} + {_0, _6494};
  wire [2:0] _23770 = {_0, _23768} + {_0, _23769};
  wire [1:0] _23771 = {_0, _8863} + {_0, _11358};
  wire [3:0] _23772 = {_0, _23770} + {_0, _0, _23771};
  wire _23773 = _12301 < _23772;
  wire _23774 = r773 ^ _23773;
  wire _23775 = _12298 ? coded_block[773] : r773;
  wire _23776 = _12296 ? _23774 : _23775;
  always @ (posedge reset or posedge clock) if (reset) r773 <= 1'd0; else if (_12300) r773 <= _23776;
  wire [1:0] _23777 = {_0, _1695} + {_0, _2526};
  wire [1:0] _23778 = {_0, _5853} + {_0, _6942};
  wire [2:0] _23779 = {_0, _23777} + {_0, _23778};
  wire [1:0] _23780 = {_0, _9534} + {_0, _10654};
  wire [3:0] _23781 = {_0, _23779} + {_0, _0, _23780};
  wire _23782 = _12301 < _23781;
  wire _23783 = r772 ^ _23782;
  wire _23784 = _12298 ? coded_block[772] : r772;
  wire _23785 = _12296 ? _23783 : _23784;
  always @ (posedge reset or posedge clock) if (reset) r772 <= 1'd0; else if (_12300) r772 <= _23785;
  wire [1:0] _23786 = {_0, _1726} + {_0, _3709};
  wire [1:0] _23787 = {_0, _4605} + {_0, _7931};
  wire [2:0] _23788 = {_0, _23786} + {_0, _23787};
  wire [1:0] _23789 = {_0, _9022} + {_0, _11613};
  wire [3:0] _23790 = {_0, _23788} + {_0, _0, _23789};
  wire _23791 = _12301 < _23790;
  wire _23792 = r771 ^ _23791;
  wire _23793 = _12298 ? coded_block[771] : r771;
  wire _23794 = _12296 ? _23792 : _23793;
  always @ (posedge reset or posedge clock) if (reset) r771 <= 1'd0; else if (_12300) r771 <= _23794;
  wire [1:0] _23795 = {_0, _1758} + {_0, _3231};
  wire [1:0] _23796 = {_0, _5790} + {_0, _6687};
  wire [2:0] _23797 = {_0, _23795} + {_0, _23796};
  wire [1:0] _23798 = {_0, _10014} + {_0, _11101};
  wire [3:0] _23799 = {_0, _23797} + {_0, _0, _23798};
  wire _23800 = _12301 < _23799;
  wire _23801 = r770 ^ _23800;
  wire _23802 = _12298 ? coded_block[770] : r770;
  wire _23803 = _12296 ? _23801 : _23802;
  always @ (posedge reset or posedge clock) if (reset) r770 <= 1'd0; else if (_12300) r770 <= _23803;
  wire [1:0] _23804 = {_0, _1789} + {_0, _3359};
  wire [1:0] _23805 = {_0, _5310} + {_0, _7868};
  wire [2:0] _23806 = {_0, _23804} + {_0, _23805};
  wire [1:0] _23807 = {_0, _8767} + {_0, _12092};
  wire [3:0] _23808 = {_0, _23806} + {_0, _0, _23807};
  wire _23809 = _12301 < _23808;
  wire _23810 = r769 ^ _23809;
  wire _23811 = _12298 ? coded_block[769] : r769;
  wire _23812 = _12296 ? _23810 : _23811;
  always @ (posedge reset or posedge clock) if (reset) r769 <= 1'd0; else if (_12300) r769 <= _23812;
  wire [1:0] _23813 = {_0, _1854} + {_0, _3933};
  wire [1:0] _23814 = {_0, _4767} + {_0, _7517};
  wire [2:0] _23815 = {_0, _23813} + {_0, _23814};
  wire [1:0] _23816 = {_0, _9469} + {_0, _12027};
  wire [3:0] _23817 = {_0, _23815} + {_0, _0, _23816};
  wire _23818 = _12301 < _23817;
  wire _23819 = r768 ^ _23818;
  wire _23820 = _12298 ? coded_block[768] : r768;
  wire _23821 = _12296 ? _23819 : _23820;
  always @ (posedge reset or posedge clock) if (reset) r768 <= 1'd0; else if (_12300) r768 <= _23821;
  wire [1:0] _23822 = {_0, _1886} + {_0, _3901};
  wire [1:0] _23823 = {_0, _6012} + {_0, _6845};
  wire [2:0] _23824 = {_0, _23822} + {_0, _23823};
  wire [1:0] _23825 = {_0, _9597} + {_0, _11550};
  wire [3:0] _23826 = {_0, _23824} + {_0, _0, _23825};
  wire _23827 = _12301 < _23826;
  wire _23828 = r767 ^ _23827;
  wire _23829 = _12298 ? coded_block[767] : r767;
  wire _23830 = _12296 ? _23828 : _23829;
  always @ (posedge reset or posedge clock) if (reset) r767 <= 1'd0; else if (_12300) r767 <= _23830;
  wire [1:0] _23831 = {_0, _1917} + {_0, _2719};
  wire [1:0] _23832 = {_0, _5981} + {_0, _8092};
  wire [2:0] _23833 = {_0, _23831} + {_0, _23832};
  wire [1:0] _23834 = {_0, _8926} + {_0, _11677};
  wire [3:0] _23835 = {_0, _23833} + {_0, _0, _23834};
  wire _23836 = _12301 < _23835;
  wire _23837 = r766 ^ _23836;
  wire _23838 = _12298 ? coded_block[766] : r766;
  wire _23839 = _12296 ? _23837 : _23838;
  always @ (posedge reset or posedge clock) if (reset) r766 <= 1'd0; else if (_12300) r766 <= _23839;
  wire [1:0] _23840 = {_0, _1950} + {_0, _3005};
  wire [1:0] _23841 = {_0, _4798} + {_0, _8059};
  wire [2:0] _23842 = {_0, _23840} + {_0, _23841};
  wire [1:0] _23843 = {_0, _10172} + {_0, _11004};
  wire [3:0] _23844 = {_0, _23842} + {_0, _0, _23843};
  wire _23845 = _12301 < _23844;
  wire _23846 = r765 ^ _23845;
  wire _23847 = _12298 ? coded_block[765] : r765;
  wire _23848 = _12296 ? _23846 : _23847;
  always @ (posedge reset or posedge clock) if (reset) r765 <= 1'd0; else if (_12300) r765 <= _23848;
  wire [1:0] _23849 = {_0, _1981} + {_0, _2399};
  wire [1:0] _23850 = {_0, _5085} + {_0, _6877};
  wire [2:0] _23851 = {_0, _23849} + {_0, _23850};
  wire [1:0] _23852 = {_0, _10141} + {_0, _12251};
  wire [3:0] _23853 = {_0, _23851} + {_0, _0, _23852};
  wire _23854 = _12301 < _23853;
  wire _23855 = r764 ^ _23854;
  wire _23856 = _12298 ? coded_block[764] : r764;
  wire _23857 = _12296 ? _23855 : _23856;
  always @ (posedge reset or posedge clock) if (reset) r764 <= 1'd0; else if (_12300) r764 <= _23857;
  wire [1:0] _23858 = {_0, _2044} + {_0, _2081};
  wire [1:0] _23859 = {_0, _4319} + {_0, _6558};
  wire [2:0] _23860 = {_0, _23858} + {_0, _23859};
  wire [1:0] _23861 = {_0, _9248} + {_0, _11038};
  wire [3:0] _23862 = {_0, _23860} + {_0, _0, _23861};
  wire _23863 = _12301 < _23862;
  wire _23864 = r763 ^ _23863;
  wire _23865 = _12298 ? coded_block[763] : r763;
  wire _23866 = _12296 ? _23864 : _23865;
  always @ (posedge reset or posedge clock) if (reset) r763 <= 1'd0; else if (_12300) r763 <= _23866;
  wire [1:0] _23867 = {_0, _65} + {_0, _2271};
  wire [1:0] _23868 = {_0, _4129} + {_0, _6397};
  wire [2:0] _23869 = {_0, _23867} + {_0, _23868};
  wire [1:0] _23870 = {_0, _8638} + {_0, _11326};
  wire [3:0] _23871 = {_0, _23869} + {_0, _0, _23870};
  wire _23872 = _12301 < _23871;
  wire _23873 = r762 ^ _23872;
  wire _23874 = _12298 ? coded_block[762] : r762;
  wire _23875 = _12296 ? _23873 : _23874;
  always @ (posedge reset or posedge clock) if (reset) r762 <= 1'd0; else if (_12300) r762 <= _23875;
  wire [1:0] _23876 = {_0, _97} + {_0, _2463};
  wire [1:0] _23877 = {_0, _4350} + {_0, _6176};
  wire [2:0] _23878 = {_0, _23876} + {_0, _23877};
  wire [1:0] _23879 = {_0, _8480} + {_0, _10717};
  wire [3:0] _23880 = {_0, _23878} + {_0, _0, _23879};
  wire _23881 = _12301 < _23880;
  wire _23882 = r761 ^ _23881;
  wire _23883 = _12298 ? coded_block[761] : r761;
  wire _23884 = _12296 ? _23882 : _23883;
  always @ (posedge reset or posedge clock) if (reset) r761 <= 1'd0; else if (_12300) r761 <= _23884;
  wire [1:0] _23885 = {_0, _128} + {_0, _3104};
  wire [1:0] _23886 = {_0, _4542} + {_0, _6431};
  wire [2:0] _23887 = {_0, _23885} + {_0, _23886};
  wire [1:0] _23888 = {_0, _8225} + {_0, _10558};
  wire [3:0] _23889 = {_0, _23887} + {_0, _0, _23888};
  wire _23890 = _12301 < _23889;
  wire _23891 = r760 ^ _23890;
  wire _23892 = _12298 ? coded_block[760] : r760;
  wire _23893 = _12296 ? _23891 : _23892;
  always @ (posedge reset or posedge clock) if (reset) r760 <= 1'd0; else if (_12300) r760 <= _23893;
  wire [1:0] _23894 = {_0, _161} + {_0, _2847};
  wire [1:0] _23895 = {_0, _5183} + {_0, _6621};
  wire [2:0] _23896 = {_0, _23894} + {_0, _23895};
  wire [1:0] _23897 = {_0, _8511} + {_0, _10272};
  wire [3:0] _23898 = {_0, _23896} + {_0, _0, _23897};
  wire _23899 = _12301 < _23898;
  wire _23900 = r759 ^ _23899;
  wire _23901 = _12298 ? coded_block[759] : r759;
  wire _23902 = _12296 ? _23900 : _23901;
  always @ (posedge reset or posedge clock) if (reset) r759 <= 1'd0; else if (_12300) r759 <= _23902;
  wire [1:0] _23903 = {_0, _192} + {_0, _4060};
  wire [1:0] _23904 = {_0, _4926} + {_0, _7262};
  wire [2:0] _23905 = {_0, _23903} + {_0, _23904};
  wire [1:0] _23906 = {_0, _8701} + {_0, _10590};
  wire [3:0] _23907 = {_0, _23905} + {_0, _0, _23906};
  wire _23908 = _12301 < _23907;
  wire _23909 = r758 ^ _23908;
  wire _23910 = _12298 ? coded_block[758] : r758;
  wire _23911 = _12296 ? _23909 : _23910;
  always @ (posedge reset or posedge clock) if (reset) r758 <= 1'd0; else if (_12300) r758 <= _23911;
  wire [1:0] _23912 = {_0, _224} + {_0, _2112};
  wire [1:0] _23913 = {_0, _6139} + {_0, _7005};
  wire [2:0] _23914 = {_0, _23912} + {_0, _23913};
  wire [1:0] _23915 = {_0, _9342} + {_0, _10783};
  wire [3:0] _23916 = {_0, _23914} + {_0, _0, _23915};
  wire _23917 = _12301 < _23916;
  wire _23918 = r757 ^ _23917;
  wire _23919 = _12298 ? coded_block[757] : r757;
  wire _23920 = _12296 ? _23918 : _23919;
  always @ (posedge reset or posedge clock) if (reset) r757 <= 1'd0; else if (_12300) r757 <= _23920;
  wire [1:0] _23921 = {_0, _255} + {_0, _2910};
  wire [1:0] _23922 = {_0, _4192} + {_0, _6207};
  wire [2:0] _23923 = {_0, _23921} + {_0, _23922};
  wire [1:0] _23924 = {_0, _9085} + {_0, _11422};
  wire [3:0] _23925 = {_0, _23923} + {_0, _0, _23924};
  wire _23926 = _12301 < _23925;
  wire _23927 = r756 ^ _23926;
  wire _23928 = _12298 ? coded_block[756] : r756;
  wire _23929 = _12296 ? _23927 : _23928;
  always @ (posedge reset or posedge clock) if (reset) r756 <= 1'd0; else if (_12300) r756 <= _23929;
  wire [1:0] _23930 = {_0, _289} + {_0, _3615};
  wire [1:0] _23931 = {_0, _4989} + {_0, _6270};
  wire [2:0] _23932 = {_0, _23930} + {_0, _23931};
  wire [1:0] _23933 = {_0, _8288} + {_0, _11165};
  wire [3:0] _23934 = {_0, _23932} + {_0, _0, _23933};
  wire _23935 = _12301 < _23934;
  wire _23936 = r755 ^ _23935;
  wire _23937 = _12298 ? coded_block[755] : r755;
  wire _23938 = _12296 ? _23936 : _23937;
  always @ (posedge reset or posedge clock) if (reset) r755 <= 1'd0; else if (_12300) r755 <= _23938;
  wire [1:0] _23939 = {_0, _320} + {_0, _3517};
  wire [1:0] _23940 = {_0, _5694} + {_0, _7069};
  wire [2:0] _23941 = {_0, _23939} + {_0, _23940};
  wire [1:0] _23942 = {_0, _8352} + {_0, _10366};
  wire [3:0] _23943 = {_0, _23941} + {_0, _0, _23942};
  wire _23944 = _12301 < _23943;
  wire _23945 = r754 ^ _23944;
  wire _23946 = _12298 ? coded_block[754] : r754;
  wire _23947 = _12296 ? _23945 : _23946;
  always @ (posedge reset or posedge clock) if (reset) r754 <= 1'd0; else if (_12300) r754 <= _23947;
  wire [1:0] _23948 = {_0, _352} + {_0, _4028};
  wire [1:0] _23949 = {_0, _5597} + {_0, _7773};
  wire [2:0] _23950 = {_0, _23948} + {_0, _23949};
  wire [1:0] _23951 = {_0, _9149} + {_0, _10430};
  wire [3:0] _23952 = {_0, _23950} + {_0, _0, _23951};
  wire _23953 = _12301 < _23952;
  wire _23954 = r753 ^ _23953;
  wire _23955 = _12298 ? coded_block[753] : r753;
  wire _23956 = _12296 ? _23954 : _23955;
  always @ (posedge reset or posedge clock) if (reset) r753 <= 1'd0; else if (_12300) r753 <= _23956;
  wire [1:0] _23957 = {_0, _383} + {_0, _2878};
  wire [1:0] _23958 = {_0, _6108} + {_0, _7675};
  wire [2:0] _23959 = {_0, _23957} + {_0, _23958};
  wire [1:0] _23960 = {_0, _9853} + {_0, _11228};
  wire [3:0] _23961 = {_0, _23959} + {_0, _0, _23960};
  wire _23962 = _12301 < _23961;
  wire _23963 = r752 ^ _23962;
  wire _23964 = _12298 ? coded_block[752] : r752;
  wire _23965 = _12296 ? _23963 : _23964;
  always @ (posedge reset or posedge clock) if (reset) r752 <= 1'd0; else if (_12300) r752 <= _23965;
  wire [1:0] _23966 = {_0, _416} + {_0, _2144};
  wire [1:0] _23967 = {_0, _4958} + {_0, _8186};
  wire [2:0] _23968 = {_0, _23966} + {_0, _23967};
  wire [1:0] _23969 = {_0, _9759} + {_0, _11933};
  wire [3:0] _23970 = {_0, _23968} + {_0, _0, _23969};
  wire _23971 = _12301 < _23970;
  wire _23972 = r751 ^ _23971;
  wire _23973 = _12298 ? coded_block[751] : r751;
  wire _23974 = _12296 ? _23972 : _23973;
  always @ (posedge reset or posedge clock) if (reset) r751 <= 1'd0; else if (_12300) r751 <= _23974;
  wire [1:0] _23975 = {_0, _447} + {_0, _3198};
  wire [1:0] _23976 = {_0, _4223} + {_0, _7036};
  wire [2:0] _23977 = {_0, _23975} + {_0, _23976};
  wire [1:0] _23978 = {_0, _8256} + {_0, _11837};
  wire [3:0] _23979 = {_0, _23977} + {_0, _0, _23978};
  wire _23980 = _12301 < _23979;
  wire _23981 = r750 ^ _23980;
  wire _23982 = _12298 ? coded_block[750] : r750;
  wire _23983 = _12296 ? _23981 : _23982;
  always @ (posedge reset or posedge clock) if (reset) r750 <= 1'd0; else if (_12300) r750 <= _23983;
  wire [1:0] _23984 = {_0, _479} + {_0, _3742};
  wire [1:0] _23985 = {_0, _5279} + {_0, _6303};
  wire [2:0] _23986 = {_0, _23984} + {_0, _23985};
  wire [1:0] _23987 = {_0, _9118} + {_0, _10335};
  wire [3:0] _23988 = {_0, _23986} + {_0, _0, _23987};
  wire _23989 = _12301 < _23988;
  wire _23990 = r749 ^ _23989;
  wire _23991 = _12298 ? coded_block[749] : r749;
  wire _23992 = _12296 ? _23990 : _23991;
  always @ (posedge reset or posedge clock) if (reset) r749 <= 1'd0; else if (_12300) r749 <= _23992;
  wire [1:0] _23993 = {_0, _545} + {_0, _3135};
  wire [1:0] _23994 = {_0, _4895} + {_0, _7900};
  wire [2:0] _23995 = {_0, _23993} + {_0, _23994};
  wire [1:0] _23996 = {_0, _9438} + {_0, _10462};
  wire [3:0] _23997 = {_0, _23995} + {_0, _0, _23996};
  wire _23998 = _12301 < _23997;
  wire _23999 = r748 ^ _23998;
  wire _24000 = _12298 ? coded_block[748] : r748;
  wire _24001 = _12296 ? _23999 : _24000;
  always @ (posedge reset or posedge clock) if (reset) r748 <= 1'd0; else if (_12300) r748 <= _24001;
  wire [1:0] _24002 = {_0, _576} + {_0, _3580};
  wire [1:0] _24003 = {_0, _5215} + {_0, _6973};
  wire [2:0] _24004 = {_0, _24002} + {_0, _24003};
  wire [1:0] _24005 = {_0, _9980} + {_0, _11516};
  wire [3:0] _24006 = {_0, _24004} + {_0, _0, _24005};
  wire _24007 = _12301 < _24006;
  wire _24008 = r747 ^ _24007;
  wire _24009 = _12298 ? coded_block[747] : r747;
  wire _24010 = _12296 ? _24008 : _24009;
  always @ (posedge reset or posedge clock) if (reset) r747 <= 1'd0; else if (_12300) r747 <= _24010;
  wire [1:0] _24011 = {_0, _608} + {_0, _2941};
  wire [1:0] _24012 = {_0, _5663} + {_0, _7293};
  wire [2:0] _24013 = {_0, _24011} + {_0, _24012};
  wire [1:0] _24014 = {_0, _9054} + {_0, _12061};
  wire [3:0] _24015 = {_0, _24013} + {_0, _0, _24014};
  wire _24016 = _12301 < _24015;
  wire _24017 = r746 ^ _24016;
  wire _24018 = _12298 ? coded_block[746] : r746;
  wire _24019 = _12296 ? _24017 : _24018;
  always @ (posedge reset or posedge clock) if (reset) r746 <= 1'd0; else if (_12300) r746 <= _24019;
  wire [1:0] _24020 = {_0, _639} + {_0, _3870};
  wire [1:0] _24021 = {_0, _5022} + {_0, _7741};
  wire [2:0] _24022 = {_0, _24020} + {_0, _24021};
  wire [1:0] _24023 = {_0, _9375} + {_0, _11132};
  wire [3:0] _24024 = {_0, _24022} + {_0, _0, _24023};
  wire _24025 = _12301 < _24024;
  wire _24026 = r745 ^ _24025;
  wire _24027 = _12298 ? coded_block[745] : r745;
  wire _24028 = _12296 ? _24026 : _24027;
  always @ (posedge reset or posedge clock) if (reset) r745 <= 1'd0; else if (_12300) r745 <= _24028;
  wire [1:0] _24029 = {_0, _703} + {_0, _3422};
  wire [1:0] _24030 = {_0, _6045} + {_0, _8028};
  wire [2:0] _24031 = {_0, _24029} + {_0, _24030};
  wire [1:0] _24032 = {_0, _9181} + {_0, _11900};
  wire [3:0] _24033 = {_0, _24031} + {_0, _0, _24032};
  wire _24034 = _12301 < _24033;
  wire _24035 = r744 ^ _24034;
  wire _24036 = _12298 ? coded_block[744] : r744;
  wire _24037 = _12296 ? _24035 : _24036;
  always @ (posedge reset or posedge clock) if (reset) r744 <= 1'd0; else if (_12300) r744 <= _24037;
  wire [1:0] _24038 = {_0, _735} + {_0, _3678};
  wire [1:0] _24039 = {_0, _5501} + {_0, _8123};
  wire [2:0] _24040 = {_0, _24038} + {_0, _24039};
  wire [1:0] _24041 = {_0, _10108} + {_0, _11259};
  wire [3:0] _24042 = {_0, _24040} + {_0, _0, _24041};
  wire _24043 = _12301 < _24042;
  wire _24044 = r743 ^ _24043;
  wire _24045 = _12298 ? coded_block[743] : r743;
  wire _24046 = _12296 ? _24044 : _24045;
  always @ (posedge reset or posedge clock) if (reset) r743 <= 1'd0; else if (_12300) r743 <= _24046;
  wire [1:0] _24047 = {_0, _766} + {_0, _2557};
  wire [1:0] _24048 = {_0, _5757} + {_0, _7581};
  wire [2:0] _24049 = {_0, _24047} + {_0, _24048};
  wire [1:0] _24050 = {_0, _10204} + {_0, _12188};
  wire [3:0] _24051 = {_0, _24049} + {_0, _0, _24050};
  wire _24052 = _12301 < _24051;
  wire _24053 = r742 ^ _24052;
  wire _24054 = _12298 ? coded_block[742] : r742;
  wire _24055 = _12296 ? _24053 : _24054;
  always @ (posedge reset or posedge clock) if (reset) r742 <= 1'd0; else if (_12300) r742 <= _24055;
  wire [1:0] _24056 = {_0, _800} + {_0, _2208};
  wire [1:0] _24057 = {_0, _4640} + {_0, _7837};
  wire [2:0] _24058 = {_0, _24056} + {_0, _24057};
  wire [1:0] _24059 = {_0, _9661} + {_0, _12282};
  wire [3:0] _24060 = {_0, _24058} + {_0, _0, _24059};
  wire _24061 = _12301 < _24060;
  wire _24062 = r741 ^ _24061;
  wire _24063 = _12298 ? coded_block[741] : r741;
  wire _24064 = _12296 ? _24062 : _24063;
  always @ (posedge reset or posedge clock) if (reset) r741 <= 1'd0; else if (_12300) r741 <= _24064;
  wire [1:0] _24065 = {_0, _831} + {_0, _2430};
  wire [1:0] _24066 = {_0, _4287} + {_0, _6718};
  wire [2:0] _24067 = {_0, _24065} + {_0, _24066};
  wire [1:0] _24068 = {_0, _9917} + {_0, _11740};
  wire [3:0] _24069 = {_0, _24067} + {_0, _0, _24068};
  wire _24070 = _12301 < _24069;
  wire _24071 = r740 ^ _24070;
  wire _24072 = _12298 ? coded_block[740] : r740;
  wire _24073 = _12296 ? _24071 : _24072;
  always @ (posedge reset or posedge clock) if (reset) r740 <= 1'd0; else if (_12300) r740 <= _24073;
  wire [1:0] _24074 = {_0, _863} + {_0, _2302};
  wire [1:0] _24075 = {_0, _4511} + {_0, _6366};
  wire [2:0] _24076 = {_0, _24074} + {_0, _24075};
  wire [1:0] _24077 = {_0, _8799} + {_0, _11996};
  wire [3:0] _24078 = {_0, _24076} + {_0, _0, _24077};
  wire _24079 = _12301 < _24078;
  wire _24080 = r739 ^ _24079;
  wire _24081 = _12298 ? coded_block[739] : r739;
  wire _24082 = _12296 ? _24080 : _24081;
  always @ (posedge reset or posedge clock) if (reset) r739 <= 1'd0; else if (_12300) r739 <= _24082;
  wire [1:0] _24083 = {_0, _894} + {_0, _2655};
  wire [1:0] _24084 = {_0, _4384} + {_0, _6589};
  wire [2:0] _24085 = {_0, _24083} + {_0, _24084};
  wire [1:0] _24086 = {_0, _8446} + {_0, _10877};
  wire [3:0] _24087 = {_0, _24085} + {_0, _0, _24086};
  wire _24088 = _12301 < _24087;
  wire _24089 = r738 ^ _24088;
  wire _24090 = _12298 ? coded_block[738] : r738;
  wire _24091 = _12296 ? _24089 : _24090;
  always @ (posedge reset or posedge clock) if (reset) r738 <= 1'd0; else if (_12300) r738 <= _24091;
  wire [1:0] _24092 = {_0, _927} + {_0, _3390};
  wire [1:0] _24093 = {_0, _4734} + {_0, _6462};
  wire [2:0] _24094 = {_0, _24092} + {_0, _24093};
  wire [1:0] _24095 = {_0, _8670} + {_0, _10527};
  wire [3:0] _24096 = {_0, _24094} + {_0, _0, _24095};
  wire _24097 = _12301 < _24096;
  wire _24098 = r737 ^ _24097;
  wire _24099 = _12298 ? coded_block[737] : r737;
  wire _24100 = _12296 ? _24098 : _24099;
  always @ (posedge reset or posedge clock) if (reset) r737 <= 1'd0; else if (_12300) r737 <= _24100;
  wire [1:0] _24101 = {_0, _990} + {_0, _3549};
  wire [1:0] _24102 = {_0, _6076} + {_0, _7548};
  wire [2:0] _24103 = {_0, _24101} + {_0, _24102};
  wire [1:0] _24104 = {_0, _8894} + {_0, _10621};
  wire [3:0] _24105 = {_0, _24103} + {_0, _0, _24104};
  wire _24106 = _12301 < _24105;
  wire _24107 = r736 ^ _24106;
  wire _24108 = _12298 ? coded_block[736] : r736;
  wire _24109 = _12296 ? _24107 : _24108;
  always @ (posedge reset or posedge clock) if (reset) r736 <= 1'd0; else if (_12300) r736 <= _24109;
  wire [1:0] _24110 = {_0, _1021} + {_0, _3167};
  wire [1:0] _24111 = {_0, _5628} + {_0, _8155};
  wire [2:0] _24112 = {_0, _24110} + {_0, _24111};
  wire [1:0] _24113 = {_0, _9630} + {_0, _10973};
  wire [3:0] _24114 = {_0, _24112} + {_0, _0, _24113};
  wire _24115 = _12301 < _24114;
  wire _24116 = r735 ^ _24115;
  wire _24117 = _12298 ? coded_block[735] : r735;
  wire _24118 = _12296 ? _24116 : _24117;
  always @ (posedge reset or posedge clock) if (reset) r735 <= 1'd0; else if (_12300) r735 <= _24118;
  wire [1:0] _24119 = {_0, _1057} + {_0, _2175};
  wire [1:0] _24120 = {_0, _5246} + {_0, _7710};
  wire [2:0] _24121 = {_0, _24119} + {_0, _24120};
  wire [1:0] _24122 = {_0, _10235} + {_0, _11708};
  wire [3:0] _24123 = {_0, _24121} + {_0, _0, _24122};
  wire _24124 = _12301 < _24123;
  wire _24125 = r734 ^ _24124;
  wire _24126 = _12298 ? coded_block[734] : r734;
  wire _24127 = _12296 ? _24125 : _24126;
  always @ (posedge reset or posedge clock) if (reset) r734 <= 1'd0; else if (_12300) r734 <= _24127;
  wire [1:0] _24128 = {_0, _1088} + {_0, _2592};
  wire [1:0] _24129 = {_0, _4256} + {_0, _7326};
  wire [2:0] _24130 = {_0, _24128} + {_0, _24129};
  wire [1:0] _24131 = {_0, _9790} + {_0, _10303};
  wire [3:0] _24132 = {_0, _24130} + {_0, _0, _24131};
  wire _24133 = _12301 < _24132;
  wire _24134 = r733 ^ _24133;
  wire _24135 = _12298 ? coded_block[733] : r733;
  wire _24136 = _12296 ? _24134 : _24135;
  always @ (posedge reset or posedge clock) if (reset) r733 <= 1'd0; else if (_12300) r733 <= _24136;
  wire [1:0] _24137 = {_0, _1120} + {_0, _3068};
  wire [1:0] _24138 = {_0, _4671} + {_0, _6334};
  wire [2:0] _24139 = {_0, _24137} + {_0, _24138};
  wire [1:0] _24140 = {_0, _9406} + {_0, _11869};
  wire [3:0] _24141 = {_0, _24139} + {_0, _0, _24140};
  wire _24142 = _12301 < _24141;
  wire _24143 = r732 ^ _24142;
  wire _24144 = _12298 ? coded_block[732] : r732;
  wire _24145 = _12296 ? _24143 : _24144;
  always @ (posedge reset or posedge clock) if (reset) r732 <= 1'd0; else if (_12300) r732 <= _24145;
  wire [1:0] _24146 = {_0, _1151} + {_0, _2494};
  wire [1:0] _24147 = {_0, _5152} + {_0, _6750};
  wire [2:0] _24148 = {_0, _24146} + {_0, _24147};
  wire [1:0] _24149 = {_0, _8415} + {_0, _11485};
  wire [3:0] _24150 = {_0, _24148} + {_0, _0, _24149};
  wire _24151 = _12301 < _24150;
  wire _24152 = r731 ^ _24151;
  wire _24153 = _12298 ? coded_block[731] : r731;
  wire _24154 = _12296 ? _24152 : _24153;
  always @ (posedge reset or posedge clock) if (reset) r731 <= 1'd0; else if (_12300) r731 <= _24154;
  wire [1:0] _24155 = {_0, _1215} + {_0, _3486};
  wire [1:0] _24156 = {_0, _5884} + {_0, _6652};
  wire [2:0] _24157 = {_0, _24155} + {_0, _24156};
  wire [1:0] _24158 = {_0, _9311} + {_0, _10910};
  wire [3:0] _24159 = {_0, _24157} + {_0, _0, _24158};
  wire _24160 = _12301 < _24159;
  wire _24161 = r730 ^ _24160;
  wire _24162 = _12298 ? coded_block[730] : r730;
  wire _24163 = _12296 ? _24161 : _24162;
  always @ (posedge reset or posedge clock) if (reset) r730 <= 1'd0; else if (_12300) r730 <= _24163;
  wire [1:0] _24164 = {_0, _1247} + {_0, _3646};
  wire [1:0] _24165 = {_0, _5565} + {_0, _7965};
  wire [2:0] _24166 = {_0, _24164} + {_0, _24165};
  wire [1:0] _24167 = {_0, _8736} + {_0, _11389};
  wire [3:0] _24168 = {_0, _24166} + {_0, _0, _24167};
  wire _24169 = _12301 < _24168;
  wire _24170 = r729 ^ _24169;
  wire _24171 = _12298 ? coded_block[729] : r729;
  wire _24172 = _12296 ? _24170 : _24171;
  always @ (posedge reset or posedge clock) if (reset) r729 <= 1'd0; else if (_12300) r729 <= _24172;
  wire [1:0] _24173 = {_0, _1278} + {_0, _3453};
  wire [1:0] _24174 = {_0, _5726} + {_0, _7644};
  wire [2:0] _24175 = {_0, _24173} + {_0, _24174};
  wire [1:0] _24176 = {_0, _10045} + {_0, _10814};
  wire [3:0] _24177 = {_0, _24175} + {_0, _0, _24176};
  wire _24178 = _12301 < _24177;
  wire _24179 = r728 ^ _24178;
  wire _24180 = _12298 ? coded_block[728] : r728;
  wire _24181 = _12296 ? _24179 : _24180;
  always @ (posedge reset or posedge clock) if (reset) r728 <= 1'd0; else if (_12300) r728 <= _24181;
  wire [1:0] _24182 = {_0, _1312} + {_0, _3836};
  wire [1:0] _24183 = {_0, _5534} + {_0, _7804};
  wire [2:0] _24184 = {_0, _24182} + {_0, _24183};
  wire [1:0] _24185 = {_0, _9724} + {_0, _12124};
  wire [3:0] _24186 = {_0, _24184} + {_0, _0, _24185};
  wire _24187 = _12301 < _24186;
  wire _24188 = r727 ^ _24187;
  wire _24189 = _12298 ? coded_block[727] : r727;
  wire _24190 = _12296 ? _24188 : _24189;
  always @ (posedge reset or posedge clock) if (reset) r727 <= 1'd0; else if (_12300) r727 <= _24190;
  wire [1:0] _24191 = {_0, _1343} + {_0, _2974};
  wire [1:0] _24192 = {_0, _5918} + {_0, _7612};
  wire [2:0] _24193 = {_0, _24191} + {_0, _24192};
  wire [1:0] _24194 = {_0, _9886} + {_0, _11806};
  wire [3:0] _24195 = {_0, _24193} + {_0, _0, _24194};
  wire _24196 = _12301 < _24195;
  wire _24197 = r726 ^ _24196;
  wire _24198 = _12298 ? coded_block[726] : r726;
  wire _24199 = _12296 ? _24197 : _24198;
  always @ (posedge reset or posedge clock) if (reset) r726 <= 1'd0; else if (_12300) r726 <= _24199;
  wire [1:0] _24200 = {_0, _1375} + {_0, _2750};
  wire [1:0] _24201 = {_0, _5053} + {_0, _7996};
  wire [2:0] _24202 = {_0, _24200} + {_0, _24201};
  wire [1:0] _24203 = {_0, _9693} + {_0, _11964};
  wire [3:0] _24204 = {_0, _24202} + {_0, _0, _24203};
  wire _24205 = _12301 < _24204;
  wire _24206 = r725 ^ _24205;
  wire _24207 = _12298 ? coded_block[725] : r725;
  wire _24208 = _12296 ? _24206 : _24207;
  always @ (posedge reset or posedge clock) if (reset) r725 <= 1'd0; else if (_12300) r725 <= _24208;
  wire [1:0] _24209 = {_0, _1439} + {_0, _3262};
  wire [1:0] _24210 = {_0, _5407} + {_0, _6908};
  wire [2:0] _24211 = {_0, _24209} + {_0, _24210};
  wire [1:0] _24212 = {_0, _9212} + {_0, _12155};
  wire [3:0] _24213 = {_0, _24211} + {_0, _0, _24212};
  wire _24214 = _12301 < _24213;
  wire _24215 = r724 ^ _24214;
  wire _24216 = _12298 ? coded_block[724] : r724;
  wire _24217 = _12296 ? _24215 : _24216;
  always @ (posedge reset or posedge clock) if (reset) r724 <= 1'd0; else if (_12300) r724 <= _24217;
  wire [1:0] _24218 = {_0, _1470} + {_0, _2367};
  wire [1:0] _24219 = {_0, _5342} + {_0, _7485};
  wire [2:0] _24220 = {_0, _24218} + {_0, _24219};
  wire [1:0] _24221 = {_0, _8991} + {_0, _11295};
  wire [3:0] _24222 = {_0, _24220} + {_0, _0, _24221};
  wire _24223 = _12301 < _24222;
  wire _24224 = r723 ^ _24223;
  wire _24225 = _12298 ? coded_block[723] : r723;
  wire _24226 = _12296 ? _24224 : _24225;
  always @ (posedge reset or posedge clock) if (reset) r723 <= 1'd0; else if (_12300) r723 <= _24226;
  wire [1:0] _24227 = {_0, _255} + {_0, _2494};
  wire [1:0] _24228 = {_0, _4734} + {_0, _7420};
  wire [2:0] _24229 = {_0, _24227} + {_0, _24228};
  wire [1:0] _24230 = {_0, _9212} + {_0, _10462};
  wire [3:0] _24231 = {_0, _24229} + {_0, _0, _24230};
  wire _24232 = _12301 < _24231;
  wire _24233 = r722 ^ _24232;
  wire _24234 = _12298 ? coded_block[722] : r722;
  wire _24235 = _12296 ? _24233 : _24234;
  always @ (posedge reset or posedge clock) if (reset) r722 <= 1'd0; else if (_12300) r722 <= _24235;
  wire [1:0] _24236 = {_0, _863} + {_0, _2557};
  wire [1:0] _24237 = {_0, _5694} + {_0, _8059};
  wire [2:0] _24238 = {_0, _24236} + {_0, _24237};
  wire [1:0] _24239 = {_0, _8543} + {_0, _11964};
  wire [3:0] _24240 = {_0, _24238} + {_0, _0, _24239};
  wire _24241 = _12301 < _24240;
  wire _24242 = r721 ^ _24241;
  wire _24243 = _12298 ? coded_block[721] : r721;
  wire _24244 = _12296 ? _24242 : _24243;
  always @ (posedge reset or posedge clock) if (reset) r721 <= 1'd0; else if (_12300) r721 <= _24244;
  wire [1:0] _24245 = {_0, _894} + {_0, _4060};
  wire [1:0] _24246 = {_0, _4640} + {_0, _7773};
  wire [2:0] _24247 = {_0, _24245} + {_0, _24246};
  wire [1:0] _24248 = {_0, _10141} + {_0, _10621};
  wire [3:0] _24249 = {_0, _24247} + {_0, _0, _24248};
  wire _24250 = _12301 < _24249;
  wire _24251 = r720 ^ _24250;
  wire _24252 = _12298 ? coded_block[720] : r720;
  wire _24253 = _12296 ? _24251 : _24252;
  always @ (posedge reset or posedge clock) if (reset) r720 <= 1'd0; else if (_12300) r720 <= _24253;
  wire [1:0] _24254 = {_0, _927} + {_0, _3037};
  wire [1:0] _24255 = {_0, _6139} + {_0, _6718};
  wire [2:0] _24256 = {_0, _24254} + {_0, _24255};
  wire [1:0] _24257 = {_0, _9853} + {_0, _12219};
  wire [3:0] _24258 = {_0, _24256} + {_0, _0, _24257};
  wire _24259 = _12301 < _24258;
  wire _24260 = r719 ^ _24259;
  wire _24261 = _12298 ? coded_block[719] : r719;
  wire _24262 = _12296 ? _24260 : _24261;
  always @ (posedge reset or posedge clock) if (reset) r719 <= 1'd0; else if (_12300) r719 <= _24262;
  wire [1:0] _24263 = {_0, _990} + {_0, _2974};
  wire [1:0] _24264 = {_0, _5884} + {_0, _7199};
  wire [2:0] _24265 = {_0, _24263} + {_0, _24264};
  wire [1:0] _24266 = {_0, _8288} + {_0, _10877};
  wire [3:0] _24267 = {_0, _24265} + {_0, _0, _24266};
  wire _24268 = _12301 < _24267;
  wire _24269 = r718 ^ _24268;
  wire _24270 = _12298 ? coded_block[718] : r718;
  wire _24271 = _12296 ? _24269 : _24270;
  always @ (posedge reset or posedge clock) if (reset) r718 <= 1'd0; else if (_12300) r718 <= _24271;
  wire [1:0] _24272 = {_0, _1021} + {_0, _2494};
  wire [1:0] _24273 = {_0, _5053} + {_0, _7965};
  wire [2:0] _24274 = {_0, _24272} + {_0, _24273};
  wire [1:0] _24275 = {_0, _9279} + {_0, _10366};
  wire [3:0] _24276 = {_0, _24274} + {_0, _0, _24275};
  wire _24277 = _12301 < _24276;
  wire _24278 = r717 ^ _24277;
  wire _24279 = _12298 ? coded_block[717] : r717;
  wire _24280 = _12296 ? _24278 : _24279;
  always @ (posedge reset or posedge clock) if (reset) r717 <= 1'd0; else if (_12300) r717 <= _24280;
  wire [1:0] _24281 = {_0, _1088} + {_0, _3964};
  wire [1:0] _24282 = {_0, _4703} + {_0, _6652};
  wire [2:0] _24283 = {_0, _24281} + {_0, _24282};
  wire [1:0] _24284 = {_0, _9212} + {_0, _12124};
  wire [3:0] _24285 = {_0, _24283} + {_0, _0, _24284};
  wire _24286 = _12301 < _24285;
  wire _24287 = r716 ^ _24286;
  wire _24288 = _12298 ? coded_block[716] : r716;
  wire _24289 = _12296 ? _24287 : _24288;
  always @ (posedge reset or posedge clock) if (reset) r716 <= 1'd0; else if (_12300) r716 <= _24289;
  wire [1:0] _24290 = {_0, _1120} + {_0, _3198};
  wire [1:0] _24291 = {_0, _6045} + {_0, _6781};
  wire [2:0] _24292 = {_0, _24290} + {_0, _24291};
  wire [1:0] _24293 = {_0, _8736} + {_0, _11295};
  wire [3:0] _24294 = {_0, _24292} + {_0, _0, _24293};
  wire _24295 = _12301 < _24294;
  wire _24296 = r715 ^ _24295;
  wire _24297 = _12298 ? coded_block[715] : r715;
  wire _24298 = _12296 ? _24296 : _24297;
  always @ (posedge reset or posedge clock) if (reset) r715 <= 1'd0; else if (_12300) r715 <= _24298;
  wire [1:0] _24299 = {_0, _1151} + {_0, _3167};
  wire [1:0] _24300 = {_0, _5279} + {_0, _8123};
  wire [2:0] _24301 = {_0, _24299} + {_0, _24300};
  wire [1:0] _24302 = {_0, _8863} + {_0, _10814};
  wire [3:0] _24303 = {_0, _24301} + {_0, _0, _24302};
  wire _24304 = _12301 < _24303;
  wire _24305 = r714 ^ _24304;
  wire _24306 = _12298 ? coded_block[714] : r714;
  wire _24307 = _12296 ? _24305 : _24306;
  always @ (posedge reset or posedge clock) if (reset) r714 <= 1'd0; else if (_12300) r714 <= _24307;
  wire [1:0] _24308 = {_0, _1215} + {_0, _2271};
  wire [1:0] _24309 = {_0, _6076} + {_0, _7326};
  wire [2:0] _24310 = {_0, _24308} + {_0, _24309};
  wire [1:0] _24311 = {_0, _9438} + {_0, _12282};
  wire [3:0] _24312 = {_0, _24310} + {_0, _0, _24311};
  wire _24313 = _12301 < _24312;
  wire _24314 = r713 ^ _24313;
  wire _24315 = _12298 ? coded_block[713] : r713;
  wire _24316 = _12296 ? _24314 : _24315;
  always @ (posedge reset or posedge clock) if (reset) r713 <= 1'd0; else if (_12300) r713 <= _24316;
  wire [1:0] _24317 = {_0, _1247} + {_0, _3678};
  wire [1:0] _24318 = {_0, _4350} + {_0, _8155};
  wire [2:0] _24319 = {_0, _24317} + {_0, _24318};
  wire [1:0] _24320 = {_0, _9406} + {_0, _11516};
  wire [3:0] _24321 = {_0, _24319} + {_0, _0, _24320};
  wire _24322 = _12301 < _24321;
  wire _24323 = r712 ^ _24322;
  wire _24324 = _12298 ? coded_block[712] : r712;
  wire _24325 = _12296 ? _24323 : _24324;
  always @ (posedge reset or posedge clock) if (reset) r712 <= 1'd0; else if (_12300) r712 <= _24325;
  wire [1:0] _24326 = {_0, _1278} + {_0, _3517};
  wire [1:0] _24327 = {_0, _5757} + {_0, _6431};
  wire [2:0] _24328 = {_0, _24326} + {_0, _24327};
  wire [1:0] _24329 = {_0, _10235} + {_0, _11485};
  wire [3:0] _24330 = {_0, _24328} + {_0, _0, _24329};
  wire _24331 = _12301 < _24330;
  wire _24332 = r711 ^ _24331;
  wire _24333 = _12298 ? coded_block[711] : r711;
  wire _24334 = _12296 ? _24332 : _24333;
  always @ (posedge reset or posedge clock) if (reset) r711 <= 1'd0; else if (_12300) r711 <= _24334;
  wire [1:0] _24335 = {_0, _1343} + {_0, _3549};
  wire [1:0] _24336 = {_0, _4129} + {_0, _7675};
  wire [2:0] _24337 = {_0, _24335} + {_0, _24336};
  wire [1:0] _24338 = {_0, _9917} + {_0, _10590};
  wire [3:0] _24339 = {_0, _24337} + {_0, _0, _24338};
  wire _24340 = _12301 < _24339;
  wire _24341 = r710 ^ _24340;
  wire _24342 = _12298 ? coded_block[710] : r710;
  wire _24343 = _12296 ? _24341 : _24342;
  always @ (posedge reset or posedge clock) if (reset) r710 <= 1'd0; else if (_12300) r710 <= _24343;
  wire [1:0] _24344 = {_0, _1375} + {_0, _3742};
  wire [1:0] _24345 = {_0, _5628} + {_0, _6176};
  wire [2:0] _24346 = {_0, _24344} + {_0, _24345};
  wire [1:0] _24347 = {_0, _9759} + {_0, _11996};
  wire [3:0] _24348 = {_0, _24346} + {_0, _0, _24347};
  wire _24349 = _12301 < _24348;
  wire _24350 = r709 ^ _24349;
  wire _24351 = _12298 ? coded_block[709] : r709;
  wire _24352 = _12296 ? _24350 : _24351;
  always @ (posedge reset or posedge clock) if (reset) r709 <= 1'd0; else if (_12300) r709 <= _24352;
  wire [1:0] _24353 = {_0, _1406} + {_0, _2367};
  wire [1:0] _24354 = {_0, _5821} + {_0, _7710};
  wire [2:0] _24355 = {_0, _24353} + {_0, _24354};
  wire [1:0] _24356 = {_0, _8225} + {_0, _11837};
  wire [3:0] _24357 = {_0, _24355} + {_0, _0, _24356};
  wire _24358 = _12301 < _24357;
  wire _24359 = r708 ^ _24358;
  wire _24360 = _12298 ? coded_block[708] : r708;
  wire _24361 = _12296 ? _24359 : _24360;
  always @ (posedge reset or posedge clock) if (reset) r708 <= 1'd0; else if (_12300) r708 <= _24361;
  wire [1:0] _24362 = {_0, _1439} + {_0, _2112};
  wire [1:0] _24363 = {_0, _4447} + {_0, _7900};
  wire [2:0] _24364 = {_0, _24362} + {_0, _24363};
  wire [1:0] _24365 = {_0, _9790} + {_0, _10272};
  wire [3:0] _24366 = {_0, _24364} + {_0, _0, _24365};
  wire _24367 = _12301 < _24366;
  wire _24368 = r707 ^ _24367;
  wire _24369 = _12298 ? coded_block[707] : r707;
  wire _24370 = _12296 ? _24368 : _24369;
  always @ (posedge reset or posedge clock) if (reset) r707 <= 1'd0; else if (_12300) r707 <= _24370;
  wire [1:0] _24371 = {_0, _1470} + {_0, _3325};
  wire [1:0] _24372 = {_0, _4192} + {_0, _6525};
  wire [2:0] _24373 = {_0, _24371} + {_0, _24372};
  wire [1:0] _24374 = {_0, _9980} + {_0, _11869};
  wire [3:0] _24375 = {_0, _24373} + {_0, _0, _24374};
  wire _24376 = _12301 < _24375;
  wire _24377 = r706 ^ _24376;
  wire _24378 = _12298 ? coded_block[706] : r706;
  wire _24379 = _12296 ? _24377 : _24378;
  always @ (posedge reset or posedge clock) if (reset) r706 <= 1'd0; else if (_12300) r706 <= _24379;
  wire [1:0] _24380 = {_0, _1502} + {_0, _3390};
  wire [1:0] _24381 = {_0, _5407} + {_0, _6270};
  wire [2:0] _24382 = {_0, _24380} + {_0, _24381};
  wire [1:0] _24383 = {_0, _8607} + {_0, _12061};
  wire [3:0] _24384 = {_0, _24382} + {_0, _0, _24383};
  wire _24385 = _12301 < _24384;
  wire _24386 = r705 ^ _24385;
  wire _24387 = _12298 ? coded_block[705] : r705;
  wire _24388 = _12296 ? _24386 : _24387;
  always @ (posedge reset or posedge clock) if (reset) r705 <= 1'd0; else if (_12300) r705 <= _24388;
  wire [1:0] _24389 = {_0, _1568} + {_0, _2878};
  wire [1:0] _24390 = {_0, _4256} + {_0, _7548};
  wire [2:0] _24391 = {_0, _24389} + {_0, _24390};
  wire [1:0] _24392 = {_0, _9566} + {_0, _10430};
  wire [3:0] _24393 = {_0, _24391} + {_0, _0, _24392};
  wire _24394 = _12301 < _24393;
  wire _24395 = r704 ^ _24394;
  wire _24396 = _12298 ? coded_block[704] : r704;
  wire _24397 = _12296 ? _24395 : _24396;
  always @ (posedge reset or posedge clock) if (reset) r704 <= 1'd0; else if (_12300) r704 <= _24397;
  wire [1:0] _24398 = {_0, _1599} + {_0, _2782};
  wire [1:0] _24399 = {_0, _4958} + {_0, _6334};
  wire [2:0] _24400 = {_0, _24398} + {_0, _24399};
  wire [1:0] _24401 = {_0, _9630} + {_0, _11644};
  wire [3:0] _24402 = {_0, _24400} + {_0, _0, _24401};
  wire _24403 = _12301 < _24402;
  wire _24404 = r703 ^ _24403;
  wire _24405 = _12298 ? coded_block[703] : r703;
  wire _24406 = _12296 ? _24404 : _24405;
  always @ (posedge reset or posedge clock) if (reset) r703 <= 1'd0; else if (_12300) r703 <= _24406;
  wire [1:0] _24407 = {_0, _1631} + {_0, _3294};
  wire [1:0] _24408 = {_0, _4861} + {_0, _7036};
  wire [2:0] _24409 = {_0, _24407} + {_0, _24408};
  wire [1:0] _24410 = {_0, _8415} + {_0, _11708};
  wire [3:0] _24411 = {_0, _24409} + {_0, _0, _24410};
  wire _24412 = _12301 < _24411;
  wire _24413 = r702 ^ _24412;
  wire _24414 = _12298 ? coded_block[702] : r702;
  wire _24415 = _12296 ? _24413 : _24414;
  always @ (posedge reset or posedge clock) if (reset) r702 <= 1'd0; else if (_12300) r702 <= _24415;
  wire [1:0] _24416 = {_0, _1662} + {_0, _2144};
  wire [1:0] _24417 = {_0, _5373} + {_0, _6942};
  wire [2:0] _24418 = {_0, _24416} + {_0, _24417};
  wire [1:0] _24419 = {_0, _9118} + {_0, _10493};
  wire [3:0] _24420 = {_0, _24418} + {_0, _0, _24419};
  wire _24421 = _12301 < _24420;
  wire _24422 = r701 ^ _24421;
  wire _24423 = _12298 ? coded_block[701] : r701;
  wire _24424 = _12296 ? _24422 : _24423;
  always @ (posedge reset or posedge clock) if (reset) r701 <= 1'd0; else if (_12300) r701 <= _24424;
  wire [1:0] _24425 = {_0, _1695} + {_0, _3422};
  wire [1:0] _24426 = {_0, _4223} + {_0, _7454};
  wire [2:0] _24427 = {_0, _24425} + {_0, _24426};
  wire [1:0] _24428 = {_0, _9022} + {_0, _11196};
  wire [3:0] _24429 = {_0, _24427} + {_0, _0, _24428};
  wire _24430 = _12301 < _24429;
  wire _24431 = r700 ^ _24430;
  wire _24432 = _12298 ? coded_block[700] : r700;
  wire _24433 = _12296 ? _24431 : _24432;
  always @ (posedge reset or posedge clock) if (reset) r700 <= 1'd0; else if (_12300) r700 <= _24433;
  wire [1:0] _24434 = {_0, _1726} + {_0, _2463};
  wire [1:0] _24435 = {_0, _5501} + {_0, _6303};
  wire [2:0] _24436 = {_0, _24434} + {_0, _24435};
  wire [1:0] _24437 = {_0, _9534} + {_0, _11101};
  wire [3:0] _24438 = {_0, _24436} + {_0, _0, _24437};
  wire _24439 = _12301 < _24438;
  wire _24440 = r699 ^ _24439;
  wire _24441 = _12298 ? coded_block[699] : r699;
  wire _24442 = _12296 ? _24440 : _24441;
  always @ (posedge reset or posedge clock) if (reset) r699 <= 1'd0; else if (_12300) r699 <= _24442;
  wire [1:0] _24443 = {_0, _1758} + {_0, _3005};
  wire [1:0] _24444 = {_0, _4542} + {_0, _7581};
  wire [2:0] _24445 = {_0, _24443} + {_0, _24444};
  wire [1:0] _24446 = {_0, _8383} + {_0, _11613};
  wire [3:0] _24447 = {_0, _24445} + {_0, _0, _24446};
  wire _24448 = _12301 < _24447;
  wire _24449 = r698 ^ _24448;
  wire _24450 = _12298 ? coded_block[698] : r698;
  wire _24451 = _12296 ? _24449 : _24450;
  always @ (posedge reset or posedge clock) if (reset) r698 <= 1'd0; else if (_12300) r698 <= _24451;
  wire [1:0] _24452 = {_0, _1789} + {_0, _4091};
  wire [1:0] _24453 = {_0, _5085} + {_0, _6621};
  wire [2:0] _24454 = {_0, _24452} + {_0, _24453};
  wire [1:0] _24455 = {_0, _9661} + {_0, _10462};
  wire [3:0] _24456 = {_0, _24454} + {_0, _0, _24455};
  wire _24457 = _12301 < _24456;
  wire _24458 = r697 ^ _24457;
  wire _24459 = _12298 ? coded_block[697] : r697;
  wire _24460 = _12296 ? _24458 : _24459;
  always @ (posedge reset or posedge clock) if (reset) r697 <= 1'd0; else if (_12300) r697 <= _24460;
  wire [1:0] _24461 = {_0, _1823} + {_0, _2399};
  wire [1:0] _24462 = {_0, _4160} + {_0, _7163};
  wire [2:0] _24463 = {_0, _24461} + {_0, _24462};
  wire [1:0] _24464 = {_0, _8701} + {_0, _11740};
  wire [3:0] _24465 = {_0, _24463} + {_0, _0, _24464};
  wire _24466 = _12301 < _24465;
  wire _24467 = r696 ^ _24466;
  wire _24468 = _12298 ? coded_block[696] : r696;
  wire _24469 = _12296 ? _24467 : _24468;
  always @ (posedge reset or posedge clock) if (reset) r696 <= 1'd0; else if (_12300) r696 <= _24469;
  wire [1:0] _24470 = {_0, _1854} + {_0, _2847};
  wire [1:0] _24471 = {_0, _4478} + {_0, _6239};
  wire [2:0] _24472 = {_0, _24470} + {_0, _24471};
  wire [1:0] _24473 = {_0, _9248} + {_0, _10783};
  wire [3:0] _24474 = {_0, _24472} + {_0, _0, _24473};
  wire _24475 = _12301 < _24474;
  wire _24476 = r695 ^ _24475;
  wire _24477 = _12298 ? coded_block[695] : r695;
  wire _24478 = _12296 ? _24476 : _24477;
  always @ (posedge reset or posedge clock) if (reset) r695 <= 1'd0; else if (_12300) r695 <= _24478;
  wire [1:0] _24479 = {_0, _1886} + {_0, _2208};
  wire [1:0] _24480 = {_0, _4926} + {_0, _6558};
  wire [2:0] _24481 = {_0, _24479} + {_0, _24480};
  wire [1:0] _24482 = {_0, _8319} + {_0, _11326};
  wire [3:0] _24483 = {_0, _24481} + {_0, _0, _24482};
  wire _24484 = _12301 < _24483;
  wire _24485 = r694 ^ _24484;
  wire _24486 = _12298 ? coded_block[694] : r694;
  wire _24487 = _12296 ? _24485 : _24486;
  always @ (posedge reset or posedge clock) if (reset) r694 <= 1'd0; else if (_12300) r694 <= _24487;
  wire [1:0] _24488 = {_0, _1917} + {_0, _3135};
  wire [1:0] _24489 = {_0, _4287} + {_0, _7005};
  wire [2:0] _24490 = {_0, _24488} + {_0, _24489};
  wire [1:0] _24491 = {_0, _8638} + {_0, _10399};
  wire [3:0] _24492 = {_0, _24490} + {_0, _0, _24491};
  wire _24493 = _12301 < _24492;
  wire _24494 = r693 ^ _24493;
  wire _24495 = _12298 ? coded_block[693] : r693;
  wire _24496 = _12296 ? _24494 : _24495;
  always @ (posedge reset or posedge clock) if (reset) r693 <= 1'd0; else if (_12300) r693 <= _24496;
  wire [1:0] _24497 = {_0, _1950} + {_0, _3231};
  wire [1:0] _24498 = {_0, _5215} + {_0, _6366};
  wire [2:0] _24499 = {_0, _24497} + {_0, _24498};
  wire [1:0] _24500 = {_0, _9085} + {_0, _10717};
  wire [3:0] _24501 = {_0, _24499} + {_0, _0, _24500};
  wire _24502 = _12301 < _24501;
  wire _24503 = r692 ^ _24502;
  wire _24504 = _12298 ? coded_block[692] : r692;
  wire _24505 = _12296 ? _24503 : _24504;
  always @ (posedge reset or posedge clock) if (reset) r692 <= 1'd0; else if (_12300) r692 <= _24505;
  wire [1:0] _24506 = {_0, _1981} + {_0, _2686};
  wire [1:0] _24507 = {_0, _5310} + {_0, _7293};
  wire [2:0] _24508 = {_0, _24506} + {_0, _24507};
  wire [1:0] _24509 = {_0, _8446} + {_0, _11165};
  wire [3:0] _24510 = {_0, _24508} + {_0, _0, _24509};
  wire _24511 = _12301 < _24510;
  wire _24512 = r691 ^ _24511;
  wire _24513 = _12298 ? coded_block[691] : r691;
  wire _24514 = _12296 ? _24512 : _24513;
  always @ (posedge reset or posedge clock) if (reset) r691 <= 1'd0; else if (_12300) r691 <= _24514;
  wire [1:0] _24515 = {_0, _2013} + {_0, _2941};
  wire [1:0] _24516 = {_0, _4767} + {_0, _7389};
  wire [2:0] _24517 = {_0, _24515} + {_0, _24516};
  wire [1:0] _24518 = {_0, _9375} + {_0, _10527};
  wire [3:0] _24519 = {_0, _24517} + {_0, _0, _24518};
  wire _24520 = _12301 < _24519;
  wire _24521 = r690 ^ _24520;
  wire _24522 = _12298 ? coded_block[690] : r690;
  wire _24523 = _12296 ? _24521 : _24522;
  always @ (posedge reset or posedge clock) if (reset) r690 <= 1'd0; else if (_12300) r690 <= _24523;
  wire [1:0] _24524 = {_0, _65} + {_0, _3486};
  wire [1:0] _24525 = {_0, _5918} + {_0, _7100};
  wire [2:0] _24526 = {_0, _24524} + {_0, _24525};
  wire [1:0] _24527 = {_0, _8926} + {_0, _11550};
  wire [3:0] _24528 = {_0, _24526} + {_0, _0, _24527};
  wire _24529 = _12301 < _24528;
  wire _24530 = r689 ^ _24529;
  wire _24531 = _12298 ? coded_block[689] : r689;
  wire _24532 = _12296 ? _24530 : _24531;
  always @ (posedge reset or posedge clock) if (reset) r689 <= 1'd0; else if (_12300) r689 <= _24532;
  wire [1:0] _24533 = {_0, _97} + {_0, _3709};
  wire [1:0] _24534 = {_0, _5565} + {_0, _7996};
  wire [2:0] _24535 = {_0, _24533} + {_0, _24534};
  wire [1:0] _24536 = {_0, _9181} + {_0, _11004};
  wire [3:0] _24537 = {_0, _24535} + {_0, _0, _24536};
  wire _24538 = _12301 < _24537;
  wire _24539 = r688 ^ _24538;
  wire _24540 = _12298 ? coded_block[688] : r688;
  wire _24541 = _12296 ? _24539 : _24540;
  always @ (posedge reset or posedge clock) if (reset) r688 <= 1'd0; else if (_12300) r688 <= _24541;
  wire [1:0] _24542 = {_0, _128} + {_0, _3580};
  wire [1:0] _24543 = {_0, _5790} + {_0, _7644};
  wire [2:0] _24544 = {_0, _24542} + {_0, _24543};
  wire [1:0] _24545 = {_0, _10077} + {_0, _11259};
  wire [3:0] _24546 = {_0, _24544} + {_0, _0, _24545};
  wire _24547 = _12301 < _24546;
  wire _24548 = r687 ^ _24547;
  wire _24549 = _12298 ? coded_block[687] : r687;
  wire _24550 = _12296 ? _24548 : _24549;
  always @ (posedge reset or posedge clock) if (reset) r687 <= 1'd0; else if (_12300) r687 <= _24550;
  wire [1:0] _24551 = {_0, _161} + {_0, _3933};
  wire [1:0] _24552 = {_0, _5663} + {_0, _7868};
  wire [2:0] _24553 = {_0, _24551} + {_0, _24552};
  wire [1:0] _24554 = {_0, _9724} + {_0, _12155};
  wire [3:0] _24555 = {_0, _24553} + {_0, _0, _24554};
  wire _24556 = _12301 < _24555;
  wire _24557 = r686 ^ _24556;
  wire _24558 = _12298 ? coded_block[686] : r686;
  wire _24559 = _12296 ? _24557 : _24558;
  always @ (posedge reset or posedge clock) if (reset) r686 <= 1'd0; else if (_12300) r686 <= _24559;
  wire [1:0] _24560 = {_0, _192} + {_0, _2655};
  wire [1:0] _24561 = {_0, _6012} + {_0, _7741};
  wire [2:0] _24562 = {_0, _24560} + {_0, _24561};
  wire [1:0] _24563 = {_0, _9949} + {_0, _11806};
  wire [3:0] _24564 = {_0, _24562} + {_0, _0, _24563};
  wire _24565 = _12301 < _24564;
  wire _24566 = r685 ^ _24565;
  wire _24567 = _12298 ? coded_block[685] : r685;
  wire _24568 = _12296 ? _24566 : _24567;
  always @ (posedge reset or posedge clock) if (reset) r685 <= 1'd0; else if (_12300) r685 <= _24568;
  wire [1:0] _24569 = {_0, _224} + {_0, _3262};
  wire [1:0] _24570 = {_0, _4734} + {_0, _8092};
  wire [2:0] _24571 = {_0, _24569} + {_0, _24570};
  wire [1:0] _24572 = {_0, _9822} + {_0, _12027};
  wire [3:0] _24573 = {_0, _24571} + {_0, _0, _24572};
  wire _24574 = _12301 < _24573;
  wire _24575 = r684 ^ _24574;
  wire _24576 = _12298 ? coded_block[684] : r684;
  wire _24577 = _12296 ? _24575 : _24576;
  always @ (posedge reset or posedge clock) if (reset) r684 <= 1'd0; else if (_12300) r684 <= _24577;
  wire [1:0] _24578 = {_0, _255} + {_0, _2813};
  wire [1:0] _24579 = {_0, _5342} + {_0, _6814};
  wire [2:0] _24580 = {_0, _24578} + {_0, _24579};
  wire [1:0] _24581 = {_0, _10172} + {_0, _11900};
  wire [3:0] _24582 = {_0, _24580} + {_0, _0, _24581};
  wire _24583 = _12301 < _24582;
  wire _24584 = r683 ^ _24583;
  wire _24585 = _12298 ? coded_block[683] : r683;
  wire _24586 = _12296 ? _24584 : _24585;
  always @ (posedge reset or posedge clock) if (reset) r683 <= 1'd0; else if (_12300) r683 <= _24586;
  wire [1:0] _24587 = {_0, _289} + {_0, _2430};
  wire [1:0] _24588 = {_0, _4895} + {_0, _7420};
  wire [2:0] _24589 = {_0, _24587} + {_0, _24588};
  wire [1:0] _24590 = {_0, _8894} + {_0, _12251};
  wire [3:0] _24591 = {_0, _24589} + {_0, _0, _24590};
  wire _24592 = _12301 < _24591;
  wire _24593 = r682 ^ _24592;
  wire _24594 = _12298 ? coded_block[682] : r682;
  wire _24595 = _12296 ? _24593 : _24594;
  always @ (posedge reset or posedge clock) if (reset) r682 <= 1'd0; else if (_12300) r682 <= _24595;
  wire [1:0] _24596 = {_0, _320} + {_0, _3453};
  wire [1:0] _24597 = {_0, _4511} + {_0, _6973};
  wire [2:0] _24598 = {_0, _24596} + {_0, _24597};
  wire [1:0] _24599 = {_0, _9503} + {_0, _10973};
  wire [3:0] _24600 = {_0, _24598} + {_0, _0, _24599};
  wire _24601 = _12301 < _24600;
  wire _24602 = r681 ^ _24601;
  wire _24603 = _12298 ? coded_block[681] : r681;
  wire _24604 = _12296 ? _24602 : _24603;
  always @ (posedge reset or posedge clock) if (reset) r681 <= 1'd0; else if (_12300) r681 <= _24604;
  wire [1:0] _24605 = {_0, _383} + {_0, _2336};
  wire [1:0] _24606 = {_0, _5949} + {_0, _7612};
  wire [2:0] _24607 = {_0, _24605} + {_0, _24606};
  wire [1:0] _24608 = {_0, _8670} + {_0, _11132};
  wire [3:0] _24609 = {_0, _24607} + {_0, _0, _24608};
  wire _24610 = _12301 < _24609;
  wire _24611 = r680 ^ _24610;
  wire _24612 = _12298 ? coded_block[680] : r680;
  wire _24613 = _12296 ? _24611 : _24612;
  always @ (posedge reset or posedge clock) if (reset) r680 <= 1'd0; else if (_12300) r680 <= _24613;
  wire [1:0] _24614 = {_0, _416} + {_0, _3773};
  wire [1:0] _24615 = {_0, _4415} + {_0, _8028};
  wire [2:0] _24616 = {_0, _24614} + {_0, _24615};
  wire [1:0] _24617 = {_0, _9693} + {_0, _10748};
  wire [3:0] _24618 = {_0, _24616} + {_0, _0, _24617};
  wire _24619 = _12301 < _24618;
  wire _24620 = r679 ^ _24619;
  wire _24621 = _12298 ? coded_block[679] : r679;
  wire _24622 = _12296 ? _24620 : _24621;
  always @ (posedge reset or posedge clock) if (reset) r679 <= 1'd0; else if (_12300) r679 <= _24622;
  wire [1:0] _24623 = {_0, _447} + {_0, _3068};
  wire [1:0] _24624 = {_0, _5853} + {_0, _6494};
  wire [2:0] _24625 = {_0, _24623} + {_0, _24624};
  wire [1:0] _24626 = {_0, _10108} + {_0, _11771};
  wire [3:0] _24627 = {_0, _24625} + {_0, _0, _24626};
  wire _24628 = _12301 < _24627;
  wire _24629 = r678 ^ _24628;
  wire _24630 = _12298 ? coded_block[678] : r678;
  wire _24631 = _12296 ? _24629 : _24630;
  always @ (posedge reset or posedge clock) if (reset) r678 <= 1'd0; else if (_12300) r678 <= _24631;
  wire [1:0] _24632 = {_0, _479} + {_0, _2750};
  wire [1:0] _24633 = {_0, _5152} + {_0, _7931};
  wire [2:0] _24634 = {_0, _24632} + {_0, _24633};
  wire [1:0] _24635 = {_0, _8574} + {_0, _12188};
  wire [3:0] _24636 = {_0, _24634} + {_0, _0, _24635};
  wire _24637 = _12301 < _24636;
  wire _24638 = r677 ^ _24637;
  wire _24639 = _12298 ? coded_block[677] : r677;
  wire _24640 = _12296 ? _24638 : _24639;
  always @ (posedge reset or posedge clock) if (reset) r677 <= 1'd0; else if (_12300) r677 <= _24640;
  wire [1:0] _24641 = {_0, _545} + {_0, _2719};
  wire [1:0] _24642 = {_0, _4989} + {_0, _6908};
  wire [2:0] _24643 = {_0, _24641} + {_0, _24642};
  wire [1:0] _24644 = {_0, _9311} + {_0, _12092};
  wire [3:0] _24645 = {_0, _24643} + {_0, _0, _24644};
  wire _24646 = _12301 < _24645;
  wire _24647 = r676 ^ _24646;
  wire _24648 = _12298 ? coded_block[676] : r676;
  wire _24649 = _12296 ? _24647 : _24648;
  always @ (posedge reset or posedge clock) if (reset) r676 <= 1'd0; else if (_12300) r676 <= _24649;
  wire [1:0] _24650 = {_0, _576} + {_0, _3104};
  wire [1:0] _24651 = {_0, _4798} + {_0, _7069};
  wire [2:0] _24652 = {_0, _24650} + {_0, _24651};
  wire [1:0] _24653 = {_0, _8991} + {_0, _11389};
  wire [3:0] _24654 = {_0, _24652} + {_0, _0, _24653};
  wire _24655 = _12301 < _24654;
  wire _24656 = r675 ^ _24655;
  wire _24657 = _12298 ? coded_block[675] : r675;
  wire _24658 = _12296 ? _24656 : _24657;
  always @ (posedge reset or posedge clock) if (reset) r675 <= 1'd0; else if (_12300) r675 <= _24658;
  wire [1:0] _24659 = {_0, _608} + {_0, _2239};
  wire [1:0] _24660 = {_0, _5183} + {_0, _6877};
  wire [2:0] _24661 = {_0, _24659} + {_0, _24660};
  wire [1:0] _24662 = {_0, _9149} + {_0, _11069};
  wire [3:0] _24663 = {_0, _24661} + {_0, _0, _24662};
  wire _24664 = _12301 < _24663;
  wire _24665 = r674 ^ _24664;
  wire _24666 = _12298 ? coded_block[674] : r674;
  wire _24667 = _12296 ? _24665 : _24666;
  always @ (posedge reset or posedge clock) if (reset) r674 <= 1'd0; else if (_12300) r674 <= _24667;
  wire [1:0] _24668 = {_0, _672} + {_0, _2592};
  wire [1:0] _24669 = {_0, _6108} + {_0, _6397};
  wire [2:0] _24670 = {_0, _24668} + {_0, _24669};
  wire [1:0] _24671 = {_0, _9342} + {_0, _11038};
  wire [3:0] _24672 = {_0, _24670} + {_0, _0, _24671};
  wire _24673 = _12301 < _24672;
  wire _24674 = r673 ^ _24673;
  wire _24675 = _12298 ? coded_block[673] : r673;
  wire _24676 = _12296 ? _24674 : _24675;
  always @ (posedge reset or posedge clock) if (reset) r673 <= 1'd0; else if (_12300) r673 <= _24676;
  wire [1:0] _24677 = {_0, _703} + {_0, _2526};
  wire [1:0] _24678 = {_0, _4671} + {_0, _8186};
  wire [2:0] _24679 = {_0, _24677} + {_0, _24678};
  wire [1:0] _24680 = {_0, _8480} + {_0, _11422};
  wire [3:0] _24681 = {_0, _24679} + {_0, _0, _24680};
  wire _24682 = _12301 < _24681;
  wire _24683 = r672 ^ _24682;
  wire _24684 = _12298 ? coded_block[672] : r672;
  wire _24685 = _12296 ? _24683 : _24684;
  always @ (posedge reset or posedge clock) if (reset) r672 <= 1'd0; else if (_12300) r672 <= _24685;
  wire [1:0] _24686 = {_0, _735} + {_0, _3646};
  wire [1:0] _24687 = {_0, _4605} + {_0, _6750};
  wire [2:0] _24688 = {_0, _24686} + {_0, _24687};
  wire [1:0] _24689 = {_0, _8256} + {_0, _10558};
  wire [3:0] _24690 = {_0, _24688} + {_0, _0, _24689};
  wire _24691 = _12301 < _24690;
  wire _24692 = r671 ^ _24691;
  wire _24693 = _12298 ? coded_block[671] : r671;
  wire _24694 = _12296 ? _24692 : _24693;
  always @ (posedge reset or posedge clock) if (reset) r671 <= 1'd0; else if (_12300) r671 <= _24694;
  wire [1:0] _24695 = {_0, _800} + {_0, _3901};
  wire [1:0] _24696 = {_0, _4384} + {_0, _7804};
  wire [2:0] _24697 = {_0, _24695} + {_0, _24696};
  wire [1:0] _24698 = {_0, _8767} + {_0, _10910};
  wire [3:0] _24699 = {_0, _24697} + {_0, _0, _24698};
  wire _24700 = _12301 < _24699;
  wire _24701 = r670 ^ _24700;
  wire _24702 = _12298 ? coded_block[670] : r670;
  wire _24703 = _12296 ? _24701 : _24702;
  always @ (posedge reset or posedge clock) if (reset) r670 <= 1'd0; else if (_12300) r670 <= _24703;
  wire [1:0] _24704 = {_0, _831} + {_0, _3615};
  wire [1:0] _24705 = {_0, _5981} + {_0, _6462};
  wire [2:0] _24706 = {_0, _24704} + {_0, _24705};
  wire [1:0] _24707 = {_0, _9886} + {_0, _10846};
  wire [3:0] _24708 = {_0, _24706} + {_0, _0, _24707};
  wire _24709 = _12301 < _24708;
  wire _24710 = r669 ^ _24709;
  wire _24711 = _12298 ? coded_block[669] : r669;
  wire _24712 = _12296 ? _24710 : _24711;
  always @ (posedge reset or posedge clock) if (reset) r669 <= 1'd0; else if (_12300) r669 <= _24712;
  wire [1:0] _24713 = {_0, _34} + {_0, _3167};
  wire [1:0] _24714 = {_0, _5246} + {_0, _7326};
  wire [2:0] _24715 = {_0, _24713} + {_0, _24714};
  wire [1:0] _24716 = {_0, _9406} + {_0, _11485};
  wire [3:0] _24717 = {_0, _24715} + {_0, _0, _24716};
  wire _24718 = _12301 < _24717;
  wire _24719 = r668 ^ _24718;
  wire _24720 = _12298 ? coded_block[668] : r668;
  wire _24721 = _12296 ? _24719 : _24720;
  always @ (posedge reset or posedge clock) if (reset) r668 <= 1'd0; else if (_12300) r668 <= _24721;
  wire [1:0] _24722 = {_0, _161} + {_0, _3678};
  wire [1:0] _24723 = {_0, _5342} + {_0, _6397};
  wire [2:0] _24724 = {_0, _24722} + {_0, _24723};
  wire [1:0] _24725 = {_0, _8863} + {_0, _11389};
  wire [3:0] _24726 = {_0, _24724} + {_0, _0, _24725};
  wire _24727 = _12301 < _24726;
  wire _24728 = r667 ^ _24727;
  wire _24729 = _12298 ? coded_block[667] : r667;
  wire _24730 = _12296 ? _24728 : _24729;
  always @ (posedge reset or posedge clock) if (reset) r667 <= 1'd0; else if (_12300) r667 <= _24730;
  wire [1:0] _24731 = {_0, _192} + {_0, _2144};
  wire [1:0] _24732 = {_0, _5757} + {_0, _7420};
  wire [2:0] _24733 = {_0, _24731} + {_0, _24732};
  wire [1:0] _24734 = {_0, _8480} + {_0, _10941};
  wire [3:0] _24735 = {_0, _24733} + {_0, _0, _24734};
  wire _24736 = _12301 < _24735;
  wire _24737 = r666 ^ _24736;
  wire _24738 = _12298 ? coded_block[666] : r666;
  wire _24739 = _12296 ? _24737 : _24738;
  always @ (posedge reset or posedge clock) if (reset) r666 <= 1'd0; else if (_12300) r666 <= _24739;
  wire [1:0] _24740 = {_0, _224} + {_0, _3580};
  wire [1:0] _24741 = {_0, _4223} + {_0, _7837};
  wire [2:0] _24742 = {_0, _24740} + {_0, _24741};
  wire [1:0] _24743 = {_0, _9503} + {_0, _10558};
  wire [3:0] _24744 = {_0, _24742} + {_0, _0, _24743};
  wire _24745 = _12301 < _24744;
  wire _24746 = r665 ^ _24745;
  wire _24747 = _12298 ? coded_block[665] : r665;
  wire _24748 = _12296 ? _24746 : _24747;
  always @ (posedge reset or posedge clock) if (reset) r665 <= 1'd0; else if (_12300) r665 <= _24748;
  wire [1:0] _24749 = {_0, _255} + {_0, _2878};
  wire [1:0] _24750 = {_0, _5663} + {_0, _6303};
  wire [2:0] _24751 = {_0, _24749} + {_0, _24750};
  wire [1:0] _24752 = {_0, _9917} + {_0, _11581};
  wire [3:0] _24753 = {_0, _24751} + {_0, _0, _24752};
  wire _24754 = _12301 < _24753;
  wire _24755 = r664 ^ _24754;
  wire _24756 = _12298 ? coded_block[664] : r664;
  wire _24757 = _12296 ? _24755 : _24756;
  always @ (posedge reset or posedge clock) if (reset) r664 <= 1'd0; else if (_12300) r664 <= _24757;
  wire [1:0] _24758 = {_0, _320} + {_0, _2719};
  wire [1:0] _24759 = {_0, _4640} + {_0, _7036};
  wire [2:0] _24760 = {_0, _24758} + {_0, _24759};
  wire [1:0] _24761 = {_0, _9822} + {_0, _10462};
  wire [3:0] _24762 = {_0, _24760} + {_0, _0, _24761};
  wire _24763 = _12301 < _24762;
  wire _24764 = r663 ^ _24763;
  wire _24765 = _12298 ? coded_block[663] : r663;
  wire _24766 = _12296 ? _24764 : _24765;
  always @ (posedge reset or posedge clock) if (reset) r663 <= 1'd0; else if (_12300) r663 <= _24766;
  wire [1:0] _24767 = {_0, _352} + {_0, _2526};
  wire [1:0] _24768 = {_0, _4798} + {_0, _6718};
  wire [2:0] _24769 = {_0, _24767} + {_0, _24768};
  wire [1:0] _24770 = {_0, _9118} + {_0, _11900};
  wire [3:0] _24771 = {_0, _24769} + {_0, _0, _24770};
  wire _24772 = _12301 < _24771;
  wire _24773 = r662 ^ _24772;
  wire _24774 = _12298 ? coded_block[662] : r662;
  wire _24775 = _12296 ? _24773 : _24774;
  always @ (posedge reset or posedge clock) if (reset) r662 <= 1'd0; else if (_12300) r662 <= _24775;
  wire [1:0] _24776 = {_0, _383} + {_0, _2910};
  wire [1:0] _24777 = {_0, _4605} + {_0, _6877};
  wire [2:0] _24778 = {_0, _24776} + {_0, _24777};
  wire [1:0] _24779 = {_0, _8799} + {_0, _11196};
  wire [3:0] _24780 = {_0, _24778} + {_0, _0, _24779};
  wire _24781 = _12301 < _24780;
  wire _24782 = r661 ^ _24781;
  wire _24783 = _12298 ? coded_block[661] : r661;
  wire _24784 = _12296 ? _24782 : _24783;
  always @ (posedge reset or posedge clock) if (reset) r661 <= 1'd0; else if (_12300) r661 <= _24784;
  wire [1:0] _24785 = {_0, _416} + {_0, _4060};
  wire [1:0] _24786 = {_0, _4989} + {_0, _6687};
  wire [2:0] _24787 = {_0, _24785} + {_0, _24786};
  wire [1:0] _24788 = {_0, _8957} + {_0, _10877};
  wire [3:0] _24789 = {_0, _24787} + {_0, _0, _24788};
  wire _24790 = _12301 < _24789;
  wire _24791 = r660 ^ _24790;
  wire _24792 = _12298 ? coded_block[660] : r660;
  wire _24793 = _12296 ? _24791 : _24792;
  always @ (posedge reset or posedge clock) if (reset) r660 <= 1'd0; else if (_12300) r660 <= _24793;
  wire [1:0] _24794 = {_0, _447} + {_0, _3836};
  wire [1:0] _24795 = {_0, _6139} + {_0, _7069};
  wire [2:0] _24796 = {_0, _24794} + {_0, _24795};
  wire [1:0] _24797 = {_0, _8767} + {_0, _11038};
  wire [3:0] _24798 = {_0, _24796} + {_0, _0, _24797};
  wire _24799 = _12301 < _24798;
  wire _24800 = r659 ^ _24799;
  wire _24801 = _12298 ? coded_block[659] : r659;
  wire _24802 = _12296 ? _24800 : _24801;
  always @ (posedge reset or posedge clock) if (reset) r659 <= 1'd0; else if (_12300) r659 <= _24802;
  wire [1:0] _24803 = {_0, _479} + {_0, _2399};
  wire [1:0] _24804 = {_0, _5918} + {_0, _6207};
  wire [2:0] _24805 = {_0, _24803} + {_0, _24804};
  wire [1:0] _24806 = {_0, _9149} + {_0, _10846};
  wire [3:0] _24807 = {_0, _24805} + {_0, _0, _24806};
  wire _24808 = _12301 < _24807;
  wire _24809 = r658 ^ _24808;
  wire _24810 = _12298 ? coded_block[658] : r658;
  wire _24811 = _12296 ? _24809 : _24810;
  always @ (posedge reset or posedge clock) if (reset) r658 <= 1'd0; else if (_12300) r658 <= _24811;
  wire [1:0] _24812 = {_0, _510} + {_0, _2336};
  wire [1:0] _24813 = {_0, _4478} + {_0, _7996};
  wire [2:0] _24814 = {_0, _24812} + {_0, _24813};
  wire [1:0] _24815 = {_0, _8288} + {_0, _11228};
  wire [3:0] _24816 = {_0, _24814} + {_0, _0, _24815};
  wire _24817 = _12301 < _24816;
  wire _24818 = r657 ^ _24817;
  wire _24819 = _12298 ? coded_block[657] : r657;
  wire _24820 = _12296 ? _24818 : _24819;
  always @ (posedge reset or posedge clock) if (reset) r657 <= 1'd0; else if (_12300) r657 <= _24820;
  wire [1:0] _24821 = {_0, _545} + {_0, _3453};
  wire [1:0] _24822 = {_0, _4415} + {_0, _6558};
  wire [2:0] _24823 = {_0, _24821} + {_0, _24822};
  wire [1:0] _24824 = {_0, _10077} + {_0, _10366};
  wire [3:0] _24825 = {_0, _24823} + {_0, _0, _24824};
  wire _24826 = _12301 < _24825;
  wire _24827 = r656 ^ _24826;
  wire _24828 = _12298 ? coded_block[656] : r656;
  wire _24829 = _12296 ? _24827 : _24828;
  always @ (posedge reset or posedge clock) if (reset) r656 <= 1'd0; else if (_12300) r656 <= _24829;
  wire [1:0] _24830 = {_0, _576} + {_0, _2112};
  wire [1:0] _24831 = {_0, _5534} + {_0, _6494};
  wire [2:0] _24832 = {_0, _24830} + {_0, _24831};
  wire [1:0] _24833 = {_0, _8638} + {_0, _12155};
  wire [3:0] _24834 = {_0, _24832} + {_0, _0, _24833};
  wire _24835 = _12301 < _24834;
  wire _24836 = r655 ^ _24835;
  wire _24837 = _12298 ? coded_block[655] : r655;
  wire _24838 = _12296 ? _24836 : _24837;
  always @ (posedge reset or posedge clock) if (reset) r655 <= 1'd0; else if (_12300) r655 <= _24838;
  wire [1:0] _24839 = {_0, _608} + {_0, _3709};
  wire [1:0] _24840 = {_0, _4192} + {_0, _7612};
  wire [2:0] _24841 = {_0, _24839} + {_0, _24840};
  wire [1:0] _24842 = {_0, _8574} + {_0, _10717};
  wire [3:0] _24843 = {_0, _24841} + {_0, _0, _24842};
  wire _24844 = _12301 < _24843;
  wire _24845 = r654 ^ _24844;
  wire _24846 = _12298 ? coded_block[654] : r654;
  wire _24847 = _12296 ? _24845 : _24846;
  always @ (posedge reset or posedge clock) if (reset) r654 <= 1'd0; else if (_12300) r654 <= _24847;
  wire [1:0] _24848 = {_0, _703} + {_0, _3870};
  wire [1:0] _24849 = {_0, _4447} + {_0, _7581};
  wire [2:0] _24850 = {_0, _24848} + {_0, _24849};
  wire [1:0] _24851 = {_0, _9949} + {_0, _10430};
  wire [3:0] _24852 = {_0, _24850} + {_0, _0, _24851};
  wire _24853 = _12301 < _24852;
  wire _24854 = r653 ^ _24853;
  wire _24855 = _12298 ? coded_block[653] : r653;
  wire _24856 = _12296 ? _24854 : _24855;
  always @ (posedge reset or posedge clock) if (reset) r653 <= 1'd0; else if (_12300) r653 <= _24856;
  wire [1:0] _24857 = {_0, _766} + {_0, _3615};
  wire [1:0] _24858 = {_0, _4926} + {_0, _8028};
  wire [2:0] _24859 = {_0, _24857} + {_0, _24858};
  wire [1:0] _24860 = {_0, _8607} + {_0, _11740};
  wire [3:0] _24861 = {_0, _24859} + {_0, _0, _24860};
  wire _24862 = _12301 < _24861;
  wire _24863 = r652 ^ _24862;
  wire _24864 = _12298 ? coded_block[652] : r652;
  wire _24865 = _12296 ? _24863 : _24864;
  always @ (posedge reset or posedge clock) if (reset) r652 <= 1'd0; else if (_12300) r652 <= _24865;
  wire [1:0] _24866 = {_0, _800} + {_0, _2782};
  wire [1:0] _24867 = {_0, _5694} + {_0, _7005};
  wire [2:0] _24868 = {_0, _24866} + {_0, _24867};
  wire [1:0] _24869 = {_0, _10108} + {_0, _10685};
  wire [3:0] _24870 = {_0, _24868} + {_0, _0, _24869};
  wire _24871 = _12301 < _24870;
  wire _24872 = r651 ^ _24871;
  wire _24873 = _12298 ? coded_block[651] : r651;
  wire _24874 = _12296 ? _24872 : _24873;
  always @ (posedge reset or posedge clock) if (reset) r651 <= 1'd0; else if (_12300) r651 <= _24874;
  wire [1:0] _24875 = {_0, _831} + {_0, _2302};
  wire [1:0] _24876 = {_0, _4861} + {_0, _7773};
  wire [2:0] _24877 = {_0, _24875} + {_0, _24876};
  wire [1:0] _24878 = {_0, _9085} + {_0, _12188};
  wire [3:0] _24879 = {_0, _24877} + {_0, _0, _24878};
  wire _24880 = _12301 < _24879;
  wire _24881 = r650 ^ _24880;
  wire _24882 = _12298 ? coded_block[650] : r650;
  wire _24883 = _12296 ? _24881 : _24882;
  always @ (posedge reset or posedge clock) if (reset) r650 <= 1'd0; else if (_12300) r650 <= _24883;
  wire [1:0] _24884 = {_0, _863} + {_0, _2430};
  wire [1:0] _24885 = {_0, _4384} + {_0, _6942};
  wire [2:0] _24886 = {_0, _24884} + {_0, _24885};
  wire [1:0] _24887 = {_0, _9853} + {_0, _11165};
  wire [3:0] _24888 = {_0, _24886} + {_0, _0, _24887};
  wire _24889 = _12301 < _24888;
  wire _24890 = r649 ^ _24889;
  wire _24891 = _12298 ? coded_block[649] : r649;
  wire _24892 = _12296 ? _24890 : _24891;
  always @ (posedge reset or posedge clock) if (reset) r649 <= 1'd0; else if (_12300) r649 <= _24892;
  wire [1:0] _24893 = {_0, _894} + {_0, _3773};
  wire [1:0] _24894 = {_0, _4511} + {_0, _6462};
  wire [2:0] _24895 = {_0, _24893} + {_0, _24894};
  wire [1:0] _24896 = {_0, _9022} + {_0, _11933};
  wire [3:0] _24897 = {_0, _24895} + {_0, _0, _24896};
  wire _24898 = _12301 < _24897;
  wire _24899 = r648 ^ _24898;
  wire _24900 = _12298 ? coded_block[648] : r648;
  wire _24901 = _12296 ? _24899 : _24900;
  always @ (posedge reset or posedge clock) if (reset) r648 <= 1'd0; else if (_12300) r648 <= _24901;
  wire [1:0] _24902 = {_0, _927} + {_0, _3005};
  wire [1:0] _24903 = {_0, _5853} + {_0, _6589};
  wire [2:0] _24904 = {_0, _24902} + {_0, _24903};
  wire [1:0] _24905 = {_0, _8543} + {_0, _11101};
  wire [3:0] _24906 = {_0, _24904} + {_0, _0, _24905};
  wire _24907 = _12301 < _24906;
  wire _24908 = r647 ^ _24907;
  wire _24909 = _12298 ? coded_block[647] : r647;
  wire _24910 = _12296 ? _24908 : _24909;
  always @ (posedge reset or posedge clock) if (reset) r647 <= 1'd0; else if (_12300) r647 <= _24910;
  wire [1:0] _24911 = {_0, _958} + {_0, _2974};
  wire [1:0] _24912 = {_0, _5085} + {_0, _7931};
  wire [2:0] _24913 = {_0, _24911} + {_0, _24912};
  wire [1:0] _24914 = {_0, _8670} + {_0, _10621};
  wire [3:0] _24915 = {_0, _24913} + {_0, _0, _24914};
  wire _24916 = _12301 < _24915;
  wire _24917 = r646 ^ _24916;
  wire _24918 = _12298 ? coded_block[646] : r646;
  wire _24919 = _12296 ? _24917 : _24918;
  always @ (posedge reset or posedge clock) if (reset) r646 <= 1'd0; else if (_12300) r646 <= _24919;
  wire [1:0] _24920 = {_0, _990} + {_0, _3805};
  wire [1:0] _24921 = {_0, _5053} + {_0, _7163};
  wire [2:0] _24922 = {_0, _24920} + {_0, _24921};
  wire [1:0] _24923 = {_0, _10014} + {_0, _10748};
  wire [3:0] _24924 = {_0, _24922} + {_0, _0, _24923};
  wire _24925 = _12301 < _24924;
  wire _24926 = r645 ^ _24925;
  wire _24927 = _12298 ? coded_block[645] : r645;
  wire _24928 = _12296 ? _24926 : _24927;
  always @ (posedge reset or posedge clock) if (reset) r645 <= 1'd0; else if (_12300) r645 <= _24928;
  wire [1:0] _24929 = {_0, _1021} + {_0, _4091};
  wire [1:0] _24930 = {_0, _5884} + {_0, _7132};
  wire [2:0] _24931 = {_0, _24929} + {_0, _24930};
  wire [1:0] _24932 = {_0, _9248} + {_0, _12092};
  wire [3:0] _24933 = {_0, _24931} + {_0, _0, _24932};
  wire _24934 = _12301 < _24933;
  wire _24935 = r644 ^ _24934;
  wire _24936 = _12298 ? coded_block[644] : r644;
  wire _24937 = _12296 ? _24935 : _24936;
  always @ (posedge reset or posedge clock) if (reset) r644 <= 1'd0; else if (_12300) r644 <= _24937;
  wire [1:0] _24938 = {_0, _1057} + {_0, _3486};
  wire [1:0] _24939 = {_0, _4160} + {_0, _7965};
  wire [2:0] _24940 = {_0, _24938} + {_0, _24939};
  wire [1:0] _24941 = {_0, _9212} + {_0, _11326};
  wire [3:0] _24942 = {_0, _24940} + {_0, _0, _24941};
  wire _24943 = _12301 < _24942;
  wire _24944 = r643 ^ _24943;
  wire _24945 = _12298 ? coded_block[643] : r643;
  wire _24946 = _12296 ? _24944 : _24945;
  always @ (posedge reset or posedge clock) if (reset) r643 <= 1'd0; else if (_12300) r643 <= _24946;
  wire [1:0] _24947 = {_0, _1088} + {_0, _3325};
  wire [1:0] _24948 = {_0, _5565} + {_0, _6239};
  wire [2:0] _24949 = {_0, _24947} + {_0, _24948};
  wire [1:0] _24950 = {_0, _10045} + {_0, _11295};
  wire [3:0] _24951 = {_0, _24949} + {_0, _0, _24950};
  wire _24952 = _12301 < _24951;
  wire _24953 = r642 ^ _24952;
  wire _24954 = _12298 ? coded_block[642] : r642;
  wire _24955 = _12296 ? _24953 : _24954;
  always @ (posedge reset or posedge clock) if (reset) r642 <= 1'd0; else if (_12300) r642 <= _24955;
  wire [1:0] _24956 = {_0, _1120} + {_0, _2081};
  wire [1:0] _24957 = {_0, _5407} + {_0, _7644};
  wire [2:0] _24958 = {_0, _24956} + {_0, _24957};
  wire [1:0] _24959 = {_0, _8319} + {_0, _12124};
  wire [3:0] _24960 = {_0, _24958} + {_0, _0, _24959};
  wire _24961 = _12301 < _24960;
  wire _24962 = r641 ^ _24961;
  wire _24963 = _12298 ? coded_block[641] : r641;
  wire _24964 = _12296 ? _24962 : _24963;
  always @ (posedge reset or posedge clock) if (reset) r641 <= 1'd0; else if (_12300) r641 <= _24964;
  wire [1:0] _24965 = {_0, _1151} + {_0, _3359};
  wire [1:0] _24966 = {_0, _4129} + {_0, _7485};
  wire [2:0] _24967 = {_0, _24965} + {_0, _24966};
  wire [1:0] _24968 = {_0, _9724} + {_0, _10399};
  wire [3:0] _24969 = {_0, _24967} + {_0, _0, _24968};
  wire _24970 = _12301 < _24969;
  wire _24971 = r640 ^ _24970;
  wire _24972 = _12298 ? coded_block[640] : r640;
  wire _24973 = _12296 ? _24971 : _24972;
  always @ (posedge reset or posedge clock) if (reset) r640 <= 1'd0; else if (_12300) r640 <= _24973;
  wire [1:0] _24974 = {_0, _1184} + {_0, _3549};
  wire [1:0] _24975 = {_0, _5438} + {_0, _6176};
  wire [2:0] _24976 = {_0, _24974} + {_0, _24975};
  wire [1:0] _24977 = {_0, _9566} + {_0, _11806};
  wire [3:0] _24978 = {_0, _24976} + {_0, _0, _24977};
  wire _24979 = _12301 < _24978;
  wire _24980 = r639 ^ _24979;
  wire _24981 = _12298 ? coded_block[639] : r639;
  wire _24982 = _12296 ? _24980 : _24981;
  always @ (posedge reset or posedge clock) if (reset) r639 <= 1'd0; else if (_12300) r639 <= _24982;
  wire [1:0] _24983 = {_0, _1215} + {_0, _2175};
  wire [1:0] _24984 = {_0, _5628} + {_0, _7517};
  wire [2:0] _24985 = {_0, _24983} + {_0, _24984};
  wire [1:0] _24986 = {_0, _8225} + {_0, _11644};
  wire [3:0] _24987 = {_0, _24985} + {_0, _0, _24986};
  wire _24988 = _12301 < _24987;
  wire _24989 = r638 ^ _24988;
  wire _24990 = _12298 ? coded_block[638] : r638;
  wire _24991 = _12296 ? _24989 : _24990;
  always @ (posedge reset or posedge clock) if (reset) r638 <= 1'd0; else if (_12300) r638 <= _24991;
  wire [1:0] _24992 = {_0, _1247} + {_0, _3933};
  wire [1:0] _24993 = {_0, _4256} + {_0, _7710};
  wire [2:0] _24994 = {_0, _24992} + {_0, _24993};
  wire [1:0] _24995 = {_0, _9597} + {_0, _10272};
  wire [3:0] _24996 = {_0, _24994} + {_0, _0, _24995};
  wire _24997 = _12301 < _24996;
  wire _24998 = r637 ^ _24997;
  wire _24999 = _12298 ? coded_block[637] : r637;
  wire _25000 = _12296 ? _24998 : _24999;
  always @ (posedge reset or posedge clock) if (reset) r637 <= 1'd0; else if (_12300) r637 <= _25000;
  wire [1:0] _25001 = {_0, _1278} + {_0, _3135};
  wire [1:0] _25002 = {_0, _6012} + {_0, _6334};
  wire [2:0] _25003 = {_0, _25001} + {_0, _25002};
  wire [1:0] _25004 = {_0, _9790} + {_0, _11677};
  wire [3:0] _25005 = {_0, _25003} + {_0, _0, _25004};
  wire _25006 = _12301 < _25005;
  wire _25007 = r636 ^ _25006;
  wire _25008 = _12298 ? coded_block[636] : r636;
  wire _25009 = _12296 ? _25007 : _25008;
  always @ (posedge reset or posedge clock) if (reset) r636 <= 1'd0; else if (_12300) r636 <= _25009;
  wire [1:0] _25010 = {_0, _1312} + {_0, _3198};
  wire [1:0] _25011 = {_0, _5215} + {_0, _8092};
  wire [2:0] _25012 = {_0, _25010} + {_0, _25011};
  wire [1:0] _25013 = {_0, _8415} + {_0, _11869};
  wire [3:0] _25014 = {_0, _25012} + {_0, _0, _25013};
  wire _25015 = _12301 < _25014;
  wire _25016 = r635 ^ _25015;
  wire _25017 = _12298 ? coded_block[635] : r635;
  wire _25018 = _12296 ? _25016 : _25017;
  always @ (posedge reset or posedge clock) if (reset) r635 <= 1'd0; else if (_12300) r635 <= _25018;
  wire [1:0] _25019 = {_0, _1343} + {_0, _3997};
  wire [1:0] _25020 = {_0, _5279} + {_0, _7293};
  wire [2:0] _25021 = {_0, _25019} + {_0, _25020};
  wire [1:0] _25022 = {_0, _10172} + {_0, _10493};
  wire [3:0] _25023 = {_0, _25021} + {_0, _0, _25022};
  wire _25024 = _12301 < _25023;
  wire _25025 = r634 ^ _25024;
  wire _25026 = _12298 ? coded_block[634] : r634;
  wire _25027 = _12296 ? _25025 : _25026;
  always @ (posedge reset or posedge clock) if (reset) r634 <= 1'd0; else if (_12300) r634 <= _25027;
  wire [1:0] _25028 = {_0, _1375} + {_0, _2686};
  wire [1:0] _25029 = {_0, _6076} + {_0, _7357};
  wire [2:0] _25030 = {_0, _25028} + {_0, _25029};
  wire [1:0] _25031 = {_0, _9375} + {_0, _12251};
  wire [3:0] _25032 = {_0, _25030} + {_0, _0, _25031};
  wire _25033 = _12301 < _25032;
  wire _25034 = r633 ^ _25033;
  wire _25035 = _12298 ? coded_block[633] : r633;
  wire _25036 = _12296 ? _25034 : _25035;
  always @ (posedge reset or posedge clock) if (reset) r633 <= 1'd0; else if (_12300) r633 <= _25036;
  wire [1:0] _25037 = {_0, _1406} + {_0, _2592};
  wire [1:0] _25038 = {_0, _4767} + {_0, _8155};
  wire [2:0] _25039 = {_0, _25037} + {_0, _25038};
  wire [1:0] _25040 = {_0, _9438} + {_0, _11453};
  wire [3:0] _25041 = {_0, _25039} + {_0, _0, _25040};
  wire _25042 = _12301 < _25041;
  wire _25043 = r632 ^ _25042;
  wire _25044 = _12298 ? coded_block[632] : r632;
  wire _25045 = _12296 ? _25043 : _25044;
  always @ (posedge reset or posedge clock) if (reset) r632 <= 1'd0; else if (_12300) r632 <= _25045;
  wire [1:0] _25046 = {_0, _1439} + {_0, _3104};
  wire [1:0] _25047 = {_0, _4671} + {_0, _6845};
  wire [2:0] _25048 = {_0, _25046} + {_0, _25047};
  wire [1:0] _25049 = {_0, _10235} + {_0, _11516};
  wire [3:0] _25050 = {_0, _25048} + {_0, _0, _25049};
  wire _25051 = _12301 < _25050;
  wire _25052 = r631 ^ _25051;
  wire _25053 = _12298 ? coded_block[631] : r631;
  wire _25054 = _12296 ? _25052 : _25053;
  always @ (posedge reset or posedge clock) if (reset) r631 <= 1'd0; else if (_12300) r631 <= _25054;
  wire [1:0] _25055 = {_0, _1470} + {_0, _3964};
  wire [1:0] _25056 = {_0, _5183} + {_0, _6750};
  wire [2:0] _25057 = {_0, _25055} + {_0, _25056};
  wire [1:0] _25058 = {_0, _8926} + {_0, _10303};
  wire [3:0] _25059 = {_0, _25057} + {_0, _0, _25058};
  wire _25060 = _12301 < _25059;
  wire _25061 = r630 ^ _25060;
  wire _25062 = _12298 ? coded_block[630] : r630;
  wire _25063 = _12296 ? _25061 : _25062;
  always @ (posedge reset or posedge clock) if (reset) r630 <= 1'd0; else if (_12300) r630 <= _25063;
  wire [1:0] _25064 = {_0, _1533} + {_0, _2271};
  wire [1:0] _25065 = {_0, _5310} + {_0, _8123};
  wire [2:0] _25066 = {_0, _25064} + {_0, _25065};
  wire [1:0] _25067 = {_0, _9342} + {_0, _10910};
  wire [3:0] _25068 = {_0, _25066} + {_0, _0, _25067};
  wire _25069 = _12301 < _25068;
  wire _25070 = r629 ^ _25069;
  wire _25071 = _12298 ? coded_block[629] : r629;
  wire _25072 = _12296 ? _25070 : _25071;
  always @ (posedge reset or posedge clock) if (reset) r629 <= 1'd0; else if (_12300) r629 <= _25072;
  wire [1:0] _25073 = {_0, _1599} + {_0, _3901};
  wire [1:0] _25074 = {_0, _4895} + {_0, _6431};
  wire [2:0] _25075 = {_0, _25073} + {_0, _25074};
  wire [1:0] _25076 = {_0, _9469} + {_0, _12282};
  wire [3:0] _25077 = {_0, _25075} + {_0, _0, _25076};
  wire _25078 = _12301 < _25077;
  wire _25079 = r628 ^ _25078;
  wire _25080 = _12298 ? coded_block[628] : r628;
  wire _25081 = _12296 ? _25079 : _25080;
  always @ (posedge reset or posedge clock) if (reset) r628 <= 1'd0; else if (_12300) r628 <= _25081;
  wire [1:0] _25082 = {_0, _1631} + {_0, _2208};
  wire [1:0] _25083 = {_0, _5981} + {_0, _6973};
  wire [2:0] _25084 = {_0, _25082} + {_0, _25083};
  wire [1:0] _25085 = {_0, _8511} + {_0, _11550};
  wire [3:0] _25086 = {_0, _25084} + {_0, _0, _25085};
  wire _25087 = _12301 < _25086;
  wire _25088 = r627 ^ _25087;
  wire _25089 = _12298 ? coded_block[627] : r627;
  wire _25090 = _12296 ? _25088 : _25089;
  always @ (posedge reset or posedge clock) if (reset) r627 <= 1'd0; else if (_12300) r627 <= _25090;
  wire [1:0] _25091 = {_0, _1662} + {_0, _2655};
  wire [1:0] _25092 = {_0, _4287} + {_0, _8059};
  wire [2:0] _25093 = {_0, _25091} + {_0, _25092};
  wire [1:0] _25094 = {_0, _9054} + {_0, _10590};
  wire [3:0] _25095 = {_0, _25093} + {_0, _0, _25094};
  wire _25096 = _12301 < _25095;
  wire _25097 = r626 ^ _25096;
  wire _25098 = _12298 ? coded_block[626] : r626;
  wire _25099 = _12296 ? _25097 : _25098;
  always @ (posedge reset or posedge clock) if (reset) r626 <= 1'd0; else if (_12300) r626 <= _25099;
  wire [1:0] _25100 = {_0, _1695} + {_0, _4028};
  wire [1:0] _25101 = {_0, _4734} + {_0, _6366};
  wire [2:0] _25102 = {_0, _25100} + {_0, _25101};
  wire [1:0] _25103 = {_0, _10141} + {_0, _11132};
  wire [3:0] _25104 = {_0, _25102} + {_0, _0, _25103};
  wire _25105 = _12301 < _25104;
  wire _25106 = r625 ^ _25105;
  wire _25107 = _12298 ? coded_block[625] : r625;
  wire _25108 = _12296 ? _25106 : _25107;
  always @ (posedge reset or posedge clock) if (reset) r625 <= 1'd0; else if (_12300) r625 <= _25108;
  wire [1:0] _25109 = {_0, _1789} + {_0, _2494};
  wire [1:0] _25110 = {_0, _5116} + {_0, _7100};
  wire [2:0] _25111 = {_0, _25109} + {_0, _25110};
  wire [1:0] _25112 = {_0, _8256} + {_0, _10973};
  wire [3:0] _25113 = {_0, _25111} + {_0, _0, _25112};
  wire _25114 = _12301 < _25113;
  wire _25115 = r624 ^ _25114;
  wire _25116 = _12298 ? coded_block[624] : r624;
  wire _25117 = _12296 ? _25115 : _25116;
  always @ (posedge reset or posedge clock) if (reset) r624 <= 1'd0; else if (_12300) r624 <= _25117;
  wire [1:0] _25118 = {_0, _1823} + {_0, _2750};
  wire [1:0] _25119 = {_0, _4574} + {_0, _7199};
  wire [2:0] _25120 = {_0, _25118} + {_0, _25119};
  wire [1:0] _25121 = {_0, _9181} + {_0, _10335};
  wire [3:0] _25122 = {_0, _25120} + {_0, _0, _25121};
  wire _25123 = _12301 < _25122;
  wire _25124 = r623 ^ _25123;
  wire _25125 = _12298 ? coded_block[623] : r623;
  wire _25126 = _12296 ? _25124 : _25125;
  always @ (posedge reset or posedge clock) if (reset) r623 <= 1'd0; else if (_12300) r623 <= _25126;
  wire [1:0] _25127 = {_0, _1854} + {_0, _3646};
  wire [1:0] _25128 = {_0, _4830} + {_0, _6652};
  wire [2:0] _25129 = {_0, _25127} + {_0, _25128};
  wire [1:0] _25130 = {_0, _9279} + {_0, _11259};
  wire [3:0] _25131 = {_0, _25129} + {_0, _0, _25130};
  wire _25132 = _12301 < _25131;
  wire _25133 = r622 ^ _25132;
  wire _25134 = _12298 ? coded_block[622] : r622;
  wire _25135 = _12296 ? _25133 : _25134;
  always @ (posedge reset or posedge clock) if (reset) r622 <= 1'd0; else if (_12300) r622 <= _25135;
  wire [1:0] _25136 = {_0, _1886} + {_0, _3294};
  wire [1:0] _25137 = {_0, _5726} + {_0, _6908};
  wire [2:0] _25138 = {_0, _25136} + {_0, _25137};
  wire [1:0] _25139 = {_0, _8736} + {_0, _11358};
  wire [3:0] _25140 = {_0, _25138} + {_0, _0, _25139};
  wire _25141 = _12301 < _25140;
  wire _25142 = r621 ^ _25141;
  wire _25143 = _12298 ? coded_block[621] : r621;
  wire _25144 = _12296 ? _25142 : _25143;
  always @ (posedge reset or posedge clock) if (reset) r621 <= 1'd0; else if (_12300) r621 <= _25144;
  wire [1:0] _25145 = {_0, _1981} + {_0, _3742};
  wire [1:0] _25146 = {_0, _5470} + {_0, _7675};
  wire [2:0] _25147 = {_0, _25145} + {_0, _25146};
  wire [1:0] _25148 = {_0, _9534} + {_0, _11964};
  wire [3:0] _25149 = {_0, _25147} + {_0, _0, _25148};
  wire _25150 = _12301 < _25149;
  wire _25151 = r620 ^ _25150;
  wire _25152 = _12298 ? coded_block[620] : r620;
  wire _25153 = _12296 ? _25151 : _25152;
  always @ (posedge reset or posedge clock) if (reset) r620 <= 1'd0; else if (_12300) r620 <= _25153;
  wire [1:0] _25154 = {_0, _2013} + {_0, _2463};
  wire [1:0] _25155 = {_0, _5821} + {_0, _7548};
  wire [2:0] _25156 = {_0, _25154} + {_0, _25155};
  wire [1:0] _25157 = {_0, _9759} + {_0, _11613};
  wire [3:0] _25158 = {_0, _25156} + {_0, _0, _25157};
  wire _25159 = _12301 < _25158;
  wire _25160 = r619 ^ _25159;
  wire _25161 = _12298 ? coded_block[619] : r619;
  wire _25162 = _12296 ? _25160 : _25161;
  always @ (posedge reset or posedge clock) if (reset) r619 <= 1'd0; else if (_12300) r619 <= _25162;
  wire [1:0] _25163 = {_0, _2044} + {_0, _3068};
  wire [1:0] _25164 = {_0, _4542} + {_0, _7900};
  wire [2:0] _25165 = {_0, _25163} + {_0, _25164};
  wire [1:0] _25166 = {_0, _9630} + {_0, _11837};
  wire [3:0] _25167 = {_0, _25165} + {_0, _0, _25166};
  wire _25168 = _12301 < _25167;
  wire _25169 = r618 ^ _25168;
  wire _25170 = _12298 ? coded_block[618] : r618;
  wire _25171 = _12296 ? _25169 : _25170;
  always @ (posedge reset or posedge clock) if (reset) r618 <= 1'd0; else if (_12300) r618 <= _25171;
  wire [1:0] _25172 = {_0, _65} + {_0, _2623};
  wire [1:0] _25173 = {_0, _5152} + {_0, _6621};
  wire [2:0] _25174 = {_0, _25172} + {_0, _25173};
  wire [1:0] _25175 = {_0, _9980} + {_0, _11708};
  wire [3:0] _25176 = {_0, _25174} + {_0, _0, _25175};
  wire _25177 = _12301 < _25176;
  wire _25178 = r617 ^ _25177;
  wire _25179 = _12298 ? coded_block[617] : r617;
  wire _25180 = _12296 ? _25178 : _25179;
  always @ (posedge reset or posedge clock) if (reset) r617 <= 1'd0; else if (_12300) r617 <= _25180;
  wire [1:0] _25181 = {_0, _34} + {_0, _2847};
  wire [1:0] _25182 = {_0, _4926} + {_0, _7005};
  wire [2:0] _25183 = {_0, _25181} + {_0, _25182};
  wire [1:0] _25184 = {_0, _9085} + {_0, _11165};
  wire [3:0] _25185 = {_0, _25183} + {_0, _0, _25184};
  wire _25186 = _12301 < _25185;
  wire _25187 = r616 ^ _25186;
  wire _25188 = _12298 ? coded_block[616] : r616;
  wire _25189 = _12296 ? _25187 : _25188;
  always @ (posedge reset or posedge clock) if (reset) r616 <= 1'd0; else if (_12300) r616 <= _25189;
  wire [1:0] _25190 = {_0, _1502} + {_0, _2430};
  wire [1:0] _25191 = {_0, _4256} + {_0, _6877};
  wire [2:0] _25192 = {_0, _25190} + {_0, _25191};
  wire [1:0] _25193 = {_0, _8863} + {_0, _12027};
  wire [3:0] _25194 = {_0, _25192} + {_0, _0, _25193};
  wire _25195 = _12301 < _25194;
  wire _25196 = r615 ^ _25195;
  wire _25197 = _12298 ? coded_block[615] : r615;
  wire _25198 = _12296 ? _25196 : _25197;
  always @ (posedge reset or posedge clock) if (reset) r615 <= 1'd0; else if (_12300) r615 <= _25198;
  wire [1:0] _25199 = {_0, _1533} + {_0, _3325};
  wire [1:0] _25200 = {_0, _4511} + {_0, _6334};
  wire [2:0] _25201 = {_0, _25199} + {_0, _25200};
  wire [1:0] _25202 = {_0, _8957} + {_0, _10941};
  wire [3:0] _25203 = {_0, _25201} + {_0, _0, _25202};
  wire _25204 = _12301 < _25203;
  wire _25205 = r614 ^ _25204;
  wire _25206 = _12298 ? coded_block[614] : r614;
  wire _25207 = _12296 ? _25205 : _25206;
  always @ (posedge reset or posedge clock) if (reset) r614 <= 1'd0; else if (_12300) r614 <= _25207;
  wire [1:0] _25208 = {_0, _1568} + {_0, _2974};
  wire [1:0] _25209 = {_0, _5407} + {_0, _6589};
  wire [2:0] _25210 = {_0, _25208} + {_0, _25209};
  wire [1:0] _25211 = {_0, _8415} + {_0, _11038};
  wire [3:0] _25212 = {_0, _25210} + {_0, _0, _25211};
  wire _25213 = _12301 < _25212;
  wire _25214 = r613 ^ _25213;
  wire _25215 = _12298 ? coded_block[613] : r613;
  wire _25216 = _12296 ? _25214 : _25215;
  always @ (posedge reset or posedge clock) if (reset) r613 <= 1'd0; else if (_12300) r613 <= _25216;
  wire [1:0] _25217 = {_0, _1599} + {_0, _3198};
  wire [1:0] _25218 = {_0, _5053} + {_0, _7485};
  wire [2:0] _25219 = {_0, _25217} + {_0, _25218};
  wire [1:0] _25220 = {_0, _8670} + {_0, _10493};
  wire [3:0] _25221 = {_0, _25219} + {_0, _0, _25220};
  wire _25222 = _12301 < _25221;
  wire _25223 = r612 ^ _25222;
  wire _25224 = _12298 ? coded_block[612] : r612;
  wire _25225 = _12296 ? _25223 : _25224;
  always @ (posedge reset or posedge clock) if (reset) r612 <= 1'd0; else if (_12300) r612 <= _25225;
  wire [1:0] _25226 = {_0, _1631} + {_0, _3068};
  wire [1:0] _25227 = {_0, _5279} + {_0, _7132};
  wire [2:0] _25228 = {_0, _25226} + {_0, _25227};
  wire [1:0] _25229 = {_0, _9566} + {_0, _10748};
  wire [3:0] _25230 = {_0, _25228} + {_0, _0, _25229};
  wire _25231 = _12301 < _25230;
  wire _25232 = r611 ^ _25231;
  wire _25233 = _12298 ? coded_block[611] : r611;
  wire _25234 = _12296 ? _25232 : _25233;
  always @ (posedge reset or posedge clock) if (reset) r611 <= 1'd0; else if (_12300) r611 <= _25234;
  wire [1:0] _25235 = {_0, _1662} + {_0, _3422};
  wire [1:0] _25236 = {_0, _5152} + {_0, _7357};
  wire [2:0] _25237 = {_0, _25235} + {_0, _25236};
  wire [1:0] _25238 = {_0, _9212} + {_0, _11644};
  wire [3:0] _25239 = {_0, _25237} + {_0, _0, _25238};
  wire _25240 = _12301 < _25239;
  wire _25241 = r610 ^ _25240;
  wire _25242 = _12298 ? coded_block[610] : r610;
  wire _25243 = _12296 ? _25241 : _25242;
  always @ (posedge reset or posedge clock) if (reset) r610 <= 1'd0; else if (_12300) r610 <= _25243;
  wire [1:0] _25244 = {_0, _1695} + {_0, _2144};
  wire [1:0] _25245 = {_0, _5501} + {_0, _7230};
  wire [2:0] _25246 = {_0, _25244} + {_0, _25245};
  wire [1:0] _25247 = {_0, _9438} + {_0, _11295};
  wire [3:0] _25248 = {_0, _25246} + {_0, _0, _25247};
  wire _25249 = _12301 < _25248;
  wire _25250 = r609 ^ _25249;
  wire _25251 = _12298 ? coded_block[609] : r609;
  wire _25252 = _12296 ? _25250 : _25251;
  always @ (posedge reset or posedge clock) if (reset) r609 <= 1'd0; else if (_12300) r609 <= _25252;
  wire [1:0] _25253 = {_0, _1726} + {_0, _2750};
  wire [1:0] _25254 = {_0, _4223} + {_0, _7581};
  wire [2:0] _25255 = {_0, _25253} + {_0, _25254};
  wire [1:0] _25256 = {_0, _9311} + {_0, _11516};
  wire [3:0] _25257 = {_0, _25255} + {_0, _0, _25256};
  wire _25258 = _12301 < _25257;
  wire _25259 = r608 ^ _25258;
  wire _25260 = _12298 ? coded_block[608] : r608;
  wire _25261 = _12296 ? _25259 : _25260;
  always @ (posedge reset or posedge clock) if (reset) r608 <= 1'd0; else if (_12300) r608 <= _25261;
  wire [1:0] _25262 = {_0, _1789} + {_0, _3933};
  wire [1:0] _25263 = {_0, _4384} + {_0, _6908};
  wire [2:0] _25264 = {_0, _25262} + {_0, _25263};
  wire [1:0] _25265 = {_0, _8383} + {_0, _11740};
  wire [3:0] _25266 = {_0, _25264} + {_0, _0, _25265};
  wire _25267 = _12301 < _25266;
  wire _25268 = r607 ^ _25267;
  wire _25269 = _12298 ? coded_block[607] : r607;
  wire _25270 = _12296 ? _25268 : _25269;
  always @ (posedge reset or posedge clock) if (reset) r607 <= 1'd0; else if (_12300) r607 <= _25270;
  wire [1:0] _25271 = {_0, _1823} + {_0, _2941};
  wire [1:0] _25272 = {_0, _6012} + {_0, _6462};
  wire [2:0] _25273 = {_0, _25271} + {_0, _25272};
  wire [1:0] _25274 = {_0, _8991} + {_0, _10462};
  wire [3:0] _25275 = {_0, _25273} + {_0, _0, _25274};
  wire _25276 = _12301 < _25275;
  wire _25277 = r606 ^ _25276;
  wire _25278 = _12298 ? coded_block[606] : r606;
  wire _25279 = _12296 ? _25277 : _25278;
  always @ (posedge reset or posedge clock) if (reset) r606 <= 1'd0; else if (_12300) r606 <= _25279;
  wire [1:0] _25280 = {_0, _1854} + {_0, _3359};
  wire [1:0] _25281 = {_0, _5022} + {_0, _8092};
  wire [2:0] _25282 = {_0, _25280} + {_0, _25281};
  wire [1:0] _25283 = {_0, _8543} + {_0, _11069};
  wire [3:0] _25284 = {_0, _25282} + {_0, _0, _25283};
  wire _25285 = _12301 < _25284;
  wire _25286 = r605 ^ _25285;
  wire _25287 = _12298 ? coded_block[605] : r605;
  wire _25288 = _12296 ? _25286 : _25287;
  always @ (posedge reset or posedge clock) if (reset) r605 <= 1'd0; else if (_12300) r605 <= _25288;
  wire [1:0] _25289 = {_0, _1886} + {_0, _3836};
  wire [1:0] _25290 = {_0, _5438} + {_0, _7100};
  wire [2:0] _25291 = {_0, _25289} + {_0, _25290};
  wire [1:0] _25292 = {_0, _10172} + {_0, _10621};
  wire [3:0] _25293 = {_0, _25291} + {_0, _0, _25292};
  wire _25294 = _12301 < _25293;
  wire _25295 = r604 ^ _25294;
  wire _25296 = _12298 ? coded_block[604] : r604;
  wire _25297 = _12296 ? _25295 : _25296;
  always @ (posedge reset or posedge clock) if (reset) r604 <= 1'd0; else if (_12300) r604 <= _25297;
  wire [1:0] _25298 = {_0, _1917} + {_0, _3262};
  wire [1:0] _25299 = {_0, _5918} + {_0, _7517};
  wire [2:0] _25300 = {_0, _25298} + {_0, _25299};
  wire [1:0] _25301 = {_0, _9181} + {_0, _12251};
  wire [3:0] _25302 = {_0, _25300} + {_0, _0, _25301};
  wire _25303 = _12301 < _25302;
  wire _25304 = r603 ^ _25303;
  wire _25305 = _12298 ? coded_block[603] : r603;
  wire _25306 = _12296 ? _25304 : _25305;
  always @ (posedge reset or posedge clock) if (reset) r603 <= 1'd0; else if (_12300) r603 <= _25306;
  wire [1:0] _25307 = {_0, _1981} + {_0, _2239};
  wire [1:0] _25308 = {_0, _4640} + {_0, _7420};
  wire [2:0] _25309 = {_0, _25307} + {_0, _25308};
  wire [1:0] _25310 = {_0, _10077} + {_0, _11677};
  wire [3:0] _25311 = {_0, _25309} + {_0, _0, _25310};
  wire _25312 = _12301 < _25311;
  wire _25313 = r602 ^ _25312;
  wire _25314 = _12298 ? coded_block[602] : r602;
  wire _25315 = _12296 ? _25313 : _25314;
  always @ (posedge reset or posedge clock) if (reset) r602 <= 1'd0; else if (_12300) r602 <= _25315;
  wire [1:0] _25316 = {_0, _2044} + {_0, _2208};
  wire [1:0] _25317 = {_0, _4478} + {_0, _6397};
  wire [2:0] _25318 = {_0, _25316} + {_0, _25317};
  wire [1:0] _25319 = {_0, _8799} + {_0, _11581};
  wire [3:0] _25320 = {_0, _25318} + {_0, _0, _25319};
  wire _25321 = _12301 < _25320;
  wire _25322 = r601 ^ _25321;
  wire _25323 = _12298 ? coded_block[601] : r601;
  wire _25324 = _12296 ? _25322 : _25323;
  always @ (posedge reset or posedge clock) if (reset) r601 <= 1'd0; else if (_12300) r601 <= _25324;
  wire [1:0] _25325 = {_0, _65} + {_0, _2592};
  wire [1:0] _25326 = {_0, _4287} + {_0, _6558};
  wire [2:0] _25327 = {_0, _25325} + {_0, _25326};
  wire [1:0] _25328 = {_0, _8480} + {_0, _10877};
  wire [3:0] _25329 = {_0, _25327} + {_0, _0, _25328};
  wire _25330 = _12301 < _25329;
  wire _25331 = r600 ^ _25330;
  wire _25332 = _12298 ? coded_block[600] : r600;
  wire _25333 = _12296 ? _25331 : _25332;
  always @ (posedge reset or posedge clock) if (reset) r600 <= 1'd0; else if (_12300) r600 <= _25333;
  wire [1:0] _25334 = {_0, _97} + {_0, _3742};
  wire [1:0] _25335 = {_0, _4671} + {_0, _6366};
  wire [2:0] _25336 = {_0, _25334} + {_0, _25335};
  wire [1:0] _25337 = {_0, _8638} + {_0, _10558};
  wire [3:0] _25338 = {_0, _25336} + {_0, _0, _25337};
  wire _25339 = _12301 < _25338;
  wire _25340 = r599 ^ _25339;
  wire _25341 = _12298 ? coded_block[599] : r599;
  wire _25342 = _12296 ? _25340 : _25341;
  always @ (posedge reset or posedge clock) if (reset) r599 <= 1'd0; else if (_12300) r599 <= _25342;
  wire [1:0] _25343 = {_0, _128} + {_0, _3517};
  wire [1:0] _25344 = {_0, _5821} + {_0, _6750};
  wire [2:0] _25345 = {_0, _25343} + {_0, _25344};
  wire [1:0] _25346 = {_0, _8446} + {_0, _10717};
  wire [3:0] _25347 = {_0, _25345} + {_0, _0, _25346};
  wire _25348 = _12301 < _25347;
  wire _25349 = r598 ^ _25348;
  wire _25350 = _12298 ? coded_block[598] : r598;
  wire _25351 = _12296 ? _25349 : _25350;
  always @ (posedge reset or posedge clock) if (reset) r598 <= 1'd0; else if (_12300) r598 <= _25351;
  wire [1:0] _25352 = {_0, _161} + {_0, _4091};
  wire [1:0] _25353 = {_0, _5597} + {_0, _7900};
  wire [2:0] _25354 = {_0, _25352} + {_0, _25353};
  wire [1:0] _25355 = {_0, _8830} + {_0, _10527};
  wire [3:0] _25356 = {_0, _25354} + {_0, _0, _25355};
  wire _25357 = _12301 < _25356;
  wire _25358 = r597 ^ _25357;
  wire _25359 = _12298 ? coded_block[597] : r597;
  wire _25360 = _12296 ? _25358 : _25359;
  always @ (posedge reset or posedge clock) if (reset) r597 <= 1'd0; else if (_12300) r597 <= _25360;
  wire [1:0] _25361 = {_0, _192} + {_0, _4028};
  wire [1:0] _25362 = {_0, _4160} + {_0, _7675};
  wire [2:0] _25363 = {_0, _25361} + {_0, _25362};
  wire [1:0] _25364 = {_0, _9980} + {_0, _10910};
  wire [3:0] _25365 = {_0, _25363} + {_0, _0, _25364};
  wire _25366 = _12301 < _25365;
  wire _25367 = r596 ^ _25366;
  wire _25368 = _12298 ? coded_block[596] : r596;
  wire _25369 = _12296 ? _25367 : _25368;
  always @ (posedge reset or posedge clock) if (reset) r596 <= 1'd0; else if (_12300) r596 <= _25369;
  wire [1:0] _25370 = {_0, _224} + {_0, _3135};
  wire [1:0] _25371 = {_0, _6108} + {_0, _6239};
  wire [2:0] _25372 = {_0, _25370} + {_0, _25371};
  wire [1:0] _25373 = {_0, _9759} + {_0, _12061};
  wire [3:0] _25374 = {_0, _25372} + {_0, _0, _25373};
  wire _25375 = _12301 < _25374;
  wire _25376 = r595 ^ _25375;
  wire _25377 = _12298 ? coded_block[595] : r595;
  wire _25378 = _12296 ? _25376 : _25377;
  always @ (posedge reset or posedge clock) if (reset) r595 <= 1'd0; else if (_12300) r595 <= _25378;
  wire [1:0] _25379 = {_0, _255} + {_0, _3805};
  wire [1:0] _25380 = {_0, _5215} + {_0, _8186};
  wire [2:0] _25381 = {_0, _25379} + {_0, _25380};
  wire [1:0] _25382 = {_0, _8319} + {_0, _11837};
  wire [3:0] _25383 = {_0, _25381} + {_0, _0, _25382};
  wire _25384 = _12301 < _25383;
  wire _25385 = r594 ^ _25384;
  wire _25386 = _12298 ? coded_block[594] : r594;
  wire _25387 = _12296 ? _25385 : _25386;
  always @ (posedge reset or posedge clock) if (reset) r594 <= 1'd0; else if (_12300) r594 <= _25387;
  wire [1:0] _25388 = {_0, _289} + {_0, _3390};
  wire [1:0] _25389 = {_0, _5884} + {_0, _7293};
  wire [2:0] _25390 = {_0, _25388} + {_0, _25389};
  wire [1:0] _25391 = {_0, _8256} + {_0, _10399};
  wire [3:0] _25392 = {_0, _25390} + {_0, _0, _25391};
  wire _25393 = _12301 < _25392;
  wire _25394 = r593 ^ _25393;
  wire _25395 = _12298 ? coded_block[593] : r593;
  wire _25396 = _12296 ? _25394 : _25395;
  always @ (posedge reset or posedge clock) if (reset) r593 <= 1'd0; else if (_12300) r593 <= _25396;
  wire [1:0] _25397 = {_0, _320} + {_0, _3104};
  wire [1:0] _25398 = {_0, _5470} + {_0, _7965};
  wire [2:0] _25399 = {_0, _25397} + {_0, _25398};
  wire [1:0] _25400 = {_0, _9375} + {_0, _10335};
  wire [3:0] _25401 = {_0, _25399} + {_0, _0, _25400};
  wire _25402 = _12301 < _25401;
  wire _25403 = r592 ^ _25402;
  wire _25404 = _12298 ? coded_block[592] : r592;
  wire _25405 = _12296 ? _25403 : _25404;
  always @ (posedge reset or posedge clock) if (reset) r592 <= 1'd0; else if (_12300) r592 <= _25405;
  wire [1:0] _25406 = {_0, _383} + {_0, _3549};
  wire [1:0] _25407 = {_0, _6139} + {_0, _7262};
  wire [2:0] _25408 = {_0, _25406} + {_0, _25407};
  wire [1:0] _25409 = {_0, _9630} + {_0, _12124};
  wire [3:0] _25410 = {_0, _25408} + {_0, _0, _25409};
  wire _25411 = _12301 < _25410;
  wire _25412 = r591 ^ _25411;
  wire _25413 = _12298 ? coded_block[591] : r591;
  wire _25414 = _12296 ? _25412 : _25413;
  always @ (posedge reset or posedge clock) if (reset) r591 <= 1'd0; else if (_12300) r591 <= _25414;
  wire [1:0] _25415 = {_0, _416} + {_0, _2526};
  wire [1:0] _25416 = {_0, _5628} + {_0, _6207};
  wire [2:0] _25417 = {_0, _25415} + {_0, _25416};
  wire [1:0] _25418 = {_0, _9342} + {_0, _11708};
  wire [3:0] _25419 = {_0, _25417} + {_0, _0, _25418};
  wire _25420 = _12301 < _25419;
  wire _25421 = r590 ^ _25420;
  wire _25422 = _12298 ? coded_block[590] : r590;
  wire _25423 = _12296 ? _25421 : _25422;
  always @ (posedge reset or posedge clock) if (reset) r590 <= 1'd0; else if (_12300) r590 <= _25423;
  wire [1:0] _25424 = {_0, _447} + {_0, _3294};
  wire [1:0] _25425 = {_0, _4605} + {_0, _7710};
  wire [2:0] _25426 = {_0, _25424} + {_0, _25425};
  wire [1:0] _25427 = {_0, _8288} + {_0, _11422};
  wire [3:0] _25428 = {_0, _25426} + {_0, _0, _25427};
  wire _25429 = _12301 < _25428;
  wire _25430 = r589 ^ _25429;
  wire _25431 = _12298 ? coded_block[589] : r589;
  wire _25432 = _12296 ? _25430 : _25431;
  always @ (posedge reset or posedge clock) if (reset) r589 <= 1'd0; else if (_12300) r589 <= _25432;
  wire [1:0] _25433 = {_0, _479} + {_0, _2463};
  wire [1:0] _25434 = {_0, _5373} + {_0, _6687};
  wire [2:0] _25435 = {_0, _25433} + {_0, _25434};
  wire [1:0] _25436 = {_0, _9790} + {_0, _10366};
  wire [3:0] _25437 = {_0, _25435} + {_0, _0, _25436};
  wire _25438 = _12301 < _25437;
  wire _25439 = r588 ^ _25438;
  wire _25440 = _12298 ? coded_block[588] : r588;
  wire _25441 = _12296 ? _25439 : _25440;
  always @ (posedge reset or posedge clock) if (reset) r588 <= 1'd0; else if (_12300) r588 <= _25441;
  wire [1:0] _25442 = {_0, _545} + {_0, _2112};
  wire [1:0] _25443 = {_0, _6076} + {_0, _6621};
  wire [2:0] _25444 = {_0, _25442} + {_0, _25443};
  wire [1:0] _25445 = {_0, _9534} + {_0, _10846};
  wire [3:0] _25446 = {_0, _25444} + {_0, _0, _25445};
  wire _25447 = _12301 < _25446;
  wire _25448 = r587 ^ _25447;
  wire _25449 = _12298 ? coded_block[587] : r587;
  wire _25450 = _12296 ? _25448 : _25449;
  always @ (posedge reset or posedge clock) if (reset) r587 <= 1'd0; else if (_12300) r587 <= _25450;
  wire [1:0] _25451 = {_0, _576} + {_0, _3453};
  wire [1:0] _25452 = {_0, _4192} + {_0, _8155};
  wire [2:0] _25453 = {_0, _25451} + {_0, _25452};
  wire [1:0] _25454 = {_0, _8701} + {_0, _11613};
  wire [3:0] _25455 = {_0, _25453} + {_0, _0, _25454};
  wire _25456 = _12301 < _25455;
  wire _25457 = r586 ^ _25456;
  wire _25458 = _12298 ? coded_block[586] : r586;
  wire _25459 = _12296 ? _25457 : _25458;
  always @ (posedge reset or posedge clock) if (reset) r586 <= 1'd0; else if (_12300) r586 <= _25459;
  wire [1:0] _25460 = {_0, _608} + {_0, _2686};
  wire [1:0] _25461 = {_0, _5534} + {_0, _6270};
  wire [2:0] _25462 = {_0, _25460} + {_0, _25461};
  wire [1:0] _25463 = {_0, _10235} + {_0, _10783};
  wire [3:0] _25464 = {_0, _25462} + {_0, _0, _25463};
  wire _25465 = _12301 < _25464;
  wire _25466 = r585 ^ _25465;
  wire _25467 = _12298 ? coded_block[585] : r585;
  wire _25468 = _12296 ? _25466 : _25467;
  always @ (posedge reset or posedge clock) if (reset) r585 <= 1'd0; else if (_12300) r585 <= _25468;
  wire [1:0] _25469 = {_0, _639} + {_0, _2655};
  wire [1:0] _25470 = {_0, _4767} + {_0, _7612};
  wire [2:0] _25471 = {_0, _25469} + {_0, _25470};
  wire [1:0] _25472 = {_0, _8352} + {_0, _10303};
  wire [3:0] _25473 = {_0, _25471} + {_0, _0, _25472};
  wire _25474 = _12301 < _25473;
  wire _25475 = r584 ^ _25474;
  wire _25476 = _12298 ? coded_block[584] : r584;
  wire _25477 = _12296 ? _25475 : _25476;
  always @ (posedge reset or posedge clock) if (reset) r584 <= 1'd0; else if (_12300) r584 <= _25477;
  wire [1:0] _25478 = {_0, _672} + {_0, _3486};
  wire [1:0] _25479 = {_0, _4734} + {_0, _6845};
  wire [2:0] _25480 = {_0, _25478} + {_0, _25479};
  wire [1:0] _25481 = {_0, _9693} + {_0, _10430};
  wire [3:0] _25482 = {_0, _25480} + {_0, _0, _25481};
  wire _25483 = _12301 < _25482;
  wire _25484 = r583 ^ _25483;
  wire _25485 = _12298 ? coded_block[583] : r583;
  wire _25486 = _12296 ? _25484 : _25485;
  always @ (posedge reset or posedge clock) if (reset) r583 <= 1'd0; else if (_12300) r583 <= _25486;
  wire [1:0] _25487 = {_0, _735} + {_0, _3167};
  wire [1:0] _25488 = {_0, _5853} + {_0, _7644};
  wire [2:0] _25489 = {_0, _25487} + {_0, _25488};
  wire [1:0] _25490 = {_0, _8894} + {_0, _11004};
  wire [3:0] _25491 = {_0, _25489} + {_0, _0, _25490};
  wire _25492 = _12301 < _25491;
  wire _25493 = r582 ^ _25492;
  wire _25494 = _12298 ? coded_block[582] : r582;
  wire _25495 = _12296 ? _25493 : _25494;
  always @ (posedge reset or posedge clock) if (reset) r582 <= 1'd0; else if (_12300) r582 <= _25495;
  wire [1:0] _25496 = {_0, _766} + {_0, _3005};
  wire [1:0] _25497 = {_0, _5246} + {_0, _7931};
  wire [2:0] _25498 = {_0, _25496} + {_0, _25497};
  wire [1:0] _25499 = {_0, _9724} + {_0, _10973};
  wire [3:0] _25500 = {_0, _25498} + {_0, _0, _25499};
  wire _25501 = _12301 < _25500;
  wire _25502 = r581 ^ _25501;
  wire _25503 = _12298 ? coded_block[581] : r581;
  wire _25504 = _12296 ? _25502 : _25503;
  always @ (posedge reset or posedge clock) if (reset) r581 <= 1'd0; else if (_12300) r581 <= _25504;
  wire [1:0] _25505 = {_0, _800} + {_0, _2081};
  wire [1:0] _25506 = {_0, _5085} + {_0, _7326};
  wire [2:0] _25507 = {_0, _25505} + {_0, _25506};
  wire [1:0] _25508 = {_0, _10014} + {_0, _11806};
  wire [3:0] _25509 = {_0, _25507} + {_0, _0, _25508};
  wire _25510 = _12301 < _25509;
  wire _25511 = r580 ^ _25510;
  wire _25512 = _12298 ? coded_block[580] : r580;
  wire _25513 = _12296 ? _25511 : _25512;
  always @ (posedge reset or posedge clock) if (reset) r580 <= 1'd0; else if (_12300) r580 <= _25513;
  wire [1:0] _25514 = {_0, _831} + {_0, _3037};
  wire [1:0] _25515 = {_0, _4129} + {_0, _7163};
  wire [2:0] _25516 = {_0, _25514} + {_0, _25515};
  wire [1:0] _25517 = {_0, _9406} + {_0, _12092};
  wire [3:0] _25518 = {_0, _25516} + {_0, _0, _25517};
  wire _25519 = _12301 < _25518;
  wire _25520 = r579 ^ _25519;
  wire _25521 = _12298 ? coded_block[579] : r579;
  wire _25522 = _12296 ? _25520 : _25521;
  always @ (posedge reset or posedge clock) if (reset) r579 <= 1'd0; else if (_12300) r579 <= _25522;
  wire [1:0] _25523 = {_0, _863} + {_0, _3231};
  wire [1:0] _25524 = {_0, _5116} + {_0, _6176};
  wire [2:0] _25525 = {_0, _25523} + {_0, _25524};
  wire [1:0] _25526 = {_0, _9248} + {_0, _11485};
  wire [3:0] _25527 = {_0, _25525} + {_0, _0, _25526};
  wire _25528 = _12301 < _25527;
  wire _25529 = r578 ^ _25528;
  wire _25530 = _12298 ? coded_block[578] : r578;
  wire _25531 = _12296 ? _25529 : _25530;
  always @ (posedge reset or posedge clock) if (reset) r578 <= 1'd0; else if (_12300) r578 <= _25531;
  wire [1:0] _25532 = {_0, _927} + {_0, _3615};
  wire [1:0] _25533 = {_0, _5949} + {_0, _7389};
  wire [2:0] _25534 = {_0, _25532} + {_0, _25533};
  wire [1:0] _25535 = {_0, _9279} + {_0, _10272};
  wire [3:0] _25536 = {_0, _25534} + {_0, _0, _25535};
  wire _25537 = _12301 < _25536;
  wire _25538 = r577 ^ _25537;
  wire _25539 = _12298 ? coded_block[577] : r577;
  wire _25540 = _12296 ? _25538 : _25539;
  always @ (posedge reset or posedge clock) if (reset) r577 <= 1'd0; else if (_12300) r577 <= _25540;
  wire [1:0] _25541 = {_0, _958} + {_0, _2813};
  wire [1:0] _25542 = {_0, _5694} + {_0, _8028};
  wire [2:0] _25543 = {_0, _25541} + {_0, _25542};
  wire [1:0] _25544 = {_0, _9469} + {_0, _11358};
  wire [3:0] _25545 = {_0, _25543} + {_0, _0, _25544};
  wire _25546 = _12301 < _25545;
  wire _25547 = r576 ^ _25546;
  wire _25548 = _12298 ? coded_block[576] : r576;
  wire _25549 = _12296 ? _25547 : _25548;
  always @ (posedge reset or posedge clock) if (reset) r576 <= 1'd0; else if (_12300) r576 <= _25549;
  wire [1:0] _25550 = {_0, _990} + {_0, _2878};
  wire [1:0] _25551 = {_0, _4895} + {_0, _7773};
  wire [2:0] _25552 = {_0, _25550} + {_0, _25551};
  wire [1:0] _25553 = {_0, _10108} + {_0, _11550};
  wire [3:0] _25554 = {_0, _25552} + {_0, _0, _25553};
  wire _25555 = _12301 < _25554;
  wire _25556 = r575 ^ _25555;
  wire _25557 = _12298 ? coded_block[575] : r575;
  wire _25558 = _12296 ? _25556 : _25557;
  always @ (posedge reset or posedge clock) if (reset) r575 <= 1'd0; else if (_12300) r575 <= _25558;
  wire [1:0] _25559 = {_0, _1021} + {_0, _3678};
  wire [1:0] _25560 = {_0, _4958} + {_0, _6973};
  wire [2:0] _25561 = {_0, _25559} + {_0, _25560};
  wire [1:0] _25562 = {_0, _9853} + {_0, _12188};
  wire [3:0] _25563 = {_0, _25561} + {_0, _0, _25562};
  wire _25564 = _12301 < _25563;
  wire _25565 = r574 ^ _25564;
  wire _25566 = _12298 ? coded_block[574] : r574;
  wire _25567 = _12296 ? _25565 : _25566;
  always @ (posedge reset or posedge clock) if (reset) r574 <= 1'd0; else if (_12300) r574 <= _25567;
  wire [1:0] _25568 = {_0, _1057} + {_0, _2367};
  wire [1:0] _25569 = {_0, _5757} + {_0, _7036};
  wire [2:0] _25570 = {_0, _25568} + {_0, _25569};
  wire [1:0] _25571 = {_0, _9054} + {_0, _11933};
  wire [3:0] _25572 = {_0, _25570} + {_0, _0, _25571};
  wire _25573 = _12301 < _25572;
  wire _25574 = r573 ^ _25573;
  wire _25575 = _12298 ? coded_block[573] : r573;
  wire _25576 = _12296 ? _25574 : _25575;
  always @ (posedge reset or posedge clock) if (reset) r573 <= 1'd0; else if (_12300) r573 <= _25576;
  wire [1:0] _25577 = {_0, _1088} + {_0, _2271};
  wire [1:0] _25578 = {_0, _4447} + {_0, _7837};
  wire [2:0] _25579 = {_0, _25577} + {_0, _25578};
  wire [1:0] _25580 = {_0, _9118} + {_0, _11132};
  wire [3:0] _25581 = {_0, _25579} + {_0, _0, _25580};
  wire _25582 = _12301 < _25581;
  wire _25583 = r572 ^ _25582;
  wire _25584 = _12298 ? coded_block[572] : r572;
  wire _25585 = _12296 ? _25583 : _25584;
  always @ (posedge reset or posedge clock) if (reset) r572 <= 1'd0; else if (_12300) r572 <= _25585;
  wire [1:0] _25586 = {_0, _1120} + {_0, _2782};
  wire [1:0] _25587 = {_0, _4350} + {_0, _6525};
  wire [2:0] _25588 = {_0, _25586} + {_0, _25587};
  wire [1:0] _25589 = {_0, _9917} + {_0, _11196};
  wire [3:0] _25590 = {_0, _25588} + {_0, _0, _25589};
  wire _25591 = _12301 < _25590;
  wire _25592 = r571 ^ _25591;
  wire _25593 = _12298 ? coded_block[571] : r571;
  wire _25594 = _12296 ? _25592 : _25593;
  always @ (posedge reset or posedge clock) if (reset) r571 <= 1'd0; else if (_12300) r571 <= _25594;
  wire [1:0] _25595 = {_0, _1151} + {_0, _3646};
  wire [1:0] _25596 = {_0, _4861} + {_0, _6431};
  wire [2:0] _25597 = {_0, _25595} + {_0, _25596};
  wire [1:0] _25598 = {_0, _8607} + {_0, _11996};
  wire [3:0] _25599 = {_0, _25597} + {_0, _0, _25598};
  wire _25600 = _12301 < _25599;
  wire _25601 = r570 ^ _25600;
  wire _25602 = _12298 ? coded_block[570] : r570;
  wire _25603 = _12296 ? _25601 : _25602;
  always @ (posedge reset or posedge clock) if (reset) r570 <= 1'd0; else if (_12300) r570 <= _25603;
  wire [1:0] _25604 = {_0, _1215} + {_0, _3964};
  wire [1:0] _25605 = {_0, _4989} + {_0, _7804};
  wire [2:0] _25606 = {_0, _25604} + {_0, _25605};
  wire [1:0] _25607 = {_0, _9022} + {_0, _10590};
  wire [3:0] _25608 = {_0, _25606} + {_0, _0, _25607};
  wire _25609 = _12301 < _25608;
  wire _25610 = r569 ^ _25609;
  wire _25611 = _12298 ? coded_block[569] : r569;
  wire _25612 = _12296 ? _25610 : _25611;
  always @ (posedge reset or posedge clock) if (reset) r569 <= 1'd0; else if (_12300) r569 <= _25612;
  wire [1:0] _25613 = {_0, _1247} + {_0, _2494};
  wire [1:0] _25614 = {_0, _6045} + {_0, _7069};
  wire [2:0] _25615 = {_0, _25613} + {_0, _25614};
  wire [1:0] _25616 = {_0, _9886} + {_0, _11101};
  wire [3:0] _25617 = {_0, _25615} + {_0, _0, _25616};
  wire _25618 = _12301 < _25617;
  wire _25619 = r568 ^ _25618;
  wire _25620 = _12298 ? coded_block[568] : r568;
  wire _25621 = _12296 ? _25619 : _25620;
  always @ (posedge reset or posedge clock) if (reset) r568 <= 1'd0; else if (_12300) r568 <= _25621;
  wire [1:0] _25622 = {_0, _1278} + {_0, _3580};
  wire [1:0] _25623 = {_0, _4574} + {_0, _8123};
  wire [2:0] _25624 = {_0, _25622} + {_0, _25623};
  wire [1:0] _25625 = {_0, _9149} + {_0, _11964};
  wire [3:0] _25626 = {_0, _25624} + {_0, _0, _25625};
  wire _25627 = _12301 < _25626;
  wire _25628 = r567 ^ _25627;
  wire _25629 = _12298 ? coded_block[567] : r567;
  wire _25630 = _12296 ? _25628 : _25629;
  always @ (posedge reset or posedge clock) if (reset) r567 <= 1'd0; else if (_12300) r567 <= _25630;
  wire [1:0] _25631 = {_0, _1312} + {_0, _3901};
  wire [1:0] _25632 = {_0, _5663} + {_0, _6652};
  wire [2:0] _25633 = {_0, _25631} + {_0, _25632};
  wire [1:0] _25634 = {_0, _10204} + {_0, _11228};
  wire [3:0] _25635 = {_0, _25633} + {_0, _0, _25634};
  wire _25636 = _12301 < _25635;
  wire _25637 = r566 ^ _25636;
  wire _25638 = _12298 ? coded_block[566] : r566;
  wire _25639 = _12296 ? _25637 : _25638;
  always @ (posedge reset or posedge clock) if (reset) r566 <= 1'd0; else if (_12300) r566 <= _25639;
  wire [1:0] _25640 = {_0, _1343} + {_0, _2336};
  wire [1:0] _25641 = {_0, _5981} + {_0, _7741};
  wire [2:0] _25642 = {_0, _25640} + {_0, _25641};
  wire [1:0] _25643 = {_0, _8736} + {_0, _12282};
  wire [3:0] _25644 = {_0, _25642} + {_0, _0, _25643};
  wire _25645 = _12301 < _25644;
  wire _25646 = r565 ^ _25645;
  wire _25647 = _12298 ? coded_block[565] : r565;
  wire _25648 = _12296 ? _25646 : _25647;
  always @ (posedge reset or posedge clock) if (reset) r565 <= 1'd0; else if (_12300) r565 <= _25648;
  wire [1:0] _25649 = {_0, _1375} + {_0, _3709};
  wire [1:0] _25650 = {_0, _4415} + {_0, _8059};
  wire [2:0] _25651 = {_0, _25649} + {_0, _25650};
  wire [1:0] _25652 = {_0, _9822} + {_0, _10814};
  wire [3:0] _25653 = {_0, _25651} + {_0, _0, _25652};
  wire _25654 = _12301 < _25653;
  wire _25655 = r564 ^ _25654;
  wire _25656 = _12298 ? coded_block[564] : r564;
  wire _25657 = _12296 ? _25655 : _25656;
  always @ (posedge reset or posedge clock) if (reset) r564 <= 1'd0; else if (_12300) r564 <= _25657;
  wire [1:0] _25658 = {_0, _1406} + {_0, _2623};
  wire [1:0] _25659 = {_0, _5790} + {_0, _6494};
  wire [2:0] _25660 = {_0, _25658} + {_0, _25659};
  wire [1:0] _25661 = {_0, _10141} + {_0, _11900};
  wire [3:0] _25662 = {_0, _25660} + {_0, _0, _25661};
  wire _25663 = _12301 < _25662;
  wire _25664 = r563 ^ _25663;
  wire _25665 = _12298 ? coded_block[563] : r563;
  wire _25666 = _12296 ? _25664 : _25665;
  always @ (posedge reset or posedge clock) if (reset) r563 <= 1'd0; else if (_12300) r563 <= _25666;
  wire [1:0] _25667 = {_0, _1439} + {_0, _2719};
  wire [1:0] _25668 = {_0, _4703} + {_0, _7868};
  wire [2:0] _25669 = {_0, _25667} + {_0, _25668};
  wire [1:0] _25670 = {_0, _8574} + {_0, _12219};
  wire [3:0] _25671 = {_0, _25669} + {_0, _0, _25670};
  wire _25672 = _12301 < _25671;
  wire _25673 = r562 ^ _25672;
  wire _25674 = _12298 ? coded_block[562] : r562;
  wire _25675 = _12296 ? _25673 : _25674;
  always @ (posedge reset or posedge clock) if (reset) r562 <= 1'd0; else if (_12300) r562 <= _25675;
  wire [1:0] _25676 = {_0, _1470} + {_0, _2175};
  wire [1:0] _25677 = {_0, _4798} + {_0, _6781};
  wire [2:0] _25678 = {_0, _25676} + {_0, _25677};
  wire [1:0] _25679 = {_0, _9949} + {_0, _10654};
  wire [3:0] _25680 = {_0, _25678} + {_0, _0, _25679};
  wire _25681 = _12301 < _25680;
  wire _25682 = r561 ^ _25681;
  wire _25683 = _12298 ? coded_block[561] : r561;
  wire _25684 = _12296 ? _25682 : _25683;
  always @ (posedge reset or posedge clock) if (reset) r561 <= 1'd0; else if (_12300) r561 <= _25684;
  wire [1:0] _25685 = {_0, _479} + {_0, _3104};
  wire [1:0] _25686 = {_0, _5884} + {_0, _6525};
  wire [2:0] _25687 = {_0, _25685} + {_0, _25686};
  wire [1:0] _25688 = {_0, _10141} + {_0, _11806};
  wire [3:0] _25689 = {_0, _25687} + {_0, _0, _25688};
  wire _25690 = _12301 < _25689;
  wire _25691 = r560 ^ _25690;
  wire _25692 = _12298 ? coded_block[560] : r560;
  wire _25693 = _12296 ? _25691 : _25692;
  always @ (posedge reset or posedge clock) if (reset) r560 <= 1'd0; else if (_12300) r560 <= _25693;
  wire [1:0] _25694 = {_0, _510} + {_0, _2782};
  wire [1:0] _25695 = {_0, _5183} + {_0, _7965};
  wire [2:0] _25696 = {_0, _25694} + {_0, _25695};
  wire [1:0] _25697 = {_0, _8607} + {_0, _12219};
  wire [3:0] _25698 = {_0, _25696} + {_0, _0, _25697};
  wire _25699 = _12301 < _25698;
  wire _25700 = r559 ^ _25699;
  wire _25701 = _12298 ? coded_block[559] : r559;
  wire _25702 = _12296 ? _25700 : _25701;
  always @ (posedge reset or posedge clock) if (reset) r559 <= 1'd0; else if (_12300) r559 <= _25702;
  wire [1:0] _25703 = {_0, _576} + {_0, _2750};
  wire [1:0] _25704 = {_0, _5022} + {_0, _6942};
  wire [2:0] _25705 = {_0, _25703} + {_0, _25704};
  wire [1:0] _25706 = {_0, _9342} + {_0, _12124};
  wire [3:0] _25707 = {_0, _25705} + {_0, _0, _25706};
  wire _25708 = _12301 < _25707;
  wire _25709 = r558 ^ _25708;
  wire _25710 = _12298 ? coded_block[558] : r558;
  wire _25711 = _12296 ? _25709 : _25710;
  always @ (posedge reset or posedge clock) if (reset) r558 <= 1'd0; else if (_12300) r558 <= _25711;
  wire [1:0] _25712 = {_0, _608} + {_0, _3135};
  wire [1:0] _25713 = {_0, _4830} + {_0, _7100};
  wire [2:0] _25714 = {_0, _25712} + {_0, _25713};
  wire [1:0] _25715 = {_0, _9022} + {_0, _11422};
  wire [3:0] _25716 = {_0, _25714} + {_0, _0, _25715};
  wire _25717 = _12301 < _25716;
  wire _25718 = r557 ^ _25717;
  wire _25719 = _12298 ? coded_block[557] : r557;
  wire _25720 = _12296 ? _25718 : _25719;
  always @ (posedge reset or posedge clock) if (reset) r557 <= 1'd0; else if (_12300) r557 <= _25720;
  wire [1:0] _25721 = {_0, _639} + {_0, _2271};
  wire [1:0] _25722 = {_0, _5215} + {_0, _6908};
  wire [2:0] _25723 = {_0, _25721} + {_0, _25722};
  wire [1:0] _25724 = {_0, _9181} + {_0, _11101};
  wire [3:0] _25725 = {_0, _25723} + {_0, _0, _25724};
  wire _25726 = _12301 < _25725;
  wire _25727 = r556 ^ _25726;
  wire _25728 = _12298 ? coded_block[556] : r556;
  wire _25729 = _12296 ? _25727 : _25728;
  always @ (posedge reset or posedge clock) if (reset) r556 <= 1'd0; else if (_12300) r556 <= _25729;
  wire [1:0] _25730 = {_0, _672} + {_0, _4060};
  wire [1:0] _25731 = {_0, _4350} + {_0, _7293};
  wire [2:0] _25732 = {_0, _25730} + {_0, _25731};
  wire [1:0] _25733 = {_0, _8991} + {_0, _11259};
  wire [3:0] _25734 = {_0, _25732} + {_0, _0, _25733};
  wire _25735 = _12301 < _25734;
  wire _25736 = r555 ^ _25735;
  wire _25737 = _12298 ? coded_block[555] : r555;
  wire _25738 = _12296 ? _25736 : _25737;
  always @ (posedge reset or posedge clock) if (reset) r555 <= 1'd0; else if (_12300) r555 <= _25738;
  wire [1:0] _25739 = {_0, _703} + {_0, _2623};
  wire [1:0] _25740 = {_0, _6139} + {_0, _6431};
  wire [2:0] _25741 = {_0, _25739} + {_0, _25740};
  wire [1:0] _25742 = {_0, _9375} + {_0, _11069};
  wire [3:0] _25743 = {_0, _25741} + {_0, _0, _25742};
  wire _25744 = _12301 < _25743;
  wire _25745 = r554 ^ _25744;
  wire _25746 = _12298 ? coded_block[554] : r554;
  wire _25747 = _12296 ? _25745 : _25746;
  always @ (posedge reset or posedge clock) if (reset) r554 <= 1'd0; else if (_12300) r554 <= _25747;
  wire [1:0] _25748 = {_0, _766} + {_0, _3678};
  wire [1:0] _25749 = {_0, _4640} + {_0, _6781};
  wire [2:0] _25750 = {_0, _25748} + {_0, _25749};
  wire [1:0] _25751 = {_0, _8288} + {_0, _10590};
  wire [3:0] _25752 = {_0, _25750} + {_0, _0, _25751};
  wire _25753 = _12301 < _25752;
  wire _25754 = r553 ^ _25753;
  wire _25755 = _12298 ? coded_block[553] : r553;
  wire _25756 = _12296 ? _25754 : _25755;
  always @ (posedge reset or posedge clock) if (reset) r553 <= 1'd0; else if (_12300) r553 <= _25756;
  wire [1:0] _25757 = {_0, _800} + {_0, _2336};
  wire [1:0] _25758 = {_0, _5757} + {_0, _6718};
  wire [2:0] _25759 = {_0, _25757} + {_0, _25758};
  wire [1:0] _25760 = {_0, _8863} + {_0, _10366};
  wire [3:0] _25761 = {_0, _25759} + {_0, _0, _25760};
  wire _25762 = _12301 < _25761;
  wire _25763 = r552 ^ _25762;
  wire _25764 = _12298 ? coded_block[552] : r552;
  wire _25765 = _12296 ? _25763 : _25764;
  always @ (posedge reset or posedge clock) if (reset) r552 <= 1'd0; else if (_12300) r552 <= _25765;
  wire [1:0] _25766 = {_0, _831} + {_0, _3933};
  wire [1:0] _25767 = {_0, _4415} + {_0, _7837};
  wire [2:0] _25768 = {_0, _25766} + {_0, _25767};
  wire [1:0] _25769 = {_0, _8799} + {_0, _10941};
  wire [3:0] _25770 = {_0, _25768} + {_0, _0, _25769};
  wire _25771 = _12301 < _25770;
  wire _25772 = r551 ^ _25771;
  wire _25773 = _12298 ? coded_block[551] : r551;
  wire _25774 = _12296 ? _25772 : _25773;
  always @ (posedge reset or posedge clock) if (reset) r551 <= 1'd0; else if (_12300) r551 <= _25774;
  wire [1:0] _25775 = {_0, _863} + {_0, _3646};
  wire [1:0] _25776 = {_0, _6012} + {_0, _6494};
  wire [2:0] _25777 = {_0, _25775} + {_0, _25776};
  wire [1:0] _25778 = {_0, _9917} + {_0, _10877};
  wire [3:0] _25779 = {_0, _25777} + {_0, _0, _25778};
  wire _25780 = _12301 < _25779;
  wire _25781 = r550 ^ _25780;
  wire _25782 = _12298 ? coded_block[550] : r550;
  wire _25783 = _12296 ? _25781 : _25782;
  always @ (posedge reset or posedge clock) if (reset) r550 <= 1'd0; else if (_12300) r550 <= _25783;
  wire [1:0] _25784 = {_0, _894} + {_0, _2592};
  wire [1:0] _25785 = {_0, _5726} + {_0, _8092};
  wire [2:0] _25786 = {_0, _25784} + {_0, _25785};
  wire [1:0] _25787 = {_0, _8574} + {_0, _11996};
  wire [3:0] _25788 = {_0, _25786} + {_0, _0, _25787};
  wire _25789 = _12301 < _25788;
  wire _25790 = r549 ^ _25789;
  wire _25791 = _12298 ? coded_block[549] : r549;
  wire _25792 = _12296 ? _25790 : _25791;
  always @ (posedge reset or posedge clock) if (reset) r549 <= 1'd0; else if (_12300) r549 <= _25792;
  wire [1:0] _25793 = {_0, _927} + {_0, _4091};
  wire [1:0] _25794 = {_0, _4671} + {_0, _7804};
  wire [2:0] _25795 = {_0, _25793} + {_0, _25794};
  wire [1:0] _25796 = {_0, _10172} + {_0, _10654};
  wire [3:0] _25797 = {_0, _25795} + {_0, _0, _25796};
  wire _25798 = _12301 < _25797;
  wire _25799 = r548 ^ _25798;
  wire _25800 = _12298 ? coded_block[548] : r548;
  wire _25801 = _12296 ? _25799 : _25800;
  always @ (posedge reset or posedge clock) if (reset) r548 <= 1'd0; else if (_12300) r548 <= _25801;
  wire [1:0] _25802 = {_0, _958} + {_0, _3068};
  wire [1:0] _25803 = {_0, _4160} + {_0, _6750};
  wire [2:0] _25804 = {_0, _25802} + {_0, _25803};
  wire [1:0] _25805 = {_0, _9886} + {_0, _12251};
  wire [3:0] _25806 = {_0, _25804} + {_0, _0, _25805};
  wire _25807 = _12301 < _25806;
  wire _25808 = r547 ^ _25807;
  wire _25809 = _12298 ? coded_block[547] : r547;
  wire _25810 = _12296 ? _25808 : _25809;
  always @ (posedge reset or posedge clock) if (reset) r547 <= 1'd0; else if (_12300) r547 <= _25810;
  wire [1:0] _25811 = {_0, _990} + {_0, _3836};
  wire [1:0] _25812 = {_0, _5152} + {_0, _6239};
  wire [2:0] _25813 = {_0, _25811} + {_0, _25812};
  wire [1:0] _25814 = {_0, _8830} + {_0, _11964};
  wire [3:0] _25815 = {_0, _25813} + {_0, _0, _25814};
  wire _25816 = _12301 < _25815;
  wire _25817 = r546 ^ _25816;
  wire _25818 = _12298 ? coded_block[546] : r546;
  wire _25819 = _12296 ? _25817 : _25818;
  always @ (posedge reset or posedge clock) if (reset) r546 <= 1'd0; else if (_12300) r546 <= _25819;
  wire [1:0] _25820 = {_0, _1021} + {_0, _3005};
  wire [1:0] _25821 = {_0, _5918} + {_0, _7230};
  wire [2:0] _25822 = {_0, _25820} + {_0, _25821};
  wire [1:0] _25823 = {_0, _8319} + {_0, _10910};
  wire [3:0] _25824 = {_0, _25822} + {_0, _0, _25823};
  wire _25825 = _12301 < _25824;
  wire _25826 = r545 ^ _25825;
  wire _25827 = _12298 ? coded_block[545] : r545;
  wire _25828 = _12296 ? _25826 : _25827;
  always @ (posedge reset or posedge clock) if (reset) r545 <= 1'd0; else if (_12300) r545 <= _25828;
  wire [1:0] _25829 = {_0, _1057} + {_0, _2526};
  wire [1:0] _25830 = {_0, _5085} + {_0, _7996};
  wire [2:0] _25831 = {_0, _25829} + {_0, _25830};
  wire [1:0] _25832 = {_0, _9311} + {_0, _10399};
  wire [3:0] _25833 = {_0, _25831} + {_0, _0, _25832};
  wire _25834 = _12301 < _25833;
  wire _25835 = r544 ^ _25834;
  wire _25836 = _12298 ? coded_block[544] : r544;
  wire _25837 = _12296 ? _25835 : _25836;
  always @ (posedge reset or posedge clock) if (reset) r544 <= 1'd0; else if (_12300) r544 <= _25837;
  wire [1:0] _25838 = {_0, _1088} + {_0, _2655};
  wire [1:0] _25839 = {_0, _4605} + {_0, _7163};
  wire [2:0] _25840 = {_0, _25838} + {_0, _25839};
  wire [1:0] _25841 = {_0, _10077} + {_0, _11389};
  wire [3:0] _25842 = {_0, _25840} + {_0, _0, _25841};
  wire _25843 = _12301 < _25842;
  wire _25844 = r543 ^ _25843;
  wire _25845 = _12298 ? coded_block[543] : r543;
  wire _25846 = _12296 ? _25844 : _25845;
  always @ (posedge reset or posedge clock) if (reset) r543 <= 1'd0; else if (_12300) r543 <= _25846;
  wire [1:0] _25847 = {_0, _1120} + {_0, _3997};
  wire [1:0] _25848 = {_0, _4734} + {_0, _6687};
  wire [2:0] _25849 = {_0, _25847} + {_0, _25848};
  wire [1:0] _25850 = {_0, _9248} + {_0, _12155};
  wire [3:0] _25851 = {_0, _25849} + {_0, _0, _25850};
  wire _25852 = _12301 < _25851;
  wire _25853 = r542 ^ _25852;
  wire _25854 = _12298 ? coded_block[542] : r542;
  wire _25855 = _12296 ? _25853 : _25854;
  always @ (posedge reset or posedge clock) if (reset) r542 <= 1'd0; else if (_12300) r542 <= _25855;
  wire [1:0] _25856 = {_0, _1151} + {_0, _3231};
  wire [1:0] _25857 = {_0, _6076} + {_0, _6814};
  wire [2:0] _25858 = {_0, _25856} + {_0, _25857};
  wire [1:0] _25859 = {_0, _8767} + {_0, _11326};
  wire [3:0] _25860 = {_0, _25858} + {_0, _0, _25859};
  wire _25861 = _12301 < _25860;
  wire _25862 = r541 ^ _25861;
  wire _25863 = _12298 ? coded_block[541] : r541;
  wire _25864 = _12296 ? _25862 : _25863;
  always @ (posedge reset or posedge clock) if (reset) r541 <= 1'd0; else if (_12300) r541 <= _25864;
  wire [1:0] _25865 = {_0, _1184} + {_0, _3198};
  wire [1:0] _25866 = {_0, _5310} + {_0, _8155};
  wire [2:0] _25867 = {_0, _25865} + {_0, _25866};
  wire [1:0] _25868 = {_0, _8894} + {_0, _10846};
  wire [3:0] _25869 = {_0, _25867} + {_0, _0, _25868};
  wire _25870 = _12301 < _25869;
  wire _25871 = r540 ^ _25870;
  wire _25872 = _12298 ? coded_block[540] : r540;
  wire _25873 = _12296 ? _25871 : _25872;
  always @ (posedge reset or posedge clock) if (reset) r540 <= 1'd0; else if (_12300) r540 <= _25873;
  wire [1:0] _25874 = {_0, _1215} + {_0, _4028};
  wire [1:0] _25875 = {_0, _5279} + {_0, _7389};
  wire [2:0] _25876 = {_0, _25874} + {_0, _25875};
  wire [1:0] _25877 = {_0, _10235} + {_0, _10973};
  wire [3:0] _25878 = {_0, _25876} + {_0, _0, _25877};
  wire _25879 = _12301 < _25878;
  wire _25880 = r539 ^ _25879;
  wire _25881 = _12298 ? coded_block[539] : r539;
  wire _25882 = _12296 ? _25880 : _25881;
  always @ (posedge reset or posedge clock) if (reset) r539 <= 1'd0; else if (_12300) r539 <= _25882;
  wire [1:0] _25883 = {_0, _1247} + {_0, _2302};
  wire [1:0] _25884 = {_0, _6108} + {_0, _7357};
  wire [2:0] _25885 = {_0, _25883} + {_0, _25884};
  wire [1:0] _25886 = {_0, _9469} + {_0, _10303};
  wire [3:0] _25887 = {_0, _25885} + {_0, _0, _25886};
  wire _25888 = _12301 < _25887;
  wire _25889 = r538 ^ _25888;
  wire _25890 = _12298 ? coded_block[538] : r538;
  wire _25891 = _12296 ? _25889 : _25890;
  always @ (posedge reset or posedge clock) if (reset) r538 <= 1'd0; else if (_12300) r538 <= _25891;
  wire [1:0] _25892 = {_0, _1278} + {_0, _3709};
  wire [1:0] _25893 = {_0, _4384} + {_0, _8186};
  wire [2:0] _25894 = {_0, _25892} + {_0, _25893};
  wire [1:0] _25895 = {_0, _9438} + {_0, _11550};
  wire [3:0] _25896 = {_0, _25894} + {_0, _0, _25895};
  wire _25897 = _12301 < _25896;
  wire _25898 = r537 ^ _25897;
  wire _25899 = _12298 ? coded_block[537] : r537;
  wire _25900 = _12296 ? _25898 : _25899;
  always @ (posedge reset or posedge clock) if (reset) r537 <= 1'd0; else if (_12300) r537 <= _25900;
  wire [1:0] _25901 = {_0, _1312} + {_0, _3549};
  wire [1:0] _25902 = {_0, _5790} + {_0, _6462};
  wire [2:0] _25903 = {_0, _25901} + {_0, _25902};
  wire [1:0] _25904 = {_0, _8256} + {_0, _11516};
  wire [3:0] _25905 = {_0, _25903} + {_0, _0, _25904};
  wire _25906 = _12301 < _25905;
  wire _25907 = r536 ^ _25906;
  wire _25908 = _12298 ? coded_block[536] : r536;
  wire _25909 = _12296 ? _25907 : _25908;
  always @ (posedge reset or posedge clock) if (reset) r536 <= 1'd0; else if (_12300) r536 <= _25909;
  wire [1:0] _25910 = {_0, _1343} + {_0, _2081};
  wire [1:0] _25911 = {_0, _5628} + {_0, _7868};
  wire [2:0] _25912 = {_0, _25910} + {_0, _25911};
  wire [1:0] _25913 = {_0, _8543} + {_0, _10335};
  wire [3:0] _25914 = {_0, _25912} + {_0, _0, _25913};
  wire _25915 = _12301 < _25914;
  wire _25916 = r535 ^ _25915;
  wire _25917 = _12298 ? coded_block[535] : r535;
  wire _25918 = _12296 ? _25916 : _25917;
  always @ (posedge reset or posedge clock) if (reset) r535 <= 1'd0; else if (_12300) r535 <= _25918;
  wire [1:0] _25919 = {_0, _1375} + {_0, _3580};
  wire [1:0] _25920 = {_0, _4129} + {_0, _7710};
  wire [2:0] _25921 = {_0, _25919} + {_0, _25920};
  wire [1:0] _25922 = {_0, _9949} + {_0, _10621};
  wire [3:0] _25923 = {_0, _25921} + {_0, _0, _25922};
  wire _25924 = _12301 < _25923;
  wire _25925 = r534 ^ _25924;
  wire _25926 = _12298 ? coded_block[534] : r534;
  wire _25927 = _12296 ? _25925 : _25926;
  always @ (posedge reset or posedge clock) if (reset) r534 <= 1'd0; else if (_12300) r534 <= _25927;
  wire [1:0] _25928 = {_0, _1406} + {_0, _3773};
  wire [1:0] _25929 = {_0, _5663} + {_0, _6176};
  wire [2:0] _25930 = {_0, _25928} + {_0, _25929};
  wire [1:0] _25931 = {_0, _9790} + {_0, _12027};
  wire [3:0] _25932 = {_0, _25930} + {_0, _0, _25931};
  wire _25933 = _12301 < _25932;
  wire _25934 = r533 ^ _25933;
  wire _25935 = _12298 ? coded_block[533] : r533;
  wire _25936 = _12296 ? _25934 : _25935;
  always @ (posedge reset or posedge clock) if (reset) r533 <= 1'd0; else if (_12300) r533 <= _25936;
  wire [1:0] _25937 = {_0, _1439} + {_0, _2399};
  wire [1:0] _25938 = {_0, _5853} + {_0, _7741};
  wire [2:0] _25939 = {_0, _25937} + {_0, _25938};
  wire [1:0] _25940 = {_0, _8225} + {_0, _11869};
  wire [3:0] _25941 = {_0, _25939} + {_0, _0, _25940};
  wire _25942 = _12301 < _25941;
  wire _25943 = r532 ^ _25942;
  wire _25944 = _12298 ? coded_block[532] : r532;
  wire _25945 = _12296 ? _25943 : _25944;
  always @ (posedge reset or posedge clock) if (reset) r532 <= 1'd0; else if (_12300) r532 <= _25945;
  wire [1:0] _25946 = {_0, _1470} + {_0, _2144};
  wire [1:0] _25947 = {_0, _4478} + {_0, _7931};
  wire [2:0] _25948 = {_0, _25946} + {_0, _25947};
  wire [1:0] _25949 = {_0, _9822} + {_0, _10272};
  wire [3:0] _25950 = {_0, _25948} + {_0, _0, _25949};
  wire _25951 = _12301 < _25950;
  wire _25952 = r531 ^ _25951;
  wire _25953 = _12298 ? coded_block[531] : r531;
  wire _25954 = _12296 ? _25952 : _25953;
  always @ (posedge reset or posedge clock) if (reset) r531 <= 1'd0; else if (_12300) r531 <= _25954;
  wire [1:0] _25955 = {_0, _1502} + {_0, _3359};
  wire [1:0] _25956 = {_0, _4223} + {_0, _6558};
  wire [2:0] _25957 = {_0, _25955} + {_0, _25956};
  wire [1:0] _25958 = {_0, _10014} + {_0, _11900};
  wire [3:0] _25959 = {_0, _25957} + {_0, _0, _25958};
  wire _25960 = _12301 < _25959;
  wire _25961 = r530 ^ _25960;
  wire _25962 = _12298 ? coded_block[530] : r530;
  wire _25963 = _12296 ? _25961 : _25962;
  always @ (posedge reset or posedge clock) if (reset) r530 <= 1'd0; else if (_12300) r530 <= _25963;
  wire [1:0] _25964 = {_0, _1533} + {_0, _3422};
  wire [1:0] _25965 = {_0, _5438} + {_0, _6303};
  wire [2:0] _25966 = {_0, _25964} + {_0, _25965};
  wire [1:0] _25967 = {_0, _8638} + {_0, _12092};
  wire [3:0] _25968 = {_0, _25966} + {_0, _0, _25967};
  wire _25969 = _12301 < _25968;
  wire _25970 = r529 ^ _25969;
  wire _25971 = _12298 ? coded_block[529] : r529;
  wire _25972 = _12296 ? _25970 : _25971;
  always @ (posedge reset or posedge clock) if (reset) r529 <= 1'd0; else if (_12300) r529 <= _25972;
  wire [1:0] _25973 = {_0, _1568} + {_0, _2208};
  wire [1:0] _25974 = {_0, _5501} + {_0, _7517};
  wire [2:0] _25975 = {_0, _25973} + {_0, _25974};
  wire [1:0] _25976 = {_0, _8383} + {_0, _10717};
  wire [3:0] _25977 = {_0, _25975} + {_0, _0, _25976};
  wire _25978 = _12301 < _25977;
  wire _25979 = r528 ^ _25978;
  wire _25980 = _12298 ? coded_block[528] : r528;
  wire _25981 = _12296 ? _25979 : _25980;
  always @ (posedge reset or posedge clock) if (reset) r528 <= 1'd0; else if (_12300) r528 <= _25981;
  wire [1:0] _25982 = {_0, _1599} + {_0, _2910};
  wire [1:0] _25983 = {_0, _4287} + {_0, _7581};
  wire [2:0] _25984 = {_0, _25982} + {_0, _25983};
  wire [1:0] _25985 = {_0, _9597} + {_0, _10462};
  wire [3:0] _25986 = {_0, _25984} + {_0, _0, _25985};
  wire _25987 = _12301 < _25986;
  wire _25988 = r527 ^ _25987;
  wire _25989 = _12298 ? coded_block[527] : r527;
  wire _25990 = _12296 ? _25988 : _25989;
  always @ (posedge reset or posedge clock) if (reset) r527 <= 1'd0; else if (_12300) r527 <= _25990;
  wire [1:0] _25991 = {_0, _1631} + {_0, _2813};
  wire [1:0] _25992 = {_0, _4989} + {_0, _6366};
  wire [2:0] _25993 = {_0, _25991} + {_0, _25992};
  wire [1:0] _25994 = {_0, _9661} + {_0, _11677};
  wire [3:0] _25995 = {_0, _25993} + {_0, _0, _25994};
  wire _25996 = _12301 < _25995;
  wire _25997 = r526 ^ _25996;
  wire _25998 = _12298 ? coded_block[526] : r526;
  wire _25999 = _12296 ? _25997 : _25998;
  always @ (posedge reset or posedge clock) if (reset) r526 <= 1'd0; else if (_12300) r526 <= _25999;
  wire [1:0] _26000 = {_0, _1662} + {_0, _3325};
  wire [1:0] _26001 = {_0, _4895} + {_0, _7069};
  wire [2:0] _26002 = {_0, _26000} + {_0, _26001};
  wire [1:0] _26003 = {_0, _8446} + {_0, _11740};
  wire [3:0] _26004 = {_0, _26002} + {_0, _0, _26003};
  wire _26005 = _12301 < _26004;
  wire _26006 = r525 ^ _26005;
  wire _26007 = _12298 ? coded_block[525] : r525;
  wire _26008 = _12296 ? _26006 : _26007;
  always @ (posedge reset or posedge clock) if (reset) r525 <= 1'd0; else if (_12300) r525 <= _26008;
  wire [1:0] _26009 = {_0, _1695} + {_0, _2175};
  wire [1:0] _26010 = {_0, _5407} + {_0, _6973};
  wire [2:0] _26011 = {_0, _26009} + {_0, _26010};
  wire [1:0] _26012 = {_0, _9149} + {_0, _10527};
  wire [3:0] _26013 = {_0, _26011} + {_0, _0, _26012};
  wire _26014 = _12301 < _26013;
  wire _26015 = r524 ^ _26014;
  wire _26016 = _12298 ? coded_block[524] : r524;
  wire _26017 = _12296 ? _26015 : _26016;
  always @ (posedge reset or posedge clock) if (reset) r524 <= 1'd0; else if (_12300) r524 <= _26017;
  wire [1:0] _26018 = {_0, _1758} + {_0, _2494};
  wire [1:0] _26019 = {_0, _5534} + {_0, _6334};
  wire [2:0] _26020 = {_0, _26018} + {_0, _26019};
  wire [1:0] _26021 = {_0, _9566} + {_0, _11132};
  wire [3:0] _26022 = {_0, _26020} + {_0, _0, _26021};
  wire _26023 = _12301 < _26022;
  wire _26024 = r523 ^ _26023;
  wire _26025 = _12298 ? coded_block[523] : r523;
  wire _26026 = _12296 ? _26024 : _26025;
  always @ (posedge reset or posedge clock) if (reset) r523 <= 1'd0; else if (_12300) r523 <= _26026;
  wire [1:0] _26027 = {_0, _1789} + {_0, _3037};
  wire [1:0] _26028 = {_0, _4574} + {_0, _7612};
  wire [2:0] _26029 = {_0, _26027} + {_0, _26028};
  wire [1:0] _26030 = {_0, _8415} + {_0, _11644};
  wire [3:0] _26031 = {_0, _26029} + {_0, _0, _26030};
  wire _26032 = _12301 < _26031;
  wire _26033 = r522 ^ _26032;
  wire _26034 = _12298 ? coded_block[522] : r522;
  wire _26035 = _12296 ? _26033 : _26034;
  always @ (posedge reset or posedge clock) if (reset) r522 <= 1'd0; else if (_12300) r522 <= _26035;
  wire [1:0] _26036 = {_0, _1823} + {_0, _2112};
  wire [1:0] _26037 = {_0, _5116} + {_0, _6652};
  wire [2:0] _26038 = {_0, _26036} + {_0, _26037};
  wire [1:0] _26039 = {_0, _9693} + {_0, _10493};
  wire [3:0] _26040 = {_0, _26038} + {_0, _0, _26039};
  wire _26041 = _12301 < _26040;
  wire _26042 = r521 ^ _26041;
  wire _26043 = _12298 ? coded_block[521] : r521;
  wire _26044 = _12296 ? _26042 : _26043;
  always @ (posedge reset or posedge clock) if (reset) r521 <= 1'd0; else if (_12300) r521 <= _26044;
  wire [1:0] _26045 = {_0, _1854} + {_0, _2430};
  wire [1:0] _26046 = {_0, _4192} + {_0, _7199};
  wire [2:0] _26047 = {_0, _26045} + {_0, _26046};
  wire [1:0] _26048 = {_0, _8736} + {_0, _11771};
  wire [3:0] _26049 = {_0, _26047} + {_0, _0, _26048};
  wire _26050 = _12301 < _26049;
  wire _26051 = r520 ^ _26050;
  wire _26052 = _12298 ? coded_block[520] : r520;
  wire _26053 = _12296 ? _26051 : _26052;
  always @ (posedge reset or posedge clock) if (reset) r520 <= 1'd0; else if (_12300) r520 <= _26053;
  wire [1:0] _26054 = {_0, _1886} + {_0, _2878};
  wire [1:0] _26055 = {_0, _4511} + {_0, _6270};
  wire [2:0] _26056 = {_0, _26054} + {_0, _26055};
  wire [1:0] _26057 = {_0, _9279} + {_0, _10814};
  wire [3:0] _26058 = {_0, _26056} + {_0, _0, _26057};
  wire _26059 = _12301 < _26058;
  wire _26060 = r519 ^ _26059;
  wire _26061 = _12298 ? coded_block[519] : r519;
  wire _26062 = _12296 ? _26060 : _26061;
  always @ (posedge reset or posedge clock) if (reset) r519 <= 1'd0; else if (_12300) r519 <= _26062;
  wire [1:0] _26063 = {_0, _1950} + {_0, _3167};
  wire [1:0] _26064 = {_0, _4319} + {_0, _7036};
  wire [2:0] _26065 = {_0, _26063} + {_0, _26064};
  wire [1:0] _26066 = {_0, _8670} + {_0, _10430};
  wire [3:0] _26067 = {_0, _26065} + {_0, _0, _26066};
  wire _26068 = _12301 < _26067;
  wire _26069 = r518 ^ _26068;
  wire _26070 = _12298 ? coded_block[518] : r518;
  wire _26071 = _12296 ? _26069 : _26070;
  always @ (posedge reset or posedge clock) if (reset) r518 <= 1'd0; else if (_12300) r518 <= _26071;
  wire [1:0] _26072 = {_0, _1981} + {_0, _3262};
  wire [1:0] _26073 = {_0, _5246} + {_0, _6397};
  wire [2:0] _26074 = {_0, _26072} + {_0, _26073};
  wire [1:0] _26075 = {_0, _9118} + {_0, _10748};
  wire [3:0] _26076 = {_0, _26074} + {_0, _0, _26075};
  wire _26077 = _12301 < _26076;
  wire _26078 = r517 ^ _26077;
  wire _26079 = _12298 ? coded_block[517] : r517;
  wire _26080 = _12296 ? _26078 : _26079;
  always @ (posedge reset or posedge clock) if (reset) r517 <= 1'd0; else if (_12300) r517 <= _26080;
  wire [1:0] _26081 = {_0, _2044} + {_0, _2974};
  wire [1:0] _26082 = {_0, _4798} + {_0, _7420};
  wire [2:0] _26083 = {_0, _26081} + {_0, _26082};
  wire [1:0] _26084 = {_0, _9406} + {_0, _10558};
  wire [3:0] _26085 = {_0, _26083} + {_0, _0, _26084};
  wire _26086 = _12301 < _26085;
  wire _26087 = r516 ^ _26086;
  wire _26088 = _12298 ? coded_block[516] : r516;
  wire _26089 = _12296 ? _26087 : _26088;
  always @ (posedge reset or posedge clock) if (reset) r516 <= 1'd0; else if (_12300) r516 <= _26089;
  wire [1:0] _26090 = {_0, _65} + {_0, _3870};
  wire [1:0] _26091 = {_0, _5053} + {_0, _6877};
  wire [2:0] _26092 = {_0, _26090} + {_0, _26091};
  wire [1:0] _26093 = {_0, _9503} + {_0, _11485};
  wire [3:0] _26094 = {_0, _26092} + {_0, _0, _26093};
  wire _26095 = _12301 < _26094;
  wire _26096 = r515 ^ _26095;
  wire _26097 = _12298 ? coded_block[515] : r515;
  wire _26098 = _12296 ? _26096 : _26097;
  always @ (posedge reset or posedge clock) if (reset) r515 <= 1'd0; else if (_12300) r515 <= _26098;
  wire [1:0] _26099 = {_0, _128} + {_0, _3742};
  wire [1:0] _26100 = {_0, _5597} + {_0, _8028};
  wire [2:0] _26101 = {_0, _26099} + {_0, _26100};
  wire [1:0] _26102 = {_0, _9212} + {_0, _11038};
  wire [3:0] _26103 = {_0, _26101} + {_0, _0, _26102};
  wire _26104 = _12301 < _26103;
  wire _26105 = r514 ^ _26104;
  wire _26106 = _12298 ? coded_block[514] : r514;
  wire _26107 = _12296 ? _26105 : _26106;
  always @ (posedge reset or posedge clock) if (reset) r514 <= 1'd0; else if (_12300) r514 <= _26107;
  wire [1:0] _26108 = {_0, _161} + {_0, _3615};
  wire [1:0] _26109 = {_0, _5821} + {_0, _7675};
  wire [2:0] _26110 = {_0, _26108} + {_0, _26109};
  wire [1:0] _26111 = {_0, _10108} + {_0, _11295};
  wire [3:0] _26112 = {_0, _26110} + {_0, _0, _26111};
  wire _26113 = _12301 < _26112;
  wire _26114 = r513 ^ _26113;
  wire _26115 = _12298 ? coded_block[513] : r513;
  wire _26116 = _12296 ? _26114 : _26115;
  always @ (posedge reset or posedge clock) if (reset) r513 <= 1'd0; else if (_12300) r513 <= _26116;
  wire [1:0] _26117 = {_0, _192} + {_0, _3964};
  wire [1:0] _26118 = {_0, _5694} + {_0, _7900};
  wire [2:0] _26119 = {_0, _26117} + {_0, _26118};
  wire [1:0] _26120 = {_0, _9759} + {_0, _12188};
  wire [3:0] _26121 = {_0, _26119} + {_0, _0, _26120};
  wire _26122 = _12301 < _26121;
  wire _26123 = r512 ^ _26122;
  wire _26124 = _12298 ? coded_block[512] : r512;
  wire _26125 = _12296 ? _26123 : _26124;
  always @ (posedge reset or posedge clock) if (reset) r512 <= 1'd0; else if (_12300) r512 <= _26125;
  wire [1:0] _26126 = {_0, _224} + {_0, _2686};
  wire [1:0] _26127 = {_0, _6045} + {_0, _7773};
  wire [2:0] _26128 = {_0, _26126} + {_0, _26127};
  wire [1:0] _26129 = {_0, _9980} + {_0, _11837};
  wire [3:0] _26130 = {_0, _26128} + {_0, _0, _26129};
  wire _26131 = _12301 < _26130;
  wire _26132 = r511 ^ _26131;
  wire _26133 = _12298 ? coded_block[511] : r511;
  wire _26134 = _12296 ? _26132 : _26133;
  always @ (posedge reset or posedge clock) if (reset) r511 <= 1'd0; else if (_12300) r511 <= _26134;
  wire [1:0] _26135 = {_0, _255} + {_0, _3294};
  wire [1:0] _26136 = {_0, _4767} + {_0, _8123};
  wire [2:0] _26137 = {_0, _26135} + {_0, _26136};
  wire [1:0] _26138 = {_0, _9853} + {_0, _12061};
  wire [3:0] _26139 = {_0, _26137} + {_0, _0, _26138};
  wire _26140 = _12301 < _26139;
  wire _26141 = r510 ^ _26140;
  wire _26142 = _12298 ? coded_block[510] : r510;
  wire _26143 = _12296 ? _26141 : _26142;
  always @ (posedge reset or posedge clock) if (reset) r510 <= 1'd0; else if (_12300) r510 <= _26143;
  wire [1:0] _26144 = {_0, _320} + {_0, _2463};
  wire [1:0] _26145 = {_0, _4926} + {_0, _7454};
  wire [2:0] _26146 = {_0, _26144} + {_0, _26145};
  wire [1:0] _26147 = {_0, _8926} + {_0, _12282};
  wire [3:0] _26148 = {_0, _26146} + {_0, _0, _26147};
  wire _26149 = _12301 < _26148;
  wire _26150 = r509 ^ _26149;
  wire _26151 = _12298 ? coded_block[509] : r509;
  wire _26152 = _12296 ? _26150 : _26151;
  always @ (posedge reset or posedge clock) if (reset) r509 <= 1'd0; else if (_12300) r509 <= _26152;
  wire [1:0] _26153 = {_0, _352} + {_0, _3486};
  wire [1:0] _26154 = {_0, _4542} + {_0, _7005};
  wire [2:0] _26155 = {_0, _26153} + {_0, _26154};
  wire [1:0] _26156 = {_0, _9534} + {_0, _11004};
  wire [3:0] _26157 = {_0, _26155} + {_0, _0, _26156};
  wire _26158 = _12301 < _26157;
  wire _26159 = r508 ^ _26158;
  wire _26160 = _12298 ? coded_block[508] : r508;
  wire _26161 = _12296 ? _26159 : _26160;
  always @ (posedge reset or posedge clock) if (reset) r508 <= 1'd0; else if (_12300) r508 <= _26161;
  wire [1:0] _26162 = {_0, _416} + {_0, _2367};
  wire [1:0] _26163 = {_0, _5981} + {_0, _7644};
  wire [2:0] _26164 = {_0, _26162} + {_0, _26163};
  wire [1:0] _26165 = {_0, _8701} + {_0, _11165};
  wire [3:0] _26166 = {_0, _26164} + {_0, _0, _26165};
  wire _26167 = _12301 < _26166;
  wire _26168 = r507 ^ _26167;
  wire _26169 = _12298 ? coded_block[507] : r507;
  wire _26170 = _12296 ? _26168 : _26169;
  always @ (posedge reset or posedge clock) if (reset) r507 <= 1'd0; else if (_12300) r507 <= _26170;
  wire [1:0] _26171 = {_0, _447} + {_0, _3805};
  wire [1:0] _26172 = {_0, _4447} + {_0, _8059};
  wire [2:0] _26173 = {_0, _26171} + {_0, _26172};
  wire [1:0] _26174 = {_0, _9724} + {_0, _10783};
  wire [3:0] _26175 = {_0, _26173} + {_0, _0, _26174};
  wire _26176 = _12301 < _26175;
  wire _26177 = r506 ^ _26176;
  wire _26178 = _12298 ? coded_block[506] : r506;
  wire _26179 = _12296 ? _26177 : _26178;
  always @ (posedge reset or posedge clock) if (reset) r506 <= 1'd0; else if (_12300) r506 <= _26179;
  wire [1:0] _26180 = {_0, _34} + {_0, _2750};
  wire [1:0] _26181 = {_0, _4830} + {_0, _6908};
  wire [2:0] _26182 = {_0, _26180} + {_0, _26181};
  wire [1:0] _26183 = {_0, _8991} + {_0, _11069};
  wire [3:0] _26184 = {_0, _26182} + {_0, _0, _26183};
  wire _26185 = _12301 < _26184;
  wire _26186 = r505 ^ _26185;
  wire _26187 = _12298 ? coded_block[505] : r505;
  wire _26188 = _12296 ? _26186 : _26187;
  always @ (posedge reset or posedge clock) if (reset) r505 <= 1'd0; else if (_12300) r505 <= _26188;
  wire [1:0] _26189 = {_0, _1057} + {_0, _3549};
  wire [1:0] _26190 = {_0, _4767} + {_0, _6334};
  wire [2:0] _26191 = {_0, _26189} + {_0, _26190};
  wire [1:0] _26192 = {_0, _8511} + {_0, _11900};
  wire [3:0] _26193 = {_0, _26191} + {_0, _0, _26192};
  wire _26194 = _12301 < _26193;
  wire _26195 = r504 ^ _26194;
  wire _26196 = _12298 ? coded_block[504] : r504;
  wire _26197 = _12296 ? _26195 : _26196;
  always @ (posedge reset or posedge clock) if (reset) r504 <= 1'd0; else if (_12300) r504 <= _26197;
  wire [1:0] _26198 = {_0, _1088} + {_0, _2813};
  wire [1:0] _26199 = {_0, _5628} + {_0, _6845};
  wire [2:0] _26200 = {_0, _26198} + {_0, _26199};
  wire [1:0] _26201 = {_0, _8415} + {_0, _10590};
  wire [3:0] _26202 = {_0, _26200} + {_0, _0, _26201};
  wire _26203 = _12301 < _26202;
  wire _26204 = r503 ^ _26203;
  wire _26205 = _12298 ? coded_block[503] : r503;
  wire _26206 = _12296 ? _26204 : _26205;
  always @ (posedge reset or posedge clock) if (reset) r503 <= 1'd0; else if (_12300) r503 <= _26206;
  wire [1:0] _26207 = {_0, _1120} + {_0, _3870};
  wire [1:0] _26208 = {_0, _4895} + {_0, _7710};
  wire [2:0] _26209 = {_0, _26207} + {_0, _26208};
  wire [1:0] _26210 = {_0, _8926} + {_0, _10493};
  wire [3:0] _26211 = {_0, _26209} + {_0, _0, _26210};
  wire _26212 = _12301 < _26211;
  wire _26213 = r502 ^ _26212;
  wire _26214 = _12298 ? coded_block[502] : r502;
  wire _26215 = _12296 ? _26213 : _26214;
  always @ (posedge reset or posedge clock) if (reset) r502 <= 1'd0; else if (_12300) r502 <= _26215;
  wire [1:0] _26216 = {_0, _1151} + {_0, _2399};
  wire [1:0] _26217 = {_0, _5949} + {_0, _6973};
  wire [2:0] _26218 = {_0, _26216} + {_0, _26217};
  wire [1:0] _26219 = {_0, _9790} + {_0, _11004};
  wire [3:0] _26220 = {_0, _26218} + {_0, _0, _26219};
  wire _26221 = _12301 < _26220;
  wire _26222 = r501 ^ _26221;
  wire _26223 = _12298 ? coded_block[501] : r501;
  wire _26224 = _12296 ? _26222 : _26223;
  always @ (posedge reset or posedge clock) if (reset) r501 <= 1'd0; else if (_12300) r501 <= _26224;
  wire [1:0] _26225 = {_0, _1184} + {_0, _3486};
  wire [1:0] _26226 = {_0, _4478} + {_0, _8028};
  wire [2:0] _26227 = {_0, _26225} + {_0, _26226};
  wire [1:0] _26228 = {_0, _9054} + {_0, _11869};
  wire [3:0] _26229 = {_0, _26227} + {_0, _0, _26228};
  wire _26230 = _12301 < _26229;
  wire _26231 = r500 ^ _26230;
  wire _26232 = _12298 ? coded_block[500] : r500;
  wire _26233 = _12296 ? _26231 : _26232;
  always @ (posedge reset or posedge clock) if (reset) r500 <= 1'd0; else if (_12300) r500 <= _26233;
  wire [1:0] _26234 = {_0, _1215} + {_0, _3805};
  wire [1:0] _26235 = {_0, _5565} + {_0, _6558};
  wire [2:0] _26236 = {_0, _26234} + {_0, _26235};
  wire [1:0] _26237 = {_0, _10108} + {_0, _11132};
  wire [3:0] _26238 = {_0, _26236} + {_0, _0, _26237};
  wire _26239 = _12301 < _26238;
  wire _26240 = r499 ^ _26239;
  wire _26241 = _12298 ? coded_block[499] : r499;
  wire _26242 = _12296 ? _26240 : _26241;
  always @ (posedge reset or posedge clock) if (reset) r499 <= 1'd0; else if (_12300) r499 <= _26242;
  wire [1:0] _26243 = {_0, _1247} + {_0, _2239};
  wire [1:0] _26244 = {_0, _5884} + {_0, _7644};
  wire [2:0] _26245 = {_0, _26243} + {_0, _26244};
  wire [1:0] _26246 = {_0, _8638} + {_0, _12188};
  wire [3:0] _26247 = {_0, _26245} + {_0, _0, _26246};
  wire _26248 = _12301 < _26247;
  wire _26249 = r498 ^ _26248;
  wire _26250 = _12298 ? coded_block[498] : r498;
  wire _26251 = _12296 ? _26249 : _26250;
  always @ (posedge reset or posedge clock) if (reset) r498 <= 1'd0; else if (_12300) r498 <= _26251;
  wire [1:0] _26252 = {_0, _1278} + {_0, _3615};
  wire [1:0] _26253 = {_0, _4319} + {_0, _7965};
  wire [2:0] _26254 = {_0, _26252} + {_0, _26253};
  wire [1:0] _26255 = {_0, _9724} + {_0, _10717};
  wire [3:0] _26256 = {_0, _26254} + {_0, _0, _26255};
  wire _26257 = _12301 < _26256;
  wire _26258 = r497 ^ _26257;
  wire _26259 = _12298 ? coded_block[497] : r497;
  wire _26260 = _12296 ? _26258 : _26259;
  always @ (posedge reset or posedge clock) if (reset) r497 <= 1'd0; else if (_12300) r497 <= _26260;
  wire [1:0] _26261 = {_0, _1312} + {_0, _2526};
  wire [1:0] _26262 = {_0, _5694} + {_0, _6397};
  wire [2:0] _26263 = {_0, _26261} + {_0, _26262};
  wire [1:0] _26264 = {_0, _10045} + {_0, _11806};
  wire [3:0] _26265 = {_0, _26263} + {_0, _0, _26264};
  wire _26266 = _12301 < _26265;
  wire _26267 = r496 ^ _26266;
  wire _26268 = _12298 ? coded_block[496] : r496;
  wire _26269 = _12296 ? _26267 : _26268;
  always @ (posedge reset or posedge clock) if (reset) r496 <= 1'd0; else if (_12300) r496 <= _26269;
  wire [1:0] _26270 = {_0, _1343} + {_0, _2623};
  wire [1:0] _26271 = {_0, _4605} + {_0, _7773};
  wire [2:0] _26272 = {_0, _26270} + {_0, _26271};
  wire [1:0] _26273 = {_0, _8480} + {_0, _12124};
  wire [3:0] _26274 = {_0, _26272} + {_0, _0, _26273};
  wire _26275 = _12301 < _26274;
  wire _26276 = r495 ^ _26275;
  wire _26277 = _12298 ? coded_block[495] : r495;
  wire _26278 = _12296 ? _26276 : _26277;
  always @ (posedge reset or posedge clock) if (reset) r495 <= 1'd0; else if (_12300) r495 <= _26278;
  wire [1:0] _26279 = {_0, _1375} + {_0, _4091};
  wire [1:0] _26280 = {_0, _4703} + {_0, _6687};
  wire [2:0] _26281 = {_0, _26279} + {_0, _26280};
  wire [1:0] _26282 = {_0, _9853} + {_0, _10558};
  wire [3:0] _26283 = {_0, _26281} + {_0, _0, _26282};
  wire _26284 = _12301 < _26283;
  wire _26285 = r494 ^ _26284;
  wire _26286 = _12298 ? coded_block[494] : r494;
  wire _26287 = _12296 ? _26285 : _26286;
  always @ (posedge reset or posedge clock) if (reset) r494 <= 1'd0; else if (_12300) r494 <= _26287;
  wire [1:0] _26288 = {_0, _1406} + {_0, _2336};
  wire [1:0] _26289 = {_0, _4160} + {_0, _6781};
  wire [2:0] _26290 = {_0, _26288} + {_0, _26289};
  wire [1:0] _26291 = {_0, _8767} + {_0, _11933};
  wire [3:0] _26292 = {_0, _26290} + {_0, _0, _26291};
  wire _26293 = _12301 < _26292;
  wire _26294 = r493 ^ _26293;
  wire _26295 = _12298 ? coded_block[493] : r493;
  wire _26296 = _12296 ? _26294 : _26295;
  always @ (posedge reset or posedge clock) if (reset) r493 <= 1'd0; else if (_12300) r493 <= _26296;
  wire [1:0] _26297 = {_0, _1439} + {_0, _3231};
  wire [1:0] _26298 = {_0, _4415} + {_0, _6239};
  wire [2:0] _26299 = {_0, _26297} + {_0, _26298};
  wire [1:0] _26300 = {_0, _8863} + {_0, _10846};
  wire [3:0] _26301 = {_0, _26299} + {_0, _0, _26300};
  wire _26302 = _12301 < _26301;
  wire _26303 = r492 ^ _26302;
  wire _26304 = _12298 ? coded_block[492] : r492;
  wire _26305 = _12296 ? _26303 : _26304;
  always @ (posedge reset or posedge clock) if (reset) r492 <= 1'd0; else if (_12300) r492 <= _26305;
  wire [1:0] _26306 = {_0, _1470} + {_0, _2878};
  wire [1:0] _26307 = {_0, _5310} + {_0, _6494};
  wire [2:0] _26308 = {_0, _26306} + {_0, _26307};
  wire [1:0] _26309 = {_0, _8319} + {_0, _10941};
  wire [3:0] _26310 = {_0, _26308} + {_0, _0, _26309};
  wire _26311 = _12301 < _26310;
  wire _26312 = r491 ^ _26311;
  wire _26313 = _12298 ? coded_block[491] : r491;
  wire _26314 = _12296 ? _26312 : _26313;
  always @ (posedge reset or posedge clock) if (reset) r491 <= 1'd0; else if (_12300) r491 <= _26314;
  wire [1:0] _26315 = {_0, _1502} + {_0, _3104};
  wire [1:0] _26316 = {_0, _4958} + {_0, _7389};
  wire [2:0] _26317 = {_0, _26315} + {_0, _26316};
  wire [1:0] _26318 = {_0, _8574} + {_0, _10399};
  wire [3:0] _26319 = {_0, _26317} + {_0, _0, _26318};
  wire _26320 = _12301 < _26319;
  wire _26321 = r490 ^ _26320;
  wire _26322 = _12298 ? coded_block[490] : r490;
  wire _26323 = _12296 ? _26321 : _26322;
  always @ (posedge reset or posedge clock) if (reset) r490 <= 1'd0; else if (_12300) r490 <= _26323;
  wire [1:0] _26324 = {_0, _1533} + {_0, _2974};
  wire [1:0] _26325 = {_0, _5183} + {_0, _7036};
  wire [2:0] _26326 = {_0, _26324} + {_0, _26325};
  wire [1:0] _26327 = {_0, _9469} + {_0, _10654};
  wire [3:0] _26328 = {_0, _26326} + {_0, _0, _26327};
  wire _26329 = _12301 < _26328;
  wire _26330 = r489 ^ _26329;
  wire _26331 = _12298 ? coded_block[489] : r489;
  wire _26332 = _12296 ? _26330 : _26331;
  always @ (posedge reset or posedge clock) if (reset) r489 <= 1'd0; else if (_12300) r489 <= _26332;
  wire [1:0] _26333 = {_0, _1568} + {_0, _3325};
  wire [1:0] _26334 = {_0, _5053} + {_0, _7262};
  wire [2:0] _26335 = {_0, _26333} + {_0, _26334};
  wire [1:0] _26336 = {_0, _9118} + {_0, _11550};
  wire [3:0] _26337 = {_0, _26335} + {_0, _0, _26336};
  wire _26338 = _12301 < _26337;
  wire _26339 = r488 ^ _26338;
  wire _26340 = _12298 ? coded_block[488] : r488;
  wire _26341 = _12296 ? _26339 : _26340;
  always @ (posedge reset or posedge clock) if (reset) r488 <= 1'd0; else if (_12300) r488 <= _26341;
  wire [1:0] _26342 = {_0, _1599} + {_0, _4060};
  wire [1:0] _26343 = {_0, _5407} + {_0, _7132};
  wire [2:0] _26344 = {_0, _26342} + {_0, _26343};
  wire [1:0] _26345 = {_0, _9342} + {_0, _11196};
  wire [3:0] _26346 = {_0, _26344} + {_0, _0, _26345};
  wire _26347 = _12301 < _26346;
  wire _26348 = r487 ^ _26347;
  wire _26349 = _12298 ? coded_block[487] : r487;
  wire _26350 = _12296 ? _26348 : _26349;
  always @ (posedge reset or posedge clock) if (reset) r487 <= 1'd0; else if (_12300) r487 <= _26350;
  wire [1:0] _26351 = {_0, _1631} + {_0, _2655};
  wire [1:0] _26352 = {_0, _6139} + {_0, _7485};
  wire [2:0] _26353 = {_0, _26351} + {_0, _26352};
  wire [1:0] _26354 = {_0, _9212} + {_0, _11422};
  wire [3:0] _26355 = {_0, _26353} + {_0, _0, _26354};
  wire _26356 = _12301 < _26355;
  wire _26357 = r486 ^ _26356;
  wire _26358 = _12298 ? coded_block[486] : r486;
  wire _26359 = _12296 ? _26357 : _26358;
  always @ (posedge reset or posedge clock) if (reset) r486 <= 1'd0; else if (_12300) r486 <= _26359;
  wire [1:0] _26360 = {_0, _1662} + {_0, _2208};
  wire [1:0] _26361 = {_0, _4734} + {_0, _6207};
  wire [2:0] _26362 = {_0, _26360} + {_0, _26361};
  wire [1:0] _26363 = {_0, _9566} + {_0, _11295};
  wire [3:0] _26364 = {_0, _26362} + {_0, _0, _26363};
  wire _26365 = _12301 < _26364;
  wire _26366 = r485 ^ _26365;
  wire _26367 = _12298 ? coded_block[485] : r485;
  wire _26368 = _12296 ? _26366 : _26367;
  always @ (posedge reset or posedge clock) if (reset) r485 <= 1'd0; else if (_12300) r485 <= _26368;
  wire [1:0] _26369 = {_0, _1726} + {_0, _2847};
  wire [1:0] _26370 = {_0, _5918} + {_0, _6366};
  wire [2:0] _26371 = {_0, _26369} + {_0, _26370};
  wire [1:0] _26372 = {_0, _8894} + {_0, _10366};
  wire [3:0] _26373 = {_0, _26371} + {_0, _0, _26372};
  wire _26374 = _12301 < _26373;
  wire _26375 = r484 ^ _26374;
  wire _26376 = _12298 ? coded_block[484] : r484;
  wire _26377 = _12296 ? _26375 : _26376;
  always @ (posedge reset or posedge clock) if (reset) r484 <= 1'd0; else if (_12300) r484 <= _26377;
  wire [1:0] _26378 = {_0, _1789} + {_0, _3742};
  wire [1:0] _26379 = {_0, _5342} + {_0, _7005};
  wire [2:0] _26380 = {_0, _26378} + {_0, _26379};
  wire [1:0] _26381 = {_0, _10077} + {_0, _10527};
  wire [3:0] _26382 = {_0, _26380} + {_0, _0, _26381};
  wire _26383 = _12301 < _26382;
  wire _26384 = r483 ^ _26383;
  wire _26385 = _12298 ? coded_block[483] : r483;
  wire _26386 = _12296 ? _26384 : _26385;
  always @ (posedge reset or posedge clock) if (reset) r483 <= 1'd0; else if (_12300) r483 <= _26386;
  wire [1:0] _26387 = {_0, _1823} + {_0, _3167};
  wire [1:0] _26388 = {_0, _5821} + {_0, _7420};
  wire [2:0] _26389 = {_0, _26387} + {_0, _26388};
  wire [1:0] _26390 = {_0, _9085} + {_0, _12155};
  wire [3:0] _26391 = {_0, _26389} + {_0, _0, _26390};
  wire _26392 = _12301 < _26391;
  wire _26393 = r482 ^ _26392;
  wire _26394 = _12298 ? coded_block[482] : r482;
  wire _26395 = _12296 ? _26393 : _26394;
  always @ (posedge reset or posedge clock) if (reset) r482 <= 1'd0; else if (_12300) r482 <= _26395;
  wire [1:0] _26396 = {_0, _1854} + {_0, _2463};
  wire [1:0] _26397 = {_0, _5246} + {_0, _7900};
  wire [2:0] _26398 = {_0, _26396} + {_0, _26397};
  wire [1:0] _26399 = {_0, _9503} + {_0, _11165};
  wire [3:0] _26400 = {_0, _26398} + {_0, _0, _26399};
  wire _26401 = _12301 < _26400;
  wire _26402 = r481 ^ _26401;
  wire _26403 = _12298 ? coded_block[481] : r481;
  wire _26404 = _12296 ? _26402 : _26403;
  always @ (posedge reset or posedge clock) if (reset) r481 <= 1'd0; else if (_12300) r481 <= _26404;
  wire [1:0] _26405 = {_0, _1886} + {_0, _2144};
  wire [1:0] _26406 = {_0, _4542} + {_0, _7326};
  wire [2:0] _26407 = {_0, _26405} + {_0, _26406};
  wire [1:0] _26408 = {_0, _9980} + {_0, _11581};
  wire [3:0] _26409 = {_0, _26407} + {_0, _0, _26408};
  wire _26410 = _12301 < _26409;
  wire _26411 = r480 ^ _26410;
  wire _26412 = _12298 ? coded_block[480] : r480;
  wire _26413 = _12296 ? _26411 : _26412;
  always @ (posedge reset or posedge clock) if (reset) r480 <= 1'd0; else if (_12300) r480 <= _26413;
  wire [1:0] _26414 = {_0, _1917} + {_0, _2302};
  wire [1:0] _26415 = {_0, _4223} + {_0, _6621};
  wire [2:0] _26416 = {_0, _26414} + {_0, _26415};
  wire [1:0] _26417 = {_0, _9406} + {_0, _12061};
  wire [3:0] _26418 = {_0, _26416} + {_0, _0, _26417};
  wire _26419 = _12301 < _26418;
  wire _26420 = r479 ^ _26419;
  wire _26421 = _12298 ? coded_block[479] : r479;
  wire _26422 = _12296 ? _26420 : _26421;
  always @ (posedge reset or posedge clock) if (reset) r479 <= 1'd0; else if (_12300) r479 <= _26422;
  wire [1:0] _26423 = {_0, _1950} + {_0, _2112};
  wire [1:0] _26424 = {_0, _4384} + {_0, _6303};
  wire [2:0] _26425 = {_0, _26423} + {_0, _26424};
  wire [1:0] _26426 = {_0, _8701} + {_0, _11485};
  wire [3:0] _26427 = {_0, _26425} + {_0, _0, _26426};
  wire _26428 = _12301 < _26427;
  wire _26429 = r478 ^ _26428;
  wire _26430 = _12298 ? coded_block[478] : r478;
  wire _26431 = _12296 ? _26429 : _26430;
  always @ (posedge reset or posedge clock) if (reset) r478 <= 1'd0; else if (_12300) r478 <= _26431;
  wire [1:0] _26432 = {_0, _1981} + {_0, _2494};
  wire [1:0] _26433 = {_0, _4192} + {_0, _6462};
  wire [2:0] _26434 = {_0, _26432} + {_0, _26433};
  wire [1:0] _26435 = {_0, _8383} + {_0, _10783};
  wire [3:0] _26436 = {_0, _26434} + {_0, _0, _26435};
  wire _26437 = _12301 < _26436;
  wire _26438 = r477 ^ _26437;
  wire _26439 = _12298 ? coded_block[477] : r477;
  wire _26440 = _12296 ? _26438 : _26439;
  always @ (posedge reset or posedge clock) if (reset) r477 <= 1'd0; else if (_12300) r477 <= _26440;
  wire [1:0] _26441 = {_0, _65} + {_0, _3997};
  wire [1:0] _26442 = {_0, _5501} + {_0, _7804};
  wire [2:0] _26443 = {_0, _26441} + {_0, _26442};
  wire [1:0] _26444 = {_0, _8736} + {_0, _10430};
  wire [3:0] _26445 = {_0, _26443} + {_0, _0, _26444};
  wire _26446 = _12301 < _26445;
  wire _26447 = r476 ^ _26446;
  wire _26448 = _12298 ? coded_block[476] : r476;
  wire _26449 = _12296 ? _26447 : _26448;
  always @ (posedge reset or posedge clock) if (reset) r476 <= 1'd0; else if (_12300) r476 <= _26449;
  wire [1:0] _26450 = {_0, _97} + {_0, _3933};
  wire [1:0] _26451 = {_0, _6076} + {_0, _7581};
  wire [2:0] _26452 = {_0, _26450} + {_0, _26451};
  wire [1:0] _26453 = {_0, _9886} + {_0, _10814};
  wire [3:0] _26454 = {_0, _26452} + {_0, _0, _26453};
  wire _26455 = _12301 < _26454;
  wire _26456 = r475 ^ _26455;
  wire _26457 = _12298 ? coded_block[475] : r475;
  wire _26458 = _12296 ? _26456 : _26457;
  always @ (posedge reset or posedge clock) if (reset) r475 <= 1'd0; else if (_12300) r475 <= _26458;
  wire [1:0] _26459 = {_0, _128} + {_0, _3037};
  wire [1:0] _26460 = {_0, _6012} + {_0, _8155};
  wire [2:0] _26461 = {_0, _26459} + {_0, _26460};
  wire [1:0] _26462 = {_0, _9661} + {_0, _11964};
  wire [3:0] _26463 = {_0, _26461} + {_0, _0, _26462};
  wire _26464 = _12301 < _26463;
  wire _26465 = r474 ^ _26464;
  wire _26466 = _12298 ? coded_block[474] : r474;
  wire _26467 = _12296 ? _26465 : _26466;
  always @ (posedge reset or posedge clock) if (reset) r474 <= 1'd0; else if (_12300) r474 <= _26467;
  wire [1:0] _26468 = {_0, _161} + {_0, _3709};
  wire [1:0] _26469 = {_0, _5116} + {_0, _8092};
  wire [2:0] _26470 = {_0, _26468} + {_0, _26469};
  wire [1:0] _26471 = {_0, _10235} + {_0, _11740};
  wire [3:0] _26472 = {_0, _26470} + {_0, _0, _26471};
  wire _26473 = _12301 < _26472;
  wire _26474 = r473 ^ _26473;
  wire _26475 = _12298 ? coded_block[473] : r473;
  wire _26476 = _12296 ? _26474 : _26475;
  always @ (posedge reset or posedge clock) if (reset) r473 <= 1'd0; else if (_12300) r473 <= _26476;
  wire [1:0] _26477 = {_0, _192} + {_0, _3294};
  wire [1:0] _26478 = {_0, _5790} + {_0, _7199};
  wire [2:0] _26479 = {_0, _26477} + {_0, _26478};
  wire [1:0] _26480 = {_0, _10172} + {_0, _10303};
  wire [3:0] _26481 = {_0, _26479} + {_0, _0, _26480};
  wire _26482 = _12301 < _26481;
  wire _26483 = r472 ^ _26482;
  wire _26484 = _12298 ? coded_block[472] : r472;
  wire _26485 = _12296 ? _26483 : _26484;
  always @ (posedge reset or posedge clock) if (reset) r472 <= 1'd0; else if (_12300) r472 <= _26485;
  wire [1:0] _26486 = {_0, _224} + {_0, _3005};
  wire [1:0] _26487 = {_0, _5373} + {_0, _7868};
  wire [2:0] _26488 = {_0, _26486} + {_0, _26487};
  wire [1:0] _26489 = {_0, _9279} + {_0, _12251};
  wire [3:0] _26490 = {_0, _26488} + {_0, _0, _26489};
  wire _26491 = _12301 < _26490;
  wire _26492 = r471 ^ _26491;
  wire _26493 = _12298 ? coded_block[471] : r471;
  wire _26494 = _12296 ? _26492 : _26493;
  always @ (posedge reset or posedge clock) if (reset) r471 <= 1'd0; else if (_12300) r471 <= _26494;
  wire [1:0] _26495 = {_0, _255} + {_0, _3964};
  wire [1:0] _26496 = {_0, _5085} + {_0, _7454};
  wire [2:0] _26497 = {_0, _26495} + {_0, _26496};
  wire [1:0] _26498 = {_0, _9949} + {_0, _11358};
  wire [3:0] _26499 = {_0, _26497} + {_0, _0, _26498};
  wire _26500 = _12301 < _26499;
  wire _26501 = r470 ^ _26500;
  wire _26502 = _12298 ? coded_block[470] : r470;
  wire _26503 = _12296 ? _26501 : _26502;
  always @ (posedge reset or posedge clock) if (reset) r470 <= 1'd0; else if (_12300) r470 <= _26503;
  wire [1:0] _26504 = {_0, _289} + {_0, _3453};
  wire [1:0] _26505 = {_0, _6045} + {_0, _7163};
  wire [2:0] _26506 = {_0, _26504} + {_0, _26505};
  wire [1:0] _26507 = {_0, _9534} + {_0, _12027};
  wire [3:0] _26508 = {_0, _26506} + {_0, _0, _26507};
  wire _26509 = _12301 < _26508;
  wire _26510 = r469 ^ _26509;
  wire _26511 = _12298 ? coded_block[469] : r469;
  wire _26512 = _12296 ? _26510 : _26511;
  always @ (posedge reset or posedge clock) if (reset) r469 <= 1'd0; else if (_12300) r469 <= _26512;
  wire [1:0] _26513 = {_0, _320} + {_0, _2430};
  wire [1:0] _26514 = {_0, _5534} + {_0, _8123};
  wire [2:0] _26515 = {_0, _26513} + {_0, _26514};
  wire [1:0] _26516 = {_0, _9248} + {_0, _11613};
  wire [3:0] _26517 = {_0, _26515} + {_0, _0, _26516};
  wire _26518 = _12301 < _26517;
  wire _26519 = r468 ^ _26518;
  wire _26520 = _12298 ? coded_block[468] : r468;
  wire _26521 = _12296 ? _26519 : _26520;
  always @ (posedge reset or posedge clock) if (reset) r468 <= 1'd0; else if (_12300) r468 <= _26521;
  wire [1:0] _26522 = {_0, _352} + {_0, _3198};
  wire [1:0] _26523 = {_0, _4511} + {_0, _7612};
  wire [2:0] _26524 = {_0, _26522} + {_0, _26523};
  wire [1:0] _26525 = {_0, _10204} + {_0, _11326};
  wire [3:0] _26526 = {_0, _26524} + {_0, _0, _26525};
  wire _26527 = _12301 < _26526;
  wire _26528 = r467 ^ _26527;
  wire _26529 = _12298 ? coded_block[467] : r467;
  wire _26530 = _12296 ? _26528 : _26529;
  always @ (posedge reset or posedge clock) if (reset) r467 <= 1'd0; else if (_12300) r467 <= _26530;
  wire [1:0] _26531 = {_0, _416} + {_0, _3901};
  wire [1:0] _26532 = {_0, _4447} + {_0, _7357};
  wire [2:0] _26533 = {_0, _26531} + {_0, _26532};
  wire [1:0] _26534 = {_0, _8670} + {_0, _11771};
  wire [3:0] _26535 = {_0, _26533} + {_0, _0, _26534};
  wire _26536 = _12301 < _26535;
  wire _26537 = r466 ^ _26536;
  wire _26538 = _12298 ? coded_block[466] : r466;
  wire _26539 = _12296 ? _26537 : _26538;
  always @ (posedge reset or posedge clock) if (reset) r466 <= 1'd0; else if (_12300) r466 <= _26539;
  wire [1:0] _26540 = {_0, _447} + {_0, _4028};
  wire [1:0] _26541 = {_0, _5981} + {_0, _6525};
  wire [2:0] _26542 = {_0, _26540} + {_0, _26541};
  wire [1:0] _26543 = {_0, _9438} + {_0, _10748};
  wire [3:0] _26544 = {_0, _26542} + {_0, _0, _26543};
  wire _26545 = _12301 < _26544;
  wire _26546 = r465 ^ _26545;
  wire _26547 = _12298 ? coded_block[465] : r465;
  wire _26548 = _12296 ? _26546 : _26547;
  always @ (posedge reset or posedge clock) if (reset) r465 <= 1'd0; else if (_12300) r465 <= _26548;
  wire [1:0] _26549 = {_0, _479} + {_0, _3359};
  wire [1:0] _26550 = {_0, _6108} + {_0, _8059};
  wire [2:0] _26551 = {_0, _26549} + {_0, _26550};
  wire [1:0] _26552 = {_0, _8607} + {_0, _11516};
  wire [3:0] _26553 = {_0, _26551} + {_0, _0, _26552};
  wire _26554 = _12301 < _26553;
  wire _26555 = r464 ^ _26554;
  wire _26556 = _12298 ? coded_block[464] : r464;
  wire _26557 = _12296 ? _26555 : _26556;
  always @ (posedge reset or posedge clock) if (reset) r464 <= 1'd0; else if (_12300) r464 <= _26557;
  wire [1:0] _26558 = {_0, _545} + {_0, _2557};
  wire [1:0] _26559 = {_0, _4671} + {_0, _7517};
  wire [2:0] _26560 = {_0, _26558} + {_0, _26559};
  wire [1:0] _26561 = {_0, _8256} + {_0, _12219};
  wire [3:0] _26562 = {_0, _26560} + {_0, _0, _26561};
  wire _26563 = _12301 < _26562;
  wire _26564 = r463 ^ _26563;
  wire _26565 = _12298 ? coded_block[463] : r463;
  wire _26566 = _12296 ? _26564 : _26565;
  always @ (posedge reset or posedge clock) if (reset) r463 <= 1'd0; else if (_12300) r463 <= _26566;
  wire [1:0] _26567 = {_0, _576} + {_0, _3390};
  wire [1:0] _26568 = {_0, _4640} + {_0, _6750};
  wire [2:0] _26569 = {_0, _26567} + {_0, _26568};
  wire [1:0] _26570 = {_0, _9597} + {_0, _10335};
  wire [3:0] _26571 = {_0, _26569} + {_0, _0, _26570};
  wire _26572 = _12301 < _26571;
  wire _26573 = r462 ^ _26572;
  wire _26574 = _12298 ? coded_block[462] : r462;
  wire _26575 = _12296 ? _26573 : _26574;
  always @ (posedge reset or posedge clock) if (reset) r462 <= 1'd0; else if (_12300) r462 <= _26575;
  wire [1:0] _26576 = {_0, _608} + {_0, _3678};
  wire [1:0] _26577 = {_0, _5470} + {_0, _6718};
  wire [2:0] _26578 = {_0, _26576} + {_0, _26577};
  wire [1:0] _26579 = {_0, _8830} + {_0, _11677};
  wire [3:0] _26580 = {_0, _26578} + {_0, _0, _26579};
  wire _26581 = _12301 < _26580;
  wire _26582 = r461 ^ _26581;
  wire _26583 = _12298 ? coded_block[461] : r461;
  wire _26584 = _12296 ? _26582 : _26583;
  always @ (posedge reset or posedge clock) if (reset) r461 <= 1'd0; else if (_12300) r461 <= _26584;
  wire [1:0] _26585 = {_0, _639} + {_0, _3068};
  wire [1:0] _26586 = {_0, _5757} + {_0, _7548};
  wire [2:0] _26587 = {_0, _26585} + {_0, _26586};
  wire [1:0] _26588 = {_0, _8799} + {_0, _10910};
  wire [3:0] _26589 = {_0, _26587} + {_0, _0, _26588};
  wire _26590 = _12301 < _26589;
  wire _26591 = r460 ^ _26590;
  wire _26592 = _12298 ? coded_block[460] : r460;
  wire _26593 = _12296 ? _26591 : _26592;
  always @ (posedge reset or posedge clock) if (reset) r460 <= 1'd0; else if (_12300) r460 <= _26593;
  wire [1:0] _26594 = {_0, _672} + {_0, _2910};
  wire [1:0] _26595 = {_0, _5152} + {_0, _7837};
  wire [2:0] _26596 = {_0, _26594} + {_0, _26595};
  wire [1:0] _26597 = {_0, _9630} + {_0, _10877};
  wire [3:0] _26598 = {_0, _26596} + {_0, _0, _26597};
  wire _26599 = _12301 < _26598;
  wire _26600 = r459 ^ _26599;
  wire _26601 = _12298 ? coded_block[459] : r459;
  wire _26602 = _12296 ? _26600 : _26601;
  always @ (posedge reset or posedge clock) if (reset) r459 <= 1'd0; else if (_12300) r459 <= _26602;
  wire [1:0] _26603 = {_0, _703} + {_0, _2081};
  wire [1:0] _26604 = {_0, _4989} + {_0, _7230};
  wire [2:0] _26605 = {_0, _26603} + {_0, _26604};
  wire [1:0] _26606 = {_0, _9917} + {_0, _11708};
  wire [3:0] _26607 = {_0, _26605} + {_0, _0, _26606};
  wire _26608 = _12301 < _26607;
  wire _26609 = r458 ^ _26608;
  wire _26610 = _12298 ? coded_block[458] : r458;
  wire _26611 = _12296 ? _26609 : _26610;
  always @ (posedge reset or posedge clock) if (reset) r458 <= 1'd0; else if (_12300) r458 <= _26611;
  wire [1:0] _26612 = {_0, _735} + {_0, _2941};
  wire [1:0] _26613 = {_0, _4129} + {_0, _7069};
  wire [2:0] _26614 = {_0, _26612} + {_0, _26613};
  wire [1:0] _26615 = {_0, _9311} + {_0, _11996};
  wire [3:0] _26616 = {_0, _26614} + {_0, _0, _26615};
  wire _26617 = _12301 < _26616;
  wire _26618 = r457 ^ _26617;
  wire _26619 = _12298 ? coded_block[457] : r457;
  wire _26620 = _12296 ? _26618 : _26619;
  always @ (posedge reset or posedge clock) if (reset) r457 <= 1'd0; else if (_12300) r457 <= _26620;
  wire [1:0] _26621 = {_0, _766} + {_0, _3135};
  wire [1:0] _26622 = {_0, _5022} + {_0, _6176};
  wire [2:0] _26623 = {_0, _26621} + {_0, _26622};
  wire [1:0] _26624 = {_0, _9149} + {_0, _11389};
  wire [3:0] _26625 = {_0, _26623} + {_0, _0, _26624};
  wire _26626 = _12301 < _26625;
  wire _26627 = r456 ^ _26626;
  wire _26628 = _12298 ? coded_block[456] : r456;
  wire _26629 = _12296 ? _26627 : _26628;
  always @ (posedge reset or posedge clock) if (reset) r456 <= 1'd0; else if (_12300) r456 <= _26629;
  wire [1:0] _26630 = {_0, _800} + {_0, _3773};
  wire [1:0] _26631 = {_0, _5215} + {_0, _7100};
  wire [2:0] _26632 = {_0, _26630} + {_0, _26631};
  wire [1:0] _26633 = {_0, _8225} + {_0, _11228};
  wire [3:0] _26634 = {_0, _26632} + {_0, _0, _26633};
  wire _26635 = _12301 < _26634;
  wire _26636 = r455 ^ _26635;
  wire _26637 = _12298 ? coded_block[455] : r455;
  wire _26638 = _12296 ? _26636 : _26637;
  always @ (posedge reset or posedge clock) if (reset) r455 <= 1'd0; else if (_12300) r455 <= _26638;
  wire [1:0] _26639 = {_0, _831} + {_0, _3517};
  wire [1:0] _26640 = {_0, _5853} + {_0, _7293};
  wire [2:0] _26641 = {_0, _26639} + {_0, _26640};
  wire [1:0] _26642 = {_0, _9181} + {_0, _10272};
  wire [3:0] _26643 = {_0, _26641} + {_0, _0, _26642};
  wire _26644 = _12301 < _26643;
  wire _26645 = r454 ^ _26644;
  wire _26646 = _12298 ? coded_block[454] : r454;
  wire _26647 = _12296 ? _26645 : _26646;
  always @ (posedge reset or posedge clock) if (reset) r454 <= 1'd0; else if (_12300) r454 <= _26647;
  wire [1:0] _26648 = {_0, _863} + {_0, _2719};
  wire [1:0] _26649 = {_0, _5597} + {_0, _7931};
  wire [2:0] _26650 = {_0, _26648} + {_0, _26649};
  wire [1:0] _26651 = {_0, _9375} + {_0, _11259};
  wire [3:0] _26652 = {_0, _26650} + {_0, _0, _26651};
  wire _26653 = _12301 < _26652;
  wire _26654 = r453 ^ _26653;
  wire _26655 = _12298 ? coded_block[453] : r453;
  wire _26656 = _12296 ? _26654 : _26655;
  always @ (posedge reset or posedge clock) if (reset) r453 <= 1'd0; else if (_12300) r453 <= _26656;
  wire [1:0] _26657 = {_0, _894} + {_0, _2782};
  wire [1:0] _26658 = {_0, _4798} + {_0, _7675};
  wire [2:0] _26659 = {_0, _26657} + {_0, _26658};
  wire [1:0] _26660 = {_0, _10014} + {_0, _11453};
  wire [3:0] _26661 = {_0, _26659} + {_0, _0, _26660};
  wire _26662 = _12301 < _26661;
  wire _26663 = r452 ^ _26662;
  wire _26664 = _12298 ? coded_block[452] : r452;
  wire _26665 = _12296 ? _26663 : _26664;
  always @ (posedge reset or posedge clock) if (reset) r452 <= 1'd0; else if (_12300) r452 <= _26665;
  wire [1:0] _26666 = {_0, _927} + {_0, _3580};
  wire [1:0] _26667 = {_0, _4861} + {_0, _6877};
  wire [2:0] _26668 = {_0, _26666} + {_0, _26667};
  wire [1:0] _26669 = {_0, _9759} + {_0, _12092};
  wire [3:0] _26670 = {_0, _26668} + {_0, _0, _26669};
  wire _26671 = _12301 < _26670;
  wire _26672 = r451 ^ _26671;
  wire _26673 = _12298 ? coded_block[451] : r451;
  wire _26674 = _12296 ? _26672 : _26673;
  always @ (posedge reset or posedge clock) if (reset) r451 <= 1'd0; else if (_12300) r451 <= _26674;
  wire [1:0] _26675 = {_0, _958} + {_0, _2271};
  wire [1:0] _26676 = {_0, _5663} + {_0, _6942};
  wire [2:0] _26677 = {_0, _26675} + {_0, _26676};
  wire [1:0] _26678 = {_0, _8957} + {_0, _11837};
  wire [3:0] _26679 = {_0, _26677} + {_0, _0, _26678};
  wire _26680 = _12301 < _26679;
  wire _26681 = r450 ^ _26680;
  wire _26682 = _12298 ? coded_block[450] : r450;
  wire _26683 = _12296 ? _26681 : _26682;
  always @ (posedge reset or posedge clock) if (reset) r450 <= 1'd0; else if (_12300) r450 <= _26683;
  wire [1:0] _26684 = {_0, _990} + {_0, _2175};
  wire [1:0] _26685 = {_0, _4350} + {_0, _7741};
  wire [2:0] _26686 = {_0, _26684} + {_0, _26685};
  wire [1:0] _26687 = {_0, _9022} + {_0, _11038};
  wire [3:0] _26688 = {_0, _26686} + {_0, _0, _26687};
  wire _26689 = _12301 < _26688;
  wire _26690 = r449 ^ _26689;
  wire _26691 = _12298 ? coded_block[449] : r449;
  wire _26692 = _12296 ? _26690 : _26691;
  always @ (posedge reset or posedge clock) if (reset) r449 <= 1'd0; else if (_12300) r449 <= _26692;
  wire [1:0] _26693 = {_0, _1021} + {_0, _2686};
  wire [1:0] _26694 = {_0, _4256} + {_0, _6431};
  wire [2:0] _26695 = {_0, _26693} + {_0, _26694};
  wire [1:0] _26696 = {_0, _9822} + {_0, _11101};
  wire [3:0] _26697 = {_0, _26695} + {_0, _0, _26696};
  wire _26698 = _12301 < _26697;
  wire _26699 = r448 ^ _26698;
  wire _26700 = _12298 ? coded_block[448] : r448;
  wire _26701 = _12296 ? _26699 : _26700;
  always @ (posedge reset or posedge clock) if (reset) r448 <= 1'd0; else if (_12300) r448 <= _26701;
  wire [1:0] _26702 = {_0, _34} + {_0, _2910};
  wire [1:0] _26703 = {_0, _4989} + {_0, _7069};
  wire [2:0] _26704 = {_0, _26702} + {_0, _26703};
  wire [1:0] _26705 = {_0, _9149} + {_0, _11228};
  wire [3:0] _26706 = {_0, _26704} + {_0, _0, _26705};
  wire _26707 = _12301 < _26706;
  wire _26708 = r447 ^ _26707;
  wire _26709 = _12298 ? coded_block[447] : r447;
  wire _26710 = _12296 ? _26708 : _26709;
  always @ (posedge reset or posedge clock) if (reset) r447 <= 1'd0; else if (_12300) r447 <= _26710;
  wire [1:0] _26711 = {_0, _735} + {_0, _3549};
  wire [1:0] _26712 = {_0, _4798} + {_0, _6908};
  wire [2:0] _26713 = {_0, _26711} + {_0, _26712};
  wire [1:0] _26714 = {_0, _9759} + {_0, _10493};
  wire [3:0] _26715 = {_0, _26713} + {_0, _0, _26714};
  wire _26716 = _12301 < _26715;
  wire _26717 = r446 ^ _26716;
  wire _26718 = _12298 ? coded_block[446] : r446;
  wire _26719 = _12296 ? _26717 : _26718;
  always @ (posedge reset or posedge clock) if (reset) r446 <= 1'd0; else if (_12300) r446 <= _26719;
  wire [1:0] _26720 = {_0, _766} + {_0, _3836};
  wire [1:0] _26721 = {_0, _5628} + {_0, _6877};
  wire [2:0] _26722 = {_0, _26720} + {_0, _26721};
  wire [1:0] _26723 = {_0, _8991} + {_0, _11837};
  wire [3:0] _26724 = {_0, _26722} + {_0, _0, _26723};
  wire _26725 = _12301 < _26724;
  wire _26726 = r445 ^ _26725;
  wire _26727 = _12298 ? coded_block[445] : r445;
  wire _26728 = _12296 ? _26726 : _26727;
  always @ (posedge reset or posedge clock) if (reset) r445 <= 1'd0; else if (_12300) r445 <= _26728;
  wire [1:0] _26729 = {_0, _800} + {_0, _3231};
  wire [1:0] _26730 = {_0, _5918} + {_0, _7710};
  wire [2:0] _26731 = {_0, _26729} + {_0, _26730};
  wire [1:0] _26732 = {_0, _8957} + {_0, _11069};
  wire [3:0] _26733 = {_0, _26731} + {_0, _0, _26732};
  wire _26734 = _12301 < _26733;
  wire _26735 = r444 ^ _26734;
  wire _26736 = _12298 ? coded_block[444] : r444;
  wire _26737 = _12296 ? _26735 : _26736;
  always @ (posedge reset or posedge clock) if (reset) r444 <= 1'd0; else if (_12300) r444 <= _26737;
  wire [1:0] _26738 = {_0, _831} + {_0, _3068};
  wire [1:0] _26739 = {_0, _5310} + {_0, _7996};
  wire [2:0] _26740 = {_0, _26738} + {_0, _26739};
  wire [1:0] _26741 = {_0, _9790} + {_0, _11038};
  wire [3:0] _26742 = {_0, _26740} + {_0, _0, _26741};
  wire _26743 = _12301 < _26742;
  wire _26744 = r443 ^ _26743;
  wire _26745 = _12298 ? coded_block[443] : r443;
  wire _26746 = _12296 ? _26744 : _26745;
  always @ (posedge reset or posedge clock) if (reset) r443 <= 1'd0; else if (_12300) r443 <= _26746;
  wire [1:0] _26747 = {_0, _863} + {_0, _2081};
  wire [1:0] _26748 = {_0, _5152} + {_0, _7389};
  wire [2:0] _26749 = {_0, _26747} + {_0, _26748};
  wire [1:0] _26750 = {_0, _10077} + {_0, _11869};
  wire [3:0] _26751 = {_0, _26749} + {_0, _0, _26750};
  wire _26752 = _12301 < _26751;
  wire _26753 = r442 ^ _26752;
  wire _26754 = _12298 ? coded_block[442] : r442;
  wire _26755 = _12296 ? _26753 : _26754;
  always @ (posedge reset or posedge clock) if (reset) r442 <= 1'd0; else if (_12300) r442 <= _26755;
  wire [1:0] _26756 = {_0, _894} + {_0, _3104};
  wire [1:0] _26757 = {_0, _4129} + {_0, _7230};
  wire [2:0] _26758 = {_0, _26756} + {_0, _26757};
  wire [1:0] _26759 = {_0, _9469} + {_0, _12155};
  wire [3:0] _26760 = {_0, _26758} + {_0, _0, _26759};
  wire _26761 = _12301 < _26760;
  wire _26762 = r441 ^ _26761;
  wire _26763 = _12298 ? coded_block[441] : r441;
  wire _26764 = _12296 ? _26762 : _26763;
  always @ (posedge reset or posedge clock) if (reset) r441 <= 1'd0; else if (_12300) r441 <= _26764;
  wire [1:0] _26765 = {_0, _927} + {_0, _3294};
  wire [1:0] _26766 = {_0, _5183} + {_0, _6176};
  wire [2:0] _26767 = {_0, _26765} + {_0, _26766};
  wire [1:0] _26768 = {_0, _9311} + {_0, _11550};
  wire [3:0] _26769 = {_0, _26767} + {_0, _0, _26768};
  wire _26770 = _12301 < _26769;
  wire _26771 = r440 ^ _26770;
  wire _26772 = _12298 ? coded_block[440] : r440;
  wire _26773 = _12296 ? _26771 : _26772;
  always @ (posedge reset or posedge clock) if (reset) r440 <= 1'd0; else if (_12300) r440 <= _26773;
  wire [1:0] _26774 = {_0, _990} + {_0, _3678};
  wire [1:0] _26775 = {_0, _6012} + {_0, _7454};
  wire [2:0] _26776 = {_0, _26774} + {_0, _26775};
  wire [1:0] _26777 = {_0, _9342} + {_0, _10272};
  wire [3:0] _26778 = {_0, _26776} + {_0, _0, _26777};
  wire _26779 = _12301 < _26778;
  wire _26780 = r439 ^ _26779;
  wire _26781 = _12298 ? coded_block[439] : r439;
  wire _26782 = _12296 ? _26780 : _26781;
  always @ (posedge reset or posedge clock) if (reset) r439 <= 1'd0; else if (_12300) r439 <= _26782;
  wire [1:0] _26783 = {_0, _1021} + {_0, _2878};
  wire [1:0] _26784 = {_0, _5757} + {_0, _8092};
  wire [2:0] _26785 = {_0, _26783} + {_0, _26784};
  wire [1:0] _26786 = {_0, _9534} + {_0, _11422};
  wire [3:0] _26787 = {_0, _26785} + {_0, _0, _26786};
  wire _26788 = _12301 < _26787;
  wire _26789 = r438 ^ _26788;
  wire _26790 = _12298 ? coded_block[438] : r438;
  wire _26791 = _12296 ? _26789 : _26790;
  always @ (posedge reset or posedge clock) if (reset) r438 <= 1'd0; else if (_12300) r438 <= _26791;
  wire [1:0] _26792 = {_0, _1088} + {_0, _3742};
  wire [1:0] _26793 = {_0, _5022} + {_0, _7036};
  wire [2:0] _26794 = {_0, _26792} + {_0, _26793};
  wire [1:0] _26795 = {_0, _9917} + {_0, _12251};
  wire [3:0] _26796 = {_0, _26794} + {_0, _0, _26795};
  wire _26797 = _12301 < _26796;
  wire _26798 = r437 ^ _26797;
  wire _26799 = _12298 ? coded_block[437] : r437;
  wire _26800 = _12296 ? _26798 : _26799;
  always @ (posedge reset or posedge clock) if (reset) r437 <= 1'd0; else if (_12300) r437 <= _26800;
  wire [1:0] _26801 = {_0, _1120} + {_0, _2430};
  wire [1:0] _26802 = {_0, _5821} + {_0, _7100};
  wire [2:0] _26803 = {_0, _26801} + {_0, _26802};
  wire [1:0] _26804 = {_0, _9118} + {_0, _11996};
  wire [3:0] _26805 = {_0, _26803} + {_0, _0, _26804};
  wire _26806 = _12301 < _26805;
  wire _26807 = r436 ^ _26806;
  wire _26808 = _12298 ? coded_block[436] : r436;
  wire _26809 = _12296 ? _26807 : _26808;
  always @ (posedge reset or posedge clock) if (reset) r436 <= 1'd0; else if (_12300) r436 <= _26809;
  wire [1:0] _26810 = {_0, _1151} + {_0, _2336};
  wire [1:0] _26811 = {_0, _4511} + {_0, _7900};
  wire [2:0] _26812 = {_0, _26810} + {_0, _26811};
  wire [1:0] _26813 = {_0, _9181} + {_0, _11196};
  wire [3:0] _26814 = {_0, _26812} + {_0, _0, _26813};
  wire _26815 = _12301 < _26814;
  wire _26816 = r435 ^ _26815;
  wire _26817 = _12298 ? coded_block[435] : r435;
  wire _26818 = _12296 ? _26816 : _26817;
  always @ (posedge reset or posedge clock) if (reset) r435 <= 1'd0; else if (_12300) r435 <= _26818;
  wire [1:0] _26819 = {_0, _1184} + {_0, _2847};
  wire [1:0] _26820 = {_0, _4415} + {_0, _6589};
  wire [2:0] _26821 = {_0, _26819} + {_0, _26820};
  wire [1:0] _26822 = {_0, _9980} + {_0, _11259};
  wire [3:0] _26823 = {_0, _26821} + {_0, _0, _26822};
  wire _26824 = _12301 < _26823;
  wire _26825 = r434 ^ _26824;
  wire _26826 = _12298 ? coded_block[434] : r434;
  wire _26827 = _12296 ? _26825 : _26826;
  always @ (posedge reset or posedge clock) if (reset) r434 <= 1'd0; else if (_12300) r434 <= _26827;
  wire [1:0] _26828 = {_0, _1215} + {_0, _3709};
  wire [1:0] _26829 = {_0, _4926} + {_0, _6494};
  wire [2:0] _26830 = {_0, _26828} + {_0, _26829};
  wire [1:0] _26831 = {_0, _8670} + {_0, _12061};
  wire [3:0] _26832 = {_0, _26830} + {_0, _0, _26831};
  wire _26833 = _12301 < _26832;
  wire _26834 = r433 ^ _26833;
  wire _26835 = _12298 ? coded_block[433] : r433;
  wire _26836 = _12296 ? _26834 : _26835;
  always @ (posedge reset or posedge clock) if (reset) r433 <= 1'd0; else if (_12300) r433 <= _26836;
  wire [1:0] _26837 = {_0, _1247} + {_0, _2974};
  wire [1:0] _26838 = {_0, _5790} + {_0, _7005};
  wire [2:0] _26839 = {_0, _26837} + {_0, _26838};
  wire [1:0] _26840 = {_0, _8574} + {_0, _10748};
  wire [3:0] _26841 = {_0, _26839} + {_0, _0, _26840};
  wire _26842 = _12301 < _26841;
  wire _26843 = r432 ^ _26842;
  wire _26844 = _12298 ? coded_block[432] : r432;
  wire _26845 = _12296 ? _26843 : _26844;
  always @ (posedge reset or posedge clock) if (reset) r432 <= 1'd0; else if (_12300) r432 <= _26845;
  wire [1:0] _26846 = {_0, _1278} + {_0, _4028};
  wire [1:0] _26847 = {_0, _5053} + {_0, _7868};
  wire [2:0] _26848 = {_0, _26846} + {_0, _26847};
  wire [1:0] _26849 = {_0, _9085} + {_0, _10654};
  wire [3:0] _26850 = {_0, _26848} + {_0, _0, _26849};
  wire _26851 = _12301 < _26850;
  wire _26852 = r431 ^ _26851;
  wire _26853 = _12298 ? coded_block[431] : r431;
  wire _26854 = _12296 ? _26852 : _26853;
  always @ (posedge reset or posedge clock) if (reset) r431 <= 1'd0; else if (_12300) r431 <= _26854;
  wire [1:0] _26855 = {_0, _1312} + {_0, _2557};
  wire [1:0] _26856 = {_0, _6108} + {_0, _7132};
  wire [2:0] _26857 = {_0, _26855} + {_0, _26856};
  wire [1:0] _26858 = {_0, _9949} + {_0, _11165};
  wire [3:0] _26859 = {_0, _26857} + {_0, _0, _26858};
  wire _26860 = _12301 < _26859;
  wire _26861 = r430 ^ _26860;
  wire _26862 = _12298 ? coded_block[430] : r430;
  wire _26863 = _12296 ? _26861 : _26862;
  always @ (posedge reset or posedge clock) if (reset) r430 <= 1'd0; else if (_12300) r430 <= _26863;
  wire [1:0] _26864 = {_0, _1343} + {_0, _3646};
  wire [1:0] _26865 = {_0, _4640} + {_0, _8186};
  wire [2:0] _26866 = {_0, _26864} + {_0, _26865};
  wire [1:0] _26867 = {_0, _9212} + {_0, _12027};
  wire [3:0] _26868 = {_0, _26866} + {_0, _0, _26867};
  wire _26869 = _12301 < _26868;
  wire _26870 = r429 ^ _26869;
  wire _26871 = _12298 ? coded_block[429] : r429;
  wire _26872 = _12296 ? _26870 : _26871;
  always @ (posedge reset or posedge clock) if (reset) r429 <= 1'd0; else if (_12300) r429 <= _26872;
  wire [1:0] _26873 = {_0, _1375} + {_0, _3964};
  wire [1:0] _26874 = {_0, _5726} + {_0, _6718};
  wire [2:0] _26875 = {_0, _26873} + {_0, _26874};
  wire [1:0] _26876 = {_0, _8256} + {_0, _11295};
  wire [3:0] _26877 = {_0, _26875} + {_0, _0, _26876};
  wire _26878 = _12301 < _26877;
  wire _26879 = r428 ^ _26878;
  wire _26880 = _12298 ? coded_block[428] : r428;
  wire _26881 = _12296 ? _26879 : _26880;
  always @ (posedge reset or posedge clock) if (reset) r428 <= 1'd0; else if (_12300) r428 <= _26881;
  wire [1:0] _26882 = {_0, _1406} + {_0, _2399};
  wire [1:0] _26883 = {_0, _6045} + {_0, _7804};
  wire [2:0] _26884 = {_0, _26882} + {_0, _26883};
  wire [1:0] _26885 = {_0, _8799} + {_0, _10335};
  wire [3:0] _26886 = {_0, _26884} + {_0, _0, _26885};
  wire _26887 = _12301 < _26886;
  wire _26888 = r427 ^ _26887;
  wire _26889 = _12298 ? coded_block[427] : r427;
  wire _26890 = _12296 ? _26888 : _26889;
  always @ (posedge reset or posedge clock) if (reset) r427 <= 1'd0; else if (_12300) r427 <= _26890;
  wire [1:0] _26891 = {_0, _1439} + {_0, _3773};
  wire [1:0] _26892 = {_0, _4478} + {_0, _8123};
  wire [2:0] _26893 = {_0, _26891} + {_0, _26892};
  wire [1:0] _26894 = {_0, _9886} + {_0, _10877};
  wire [3:0] _26895 = {_0, _26893} + {_0, _0, _26894};
  wire _26896 = _12301 < _26895;
  wire _26897 = r426 ^ _26896;
  wire _26898 = _12298 ? coded_block[426] : r426;
  wire _26899 = _12296 ? _26897 : _26898;
  always @ (posedge reset or posedge clock) if (reset) r426 <= 1'd0; else if (_12300) r426 <= _26899;
  wire [1:0] _26900 = {_0, _1470} + {_0, _2686};
  wire [1:0] _26901 = {_0, _5853} + {_0, _6558};
  wire [2:0] _26902 = {_0, _26900} + {_0, _26901};
  wire [1:0] _26903 = {_0, _10204} + {_0, _11964};
  wire [3:0] _26904 = {_0, _26902} + {_0, _0, _26903};
  wire _26905 = _12301 < _26904;
  wire _26906 = r425 ^ _26905;
  wire _26907 = _12298 ? coded_block[425] : r425;
  wire _26908 = _12296 ? _26906 : _26907;
  always @ (posedge reset or posedge clock) if (reset) r425 <= 1'd0; else if (_12300) r425 <= _26908;
  wire [1:0] _26909 = {_0, _1502} + {_0, _2782};
  wire [1:0] _26910 = {_0, _4767} + {_0, _7931};
  wire [2:0] _26911 = {_0, _26909} + {_0, _26910};
  wire [1:0] _26912 = {_0, _8638} + {_0, _12282};
  wire [3:0] _26913 = {_0, _26911} + {_0, _0, _26912};
  wire _26914 = _12301 < _26913;
  wire _26915 = r424 ^ _26914;
  wire _26916 = _12298 ? coded_block[424] : r424;
  wire _26917 = _12296 ? _26915 : _26916;
  always @ (posedge reset or posedge clock) if (reset) r424 <= 1'd0; else if (_12300) r424 <= _26917;
  wire [1:0] _26918 = {_0, _1568} + {_0, _2494};
  wire [1:0] _26919 = {_0, _4319} + {_0, _6942};
  wire [2:0] _26920 = {_0, _26918} + {_0, _26919};
  wire [1:0] _26921 = {_0, _8926} + {_0, _12092};
  wire [3:0] _26922 = {_0, _26920} + {_0, _0, _26921};
  wire _26923 = _12301 < _26922;
  wire _26924 = r423 ^ _26923;
  wire _26925 = _12298 ? coded_block[423] : r423;
  wire _26926 = _12296 ? _26924 : _26925;
  always @ (posedge reset or posedge clock) if (reset) r423 <= 1'd0; else if (_12300) r423 <= _26926;
  wire [1:0] _26927 = {_0, _1599} + {_0, _3390};
  wire [1:0] _26928 = {_0, _4574} + {_0, _6397};
  wire [2:0] _26929 = {_0, _26927} + {_0, _26928};
  wire [1:0] _26930 = {_0, _9022} + {_0, _11004};
  wire [3:0] _26931 = {_0, _26929} + {_0, _0, _26930};
  wire _26932 = _12301 < _26931;
  wire _26933 = r422 ^ _26932;
  wire _26934 = _12298 ? coded_block[422] : r422;
  wire _26935 = _12296 ? _26933 : _26934;
  always @ (posedge reset or posedge clock) if (reset) r422 <= 1'd0; else if (_12300) r422 <= _26935;
  wire [1:0] _26936 = {_0, _1631} + {_0, _3037};
  wire [1:0] _26937 = {_0, _5470} + {_0, _6652};
  wire [2:0] _26938 = {_0, _26936} + {_0, _26937};
  wire [1:0] _26939 = {_0, _8480} + {_0, _11101};
  wire [3:0] _26940 = {_0, _26938} + {_0, _0, _26939};
  wire _26941 = _12301 < _26940;
  wire _26942 = r421 ^ _26941;
  wire _26943 = _12298 ? coded_block[421] : r421;
  wire _26944 = _12296 ? _26942 : _26943;
  always @ (posedge reset or posedge clock) if (reset) r421 <= 1'd0; else if (_12300) r421 <= _26944;
  wire [1:0] _26945 = {_0, _1662} + {_0, _3262};
  wire [1:0] _26946 = {_0, _5116} + {_0, _7548};
  wire [2:0] _26947 = {_0, _26945} + {_0, _26946};
  wire [1:0] _26948 = {_0, _8736} + {_0, _10558};
  wire [3:0] _26949 = {_0, _26947} + {_0, _0, _26948};
  wire _26950 = _12301 < _26949;
  wire _26951 = r420 ^ _26950;
  wire _26952 = _12298 ? coded_block[420] : r420;
  wire _26953 = _12296 ? _26951 : _26952;
  always @ (posedge reset or posedge clock) if (reset) r420 <= 1'd0; else if (_12300) r420 <= _26953;
  wire [1:0] _26954 = {_0, _1695} + {_0, _3135};
  wire [1:0] _26955 = {_0, _5342} + {_0, _7199};
  wire [2:0] _26956 = {_0, _26954} + {_0, _26955};
  wire [1:0] _26957 = {_0, _9630} + {_0, _10814};
  wire [3:0] _26958 = {_0, _26956} + {_0, _0, _26957};
  wire _26959 = _12301 < _26958;
  wire _26960 = r419 ^ _26959;
  wire _26961 = _12298 ? coded_block[419] : r419;
  wire _26962 = _12296 ? _26960 : _26961;
  always @ (posedge reset or posedge clock) if (reset) r419 <= 1'd0; else if (_12300) r419 <= _26962;
  wire [1:0] _26963 = {_0, _1726} + {_0, _3486};
  wire [1:0] _26964 = {_0, _5215} + {_0, _7420};
  wire [2:0] _26965 = {_0, _26963} + {_0, _26964};
  wire [1:0] _26966 = {_0, _9279} + {_0, _11708};
  wire [3:0] _26967 = {_0, _26965} + {_0, _0, _26966};
  wire _26968 = _12301 < _26967;
  wire _26969 = r418 ^ _26968;
  wire _26970 = _12298 ? coded_block[418] : r418;
  wire _26971 = _12296 ? _26969 : _26970;
  always @ (posedge reset or posedge clock) if (reset) r418 <= 1'd0; else if (_12300) r418 <= _26971;
  wire [1:0] _26972 = {_0, _1758} + {_0, _2208};
  wire [1:0] _26973 = {_0, _5565} + {_0, _7293};
  wire [2:0] _26974 = {_0, _26972} + {_0, _26973};
  wire [1:0] _26975 = {_0, _9503} + {_0, _11358};
  wire [3:0] _26976 = {_0, _26974} + {_0, _0, _26975};
  wire _26977 = _12301 < _26976;
  wire _26978 = r417 ^ _26977;
  wire _26979 = _12298 ? coded_block[417] : r417;
  wire _26980 = _12296 ? _26978 : _26979;
  always @ (posedge reset or posedge clock) if (reset) r417 <= 1'd0; else if (_12300) r417 <= _26980;
  wire [1:0] _26981 = {_0, _1789} + {_0, _2813};
  wire [1:0] _26982 = {_0, _4287} + {_0, _7644};
  wire [2:0] _26983 = {_0, _26981} + {_0, _26982};
  wire [1:0] _26984 = {_0, _9375} + {_0, _11581};
  wire [3:0] _26985 = {_0, _26983} + {_0, _0, _26984};
  wire _26986 = _12301 < _26985;
  wire _26987 = r416 ^ _26986;
  wire _26988 = _12298 ? coded_block[416] : r416;
  wire _26989 = _12296 ? _26987 : _26988;
  always @ (posedge reset or posedge clock) if (reset) r416 <= 1'd0; else if (_12300) r416 <= _26989;
  wire [1:0] _26990 = {_0, _1823} + {_0, _2367};
  wire [1:0] _26991 = {_0, _4895} + {_0, _6366};
  wire [2:0] _26992 = {_0, _26990} + {_0, _26991};
  wire [1:0] _26993 = {_0, _9724} + {_0, _11453};
  wire [3:0] _26994 = {_0, _26992} + {_0, _0, _26993};
  wire _26995 = _12301 < _26994;
  wire _26996 = r415 ^ _26995;
  wire _26997 = _12298 ? coded_block[415] : r415;
  wire _26998 = _12296 ? _26996 : _26997;
  always @ (posedge reset or posedge clock) if (reset) r415 <= 1'd0; else if (_12300) r415 <= _26998;
  wire [1:0] _26999 = {_0, _1854} + {_0, _3997};
  wire [1:0] _27000 = {_0, _4447} + {_0, _6973};
  wire [2:0] _27001 = {_0, _26999} + {_0, _27000};
  wire [1:0] _27002 = {_0, _8446} + {_0, _11806};
  wire [3:0] _27003 = {_0, _27001} + {_0, _0, _27002};
  wire _27004 = _12301 < _27003;
  wire _27005 = r414 ^ _27004;
  wire _27006 = _12298 ? coded_block[414] : r414;
  wire _27007 = _12296 ? _27005 : _27006;
  always @ (posedge reset or posedge clock) if (reset) r414 <= 1'd0; else if (_12300) r414 <= _27007;
  wire [1:0] _27008 = {_0, _1886} + {_0, _3005};
  wire [1:0] _27009 = {_0, _6076} + {_0, _6525};
  wire [2:0] _27010 = {_0, _27008} + {_0, _27009};
  wire [1:0] _27011 = {_0, _9054} + {_0, _10527};
  wire [3:0] _27012 = {_0, _27010} + {_0, _0, _27011};
  wire _27013 = _12301 < _27012;
  wire _27014 = r413 ^ _27013;
  wire _27015 = _12298 ? coded_block[413] : r413;
  wire _27016 = _12296 ? _27014 : _27015;
  always @ (posedge reset or posedge clock) if (reset) r413 <= 1'd0; else if (_12300) r413 <= _27016;
  wire [1:0] _27017 = {_0, _1917} + {_0, _3422};
  wire [1:0] _27018 = {_0, _5085} + {_0, _8155};
  wire [2:0] _27019 = {_0, _27017} + {_0, _27018};
  wire [1:0] _27020 = {_0, _8607} + {_0, _11132};
  wire [3:0] _27021 = {_0, _27019} + {_0, _0, _27020};
  wire _27022 = _12301 < _27021;
  wire _27023 = r412 ^ _27022;
  wire _27024 = _12298 ? coded_block[412] : r412;
  wire _27025 = _12296 ? _27023 : _27024;
  always @ (posedge reset or posedge clock) if (reset) r412 <= 1'd0; else if (_12300) r412 <= _27025;
  wire [1:0] _27026 = {_0, _1950} + {_0, _3901};
  wire [1:0] _27027 = {_0, _5501} + {_0, _7163};
  wire [2:0] _27028 = {_0, _27026} + {_0, _27027};
  wire [1:0] _27029 = {_0, _10235} + {_0, _10685};
  wire [3:0] _27030 = {_0, _27028} + {_0, _0, _27029};
  wire _27031 = _12301 < _27030;
  wire _27032 = r411 ^ _27031;
  wire _27033 = _12298 ? coded_block[411] : r411;
  wire _27034 = _12296 ? _27032 : _27033;
  always @ (posedge reset or posedge clock) if (reset) r411 <= 1'd0; else if (_12300) r411 <= _27034;
  wire [1:0] _27035 = {_0, _1981} + {_0, _3325};
  wire [1:0] _27036 = {_0, _5981} + {_0, _7581};
  wire [2:0] _27037 = {_0, _27035} + {_0, _27036};
  wire [1:0] _27038 = {_0, _9248} + {_0, _10303};
  wire [3:0] _27039 = {_0, _27037} + {_0, _0, _27038};
  wire _27040 = _12301 < _27039;
  wire _27041 = r410 ^ _27040;
  wire _27042 = _12298 ? coded_block[410] : r410;
  wire _27043 = _12296 ? _27041 : _27042;
  always @ (posedge reset or posedge clock) if (reset) r410 <= 1'd0; else if (_12300) r410 <= _27043;
  wire [1:0] _27044 = {_0, _2013} + {_0, _2623};
  wire [1:0] _27045 = {_0, _5407} + {_0, _8059};
  wire [2:0] _27046 = {_0, _27044} + {_0, _27045};
  wire [1:0] _27047 = {_0, _9661} + {_0, _11326};
  wire [3:0] _27048 = {_0, _27046} + {_0, _0, _27047};
  wire _27049 = _12301 < _27048;
  wire _27050 = r409 ^ _27049;
  wire _27051 = _12298 ? coded_block[409] : r409;
  wire _27052 = _12296 ? _27050 : _27051;
  always @ (posedge reset or posedge clock) if (reset) r409 <= 1'd0; else if (_12300) r409 <= _27052;
  wire [1:0] _27053 = {_0, _65} + {_0, _2463};
  wire [1:0] _27054 = {_0, _4384} + {_0, _6781};
  wire [2:0] _27055 = {_0, _27053} + {_0, _27054};
  wire [1:0] _27056 = {_0, _9566} + {_0, _12219};
  wire [3:0] _27057 = {_0, _27055} + {_0, _0, _27056};
  wire _27058 = _12301 < _27057;
  wire _27059 = r408 ^ _27058;
  wire _27060 = _12298 ? coded_block[408] : r408;
  wire _27061 = _12296 ? _27059 : _27060;
  always @ (posedge reset or posedge clock) if (reset) r408 <= 1'd0; else if (_12300) r408 <= _27061;
  wire [1:0] _27062 = {_0, _97} + {_0, _2271};
  wire [1:0] _27063 = {_0, _4542} + {_0, _6462};
  wire [2:0] _27064 = {_0, _27062} + {_0, _27063};
  wire [1:0] _27065 = {_0, _8863} + {_0, _11644};
  wire [3:0] _27066 = {_0, _27064} + {_0, _0, _27065};
  wire _27067 = _12301 < _27066;
  wire _27068 = r407 ^ _27067;
  wire _27069 = _12298 ? coded_block[407] : r407;
  wire _27070 = _12296 ? _27068 : _27069;
  always @ (posedge reset or posedge clock) if (reset) r407 <= 1'd0; else if (_12300) r407 <= _27070;
  wire [1:0] _27071 = {_0, _161} + {_0, _3805};
  wire [1:0] _27072 = {_0, _4734} + {_0, _6431};
  wire [2:0] _27073 = {_0, _27071} + {_0, _27072};
  wire [1:0] _27074 = {_0, _8701} + {_0, _10621};
  wire [3:0] _27075 = {_0, _27073} + {_0, _0, _27074};
  wire _27076 = _12301 < _27075;
  wire _27077 = r406 ^ _27076;
  wire _27078 = _12298 ? coded_block[406] : r406;
  wire _27079 = _12296 ? _27077 : _27078;
  always @ (posedge reset or posedge clock) if (reset) r406 <= 1'd0; else if (_12300) r406 <= _27079;
  wire [1:0] _27080 = {_0, _192} + {_0, _3580};
  wire [1:0] _27081 = {_0, _5884} + {_0, _6814};
  wire [2:0] _27082 = {_0, _27080} + {_0, _27081};
  wire [1:0] _27083 = {_0, _8511} + {_0, _10783};
  wire [3:0] _27084 = {_0, _27082} + {_0, _0, _27083};
  wire _27085 = _12301 < _27084;
  wire _27086 = r405 ^ _27085;
  wire _27087 = _12298 ? coded_block[405] : r405;
  wire _27088 = _12296 ? _27086 : _27087;
  always @ (posedge reset or posedge clock) if (reset) r405 <= 1'd0; else if (_12300) r405 <= _27088;
  wire [1:0] _27089 = {_0, _224} + {_0, _2144};
  wire [1:0] _27090 = {_0, _5663} + {_0, _7965};
  wire [2:0] _27091 = {_0, _27089} + {_0, _27090};
  wire [1:0] _27092 = {_0, _8894} + {_0, _10590};
  wire [3:0] _27093 = {_0, _27091} + {_0, _0, _27092};
  wire _27094 = _12301 < _27093;
  wire _27095 = r404 ^ _27094;
  wire _27096 = _12298 ? coded_block[404] : r404;
  wire _27097 = _12296 ? _27095 : _27096;
  always @ (posedge reset or posedge clock) if (reset) r404 <= 1'd0; else if (_12300) r404 <= _27097;
  wire [1:0] _27098 = {_0, _255} + {_0, _4091};
  wire [1:0] _27099 = {_0, _4223} + {_0, _7741};
  wire [2:0] _27100 = {_0, _27098} + {_0, _27099};
  wire [1:0] _27101 = {_0, _10045} + {_0, _10973};
  wire [3:0] _27102 = {_0, _27100} + {_0, _0, _27101};
  wire _27103 = _12301 < _27102;
  wire _27104 = r403 ^ _27103;
  wire _27105 = _12298 ? coded_block[403] : r403;
  wire _27106 = _12296 ? _27104 : _27105;
  always @ (posedge reset or posedge clock) if (reset) r403 <= 1'd0; else if (_12300) r403 <= _27106;
  wire [1:0] _27107 = {_0, _289} + {_0, _3198};
  wire [1:0] _27108 = {_0, _4160} + {_0, _6303};
  wire [2:0] _27109 = {_0, _27107} + {_0, _27108};
  wire [1:0] _27110 = {_0, _9822} + {_0, _12124};
  wire [3:0] _27111 = {_0, _27109} + {_0, _0, _27110};
  wire _27112 = _12301 < _27111;
  wire _27113 = r402 ^ _27112;
  wire _27114 = _12298 ? coded_block[402] : r402;
  wire _27115 = _12296 ? _27113 : _27114;
  always @ (posedge reset or posedge clock) if (reset) r402 <= 1'd0; else if (_12300) r402 <= _27115;
  wire [1:0] _27116 = {_0, _320} + {_0, _3870};
  wire [1:0] _27117 = {_0, _5279} + {_0, _6239};
  wire [2:0] _27118 = {_0, _27116} + {_0, _27117};
  wire [1:0] _27119 = {_0, _8383} + {_0, _11900};
  wire [3:0] _27120 = {_0, _27118} + {_0, _0, _27119};
  wire _27121 = _12301 < _27120;
  wire _27122 = r401 ^ _27121;
  wire _27123 = _12298 ? coded_block[401] : r401;
  wire _27124 = _12296 ? _27122 : _27123;
  always @ (posedge reset or posedge clock) if (reset) r401 <= 1'd0; else if (_12300) r401 <= _27124;
  wire [1:0] _27125 = {_0, _383} + {_0, _3167};
  wire [1:0] _27126 = {_0, _5534} + {_0, _8028};
  wire [2:0] _27127 = {_0, _27125} + {_0, _27126};
  wire [1:0] _27128 = {_0, _9438} + {_0, _10399};
  wire [3:0] _27129 = {_0, _27127} + {_0, _0, _27128};
  wire _27130 = _12301 < _27129;
  wire _27131 = r400 ^ _27130;
  wire _27132 = _12298 ? coded_block[400] : r400;
  wire _27133 = _12296 ? _27131 : _27132;
  always @ (posedge reset or posedge clock) if (reset) r400 <= 1'd0; else if (_12300) r400 <= _27133;
  wire [1:0] _27134 = {_0, _416} + {_0, _2112};
  wire [1:0] _27135 = {_0, _5246} + {_0, _7612};
  wire [2:0] _27136 = {_0, _27134} + {_0, _27135};
  wire [1:0] _27137 = {_0, _10108} + {_0, _11516};
  wire [3:0] _27138 = {_0, _27136} + {_0, _0, _27137};
  wire _27139 = _12301 < _27138;
  wire _27140 = r399 ^ _27139;
  wire _27141 = _12298 ? coded_block[399] : r399;
  wire _27142 = _12296 ? _27140 : _27141;
  always @ (posedge reset or posedge clock) if (reset) r399 <= 1'd0; else if (_12300) r399 <= _27142;
  wire [1:0] _27143 = {_0, _447} + {_0, _3615};
  wire [1:0] _27144 = {_0, _4192} + {_0, _7326};
  wire [2:0] _27145 = {_0, _27143} + {_0, _27144};
  wire [1:0] _27146 = {_0, _9693} + {_0, _12188};
  wire [3:0] _27147 = {_0, _27145} + {_0, _0, _27146};
  wire _27148 = _12301 < _27147;
  wire _27149 = r398 ^ _27148;
  wire _27150 = _12298 ? coded_block[398] : r398;
  wire _27151 = _12296 ? _27149 : _27150;
  always @ (posedge reset or posedge clock) if (reset) r398 <= 1'd0; else if (_12300) r398 <= _27151;
  wire [1:0] _27152 = {_0, _479} + {_0, _2592};
  wire [1:0] _27153 = {_0, _5694} + {_0, _6270};
  wire [2:0] _27154 = {_0, _27152} + {_0, _27153};
  wire [1:0] _27155 = {_0, _9406} + {_0, _11771};
  wire [3:0] _27156 = {_0, _27154} + {_0, _0, _27155};
  wire _27157 = _12301 < _27156;
  wire _27158 = r397 ^ _27157;
  wire _27159 = _12298 ? coded_block[397] : r397;
  wire _27160 = _12296 ? _27158 : _27159;
  always @ (posedge reset or posedge clock) if (reset) r397 <= 1'd0; else if (_12300) r397 <= _27160;
  wire [1:0] _27161 = {_0, _510} + {_0, _3359};
  wire [1:0] _27162 = {_0, _4671} + {_0, _7773};
  wire [2:0] _27163 = {_0, _27161} + {_0, _27162};
  wire [1:0] _27164 = {_0, _8352} + {_0, _11485};
  wire [3:0] _27165 = {_0, _27163} + {_0, _0, _27164};
  wire _27166 = _12301 < _27165;
  wire _27167 = r396 ^ _27166;
  wire _27168 = _12298 ? coded_block[396] : r396;
  wire _27169 = _12296 ? _27167 : _27168;
  always @ (posedge reset or posedge clock) if (reset) r396 <= 1'd0; else if (_12300) r396 <= _27169;
  wire [1:0] _27170 = {_0, _545} + {_0, _2526};
  wire [1:0] _27171 = {_0, _5438} + {_0, _6750};
  wire [2:0] _27172 = {_0, _27170} + {_0, _27171};
  wire [1:0] _27173 = {_0, _9853} + {_0, _10430};
  wire [3:0] _27174 = {_0, _27172} + {_0, _0, _27173};
  wire _27175 = _12301 < _27174;
  wire _27176 = r395 ^ _27175;
  wire _27177 = _12298 ? coded_block[395] : r395;
  wire _27178 = _12296 ? _27176 : _27177;
  always @ (posedge reset or posedge clock) if (reset) r395 <= 1'd0; else if (_12300) r395 <= _27178;
  wire [1:0] _27179 = {_0, _576} + {_0, _4060};
  wire [1:0] _27180 = {_0, _4605} + {_0, _7517};
  wire [2:0] _27181 = {_0, _27179} + {_0, _27180};
  wire [1:0] _27182 = {_0, _8830} + {_0, _11933};
  wire [3:0] _27183 = {_0, _27181} + {_0, _0, _27182};
  wire _27184 = _12301 < _27183;
  wire _27185 = r394 ^ _27184;
  wire _27186 = _12298 ? coded_block[394] : r394;
  wire _27187 = _12296 ? _27185 : _27186;
  always @ (posedge reset or posedge clock) if (reset) r394 <= 1'd0; else if (_12300) r394 <= _27187;
  wire [1:0] _27188 = {_0, _608} + {_0, _2175};
  wire [1:0] _27189 = {_0, _6139} + {_0, _6687};
  wire [2:0] _27190 = {_0, _27188} + {_0, _27189};
  wire [1:0] _27191 = {_0, _9597} + {_0, _10910};
  wire [3:0] _27192 = {_0, _27190} + {_0, _0, _27191};
  wire _27193 = _12301 < _27192;
  wire _27194 = r393 ^ _27193;
  wire _27195 = _12298 ? coded_block[393] : r393;
  wire _27196 = _12296 ? _27194 : _27195;
  always @ (posedge reset or posedge clock) if (reset) r393 <= 1'd0; else if (_12300) r393 <= _27196;
  wire [1:0] _27197 = {_0, _703} + {_0, _2719};
  wire [1:0] _27198 = {_0, _4830} + {_0, _7675};
  wire [2:0] _27199 = {_0, _27197} + {_0, _27198};
  wire [1:0] _27200 = {_0, _8415} + {_0, _10366};
  wire [3:0] _27201 = {_0, _27199} + {_0, _0, _27200};
  wire _27202 = _12301 < _27201;
  wire _27203 = r392 ^ _27202;
  wire _27204 = _12298 ? coded_block[392] : r392;
  wire _27205 = _12296 ? _27203 : _27204;
  always @ (posedge reset or posedge clock) if (reset) r392 <= 1'd0; else if (_12300) r392 <= _27205;
  wire [1:0] _27206 = {_0, _320} + {_0, _2526};
  wire [1:0] _27207 = {_0, _4129} + {_0, _6652};
  wire [2:0] _27208 = {_0, _27206} + {_0, _27207};
  wire [1:0] _27209 = {_0, _8894} + {_0, _11581};
  wire [3:0] _27210 = {_0, _27208} + {_0, _0, _27209};
  wire _27211 = _12301 < _27210;
  wire _27212 = r391 ^ _27211;
  wire _27213 = _12298 ? coded_block[391] : r391;
  wire _27214 = _12296 ? _27212 : _27213;
  always @ (posedge reset or posedge clock) if (reset) r391 <= 1'd0; else if (_12300) r391 <= _27214;
  wire [1:0] _27215 = {_0, _990} + {_0, _3742};
  wire [1:0] _27216 = {_0, _4767} + {_0, _7581};
  wire [2:0] _27217 = {_0, _27215} + {_0, _27216};
  wire [1:0] _27218 = {_0, _8799} + {_0, _10366};
  wire [3:0] _27219 = {_0, _27217} + {_0, _0, _27218};
  wire _27220 = _12301 < _27219;
  wire _27221 = r390 ^ _27220;
  wire _27222 = _12298 ? coded_block[390] : r390;
  wire _27223 = _12296 ? _27221 : _27222;
  always @ (posedge reset or posedge clock) if (reset) r390 <= 1'd0; else if (_12300) r390 <= _27223;
  wire [1:0] _27224 = {_0, _1021} + {_0, _2271};
  wire [1:0] _27225 = {_0, _5821} + {_0, _6845};
  wire [2:0] _27226 = {_0, _27224} + {_0, _27225};
  wire [1:0] _27227 = {_0, _9661} + {_0, _10877};
  wire [3:0] _27228 = {_0, _27226} + {_0, _0, _27227};
  wire _27229 = _12301 < _27228;
  wire _27230 = r389 ^ _27229;
  wire _27231 = _12298 ? coded_block[389] : r389;
  wire _27232 = _12296 ? _27230 : _27231;
  always @ (posedge reset or posedge clock) if (reset) r389 <= 1'd0; else if (_12300) r389 <= _27232;
  wire [1:0] _27233 = {_0, _1057} + {_0, _3359};
  wire [1:0] _27234 = {_0, _4350} + {_0, _7900};
  wire [2:0] _27235 = {_0, _27233} + {_0, _27234};
  wire [1:0] _27236 = {_0, _8926} + {_0, _11740};
  wire [3:0] _27237 = {_0, _27235} + {_0, _0, _27236};
  wire _27238 = _12301 < _27237;
  wire _27239 = r388 ^ _27238;
  wire _27240 = _12298 ? coded_block[388] : r388;
  wire _27241 = _12296 ? _27239 : _27240;
  always @ (posedge reset or posedge clock) if (reset) r388 <= 1'd0; else if (_12300) r388 <= _27241;
  wire [1:0] _27242 = {_0, _1088} + {_0, _3678};
  wire [1:0] _27243 = {_0, _5438} + {_0, _6431};
  wire [2:0] _27244 = {_0, _27242} + {_0, _27243};
  wire [1:0] _27245 = {_0, _9980} + {_0, _11004};
  wire [3:0] _27246 = {_0, _27244} + {_0, _0, _27245};
  wire _27247 = _12301 < _27246;
  wire _27248 = r387 ^ _27247;
  wire _27249 = _12298 ? coded_block[387] : r387;
  wire _27250 = _12296 ? _27248 : _27249;
  always @ (posedge reset or posedge clock) if (reset) r387 <= 1'd0; else if (_12300) r387 <= _27250;
  wire [1:0] _27251 = {_0, _1120} + {_0, _2112};
  wire [1:0] _27252 = {_0, _5757} + {_0, _7517};
  wire [2:0] _27253 = {_0, _27251} + {_0, _27252};
  wire [1:0] _27254 = {_0, _8511} + {_0, _12061};
  wire [3:0] _27255 = {_0, _27253} + {_0, _0, _27254};
  wire _27256 = _12301 < _27255;
  wire _27257 = r386 ^ _27256;
  wire _27258 = _12298 ? coded_block[386] : r386;
  wire _27259 = _12296 ? _27257 : _27258;
  always @ (posedge reset or posedge clock) if (reset) r386 <= 1'd0; else if (_12300) r386 <= _27259;
  wire [1:0] _27260 = {_0, _1151} + {_0, _3486};
  wire [1:0] _27261 = {_0, _4192} + {_0, _7837};
  wire [2:0] _27262 = {_0, _27260} + {_0, _27261};
  wire [1:0] _27263 = {_0, _9597} + {_0, _10590};
  wire [3:0] _27264 = {_0, _27262} + {_0, _0, _27263};
  wire _27265 = _12301 < _27264;
  wire _27266 = r385 ^ _27265;
  wire _27267 = _12298 ? coded_block[385] : r385;
  wire _27268 = _12296 ? _27266 : _27267;
  always @ (posedge reset or posedge clock) if (reset) r385 <= 1'd0; else if (_12300) r385 <= _27268;
  wire [1:0] _27269 = {_0, _1184} + {_0, _2399};
  wire [1:0] _27270 = {_0, _5565} + {_0, _6270};
  wire [2:0] _27271 = {_0, _27269} + {_0, _27270};
  wire [1:0] _27272 = {_0, _9917} + {_0, _11677};
  wire [3:0] _27273 = {_0, _27271} + {_0, _0, _27272};
  wire _27274 = _12301 < _27273;
  wire _27275 = r384 ^ _27274;
  wire _27276 = _12298 ? coded_block[384] : r384;
  wire _27277 = _12296 ? _27275 : _27276;
  always @ (posedge reset or posedge clock) if (reset) r384 <= 1'd0; else if (_12300) r384 <= _27277;
  wire [1:0] _27278 = {_0, _1215} + {_0, _2494};
  wire [1:0] _27279 = {_0, _4478} + {_0, _7644};
  wire [2:0] _27280 = {_0, _27278} + {_0, _27279};
  wire [1:0] _27281 = {_0, _8352} + {_0, _11996};
  wire [3:0] _27282 = {_0, _27280} + {_0, _0, _27281};
  wire _27283 = _12301 < _27282;
  wire _27284 = r383 ^ _27283;
  wire _27285 = _12298 ? coded_block[383] : r383;
  wire _27286 = _12296 ? _27284 : _27285;
  always @ (posedge reset or posedge clock) if (reset) r383 <= 1'd0; else if (_12300) r383 <= _27286;
  wire [1:0] _27287 = {_0, _1247} + {_0, _3964};
  wire [1:0] _27288 = {_0, _4574} + {_0, _6558};
  wire [2:0] _27289 = {_0, _27287} + {_0, _27288};
  wire [1:0] _27290 = {_0, _9724} + {_0, _10430};
  wire [3:0] _27291 = {_0, _27289} + {_0, _0, _27290};
  wire _27292 = _12301 < _27291;
  wire _27293 = r382 ^ _27292;
  wire _27294 = _12298 ? coded_block[382] : r382;
  wire _27295 = _12296 ? _27293 : _27294;
  always @ (posedge reset or posedge clock) if (reset) r382 <= 1'd0; else if (_12300) r382 <= _27295;
  wire [1:0] _27296 = {_0, _1278} + {_0, _2208};
  wire [1:0] _27297 = {_0, _6045} + {_0, _6652};
  wire [2:0] _27298 = {_0, _27296} + {_0, _27297};
  wire [1:0] _27299 = {_0, _8638} + {_0, _11806};
  wire [3:0] _27300 = {_0, _27298} + {_0, _0, _27299};
  wire _27301 = _12301 < _27300;
  wire _27302 = r381 ^ _27301;
  wire _27303 = _12298 ? coded_block[381] : r381;
  wire _27304 = _12296 ? _27302 : _27303;
  always @ (posedge reset or posedge clock) if (reset) r381 <= 1'd0; else if (_12300) r381 <= _27304;
  wire [1:0] _27305 = {_0, _1312} + {_0, _3104};
  wire [1:0] _27306 = {_0, _4287} + {_0, _8123};
  wire [2:0] _27307 = {_0, _27305} + {_0, _27306};
  wire [1:0] _27308 = {_0, _8736} + {_0, _10717};
  wire [3:0] _27309 = {_0, _27307} + {_0, _0, _27308};
  wire _27310 = _12301 < _27309;
  wire _27311 = r380 ^ _27310;
  wire _27312 = _12298 ? coded_block[380] : r380;
  wire _27313 = _12296 ? _27311 : _27312;
  always @ (posedge reset or posedge clock) if (reset) r380 <= 1'd0; else if (_12300) r380 <= _27313;
  wire [1:0] _27314 = {_0, _1343} + {_0, _2750};
  wire [1:0] _27315 = {_0, _5183} + {_0, _6366};
  wire [2:0] _27316 = {_0, _27314} + {_0, _27315};
  wire [1:0] _27317 = {_0, _10204} + {_0, _10814};
  wire [3:0] _27318 = {_0, _27316} + {_0, _0, _27317};
  wire _27319 = _12301 < _27318;
  wire _27320 = r379 ^ _27319;
  wire _27321 = _12298 ? coded_block[379] : r379;
  wire _27322 = _12296 ? _27320 : _27321;
  always @ (posedge reset or posedge clock) if (reset) r379 <= 1'd0; else if (_12300) r379 <= _27322;
  wire [1:0] _27323 = {_0, _1375} + {_0, _2974};
  wire [1:0] _27324 = {_0, _4830} + {_0, _7262};
  wire [2:0] _27325 = {_0, _27323} + {_0, _27324};
  wire [1:0] _27326 = {_0, _8446} + {_0, _12282};
  wire [3:0] _27327 = {_0, _27325} + {_0, _0, _27326};
  wire _27328 = _12301 < _27327;
  wire _27329 = r378 ^ _27328;
  wire _27330 = _12298 ? coded_block[378] : r378;
  wire _27331 = _12296 ? _27329 : _27330;
  always @ (posedge reset or posedge clock) if (reset) r378 <= 1'd0; else if (_12300) r378 <= _27331;
  wire [1:0] _27332 = {_0, _1406} + {_0, _2847};
  wire [1:0] _27333 = {_0, _5053} + {_0, _6908};
  wire [2:0] _27334 = {_0, _27332} + {_0, _27333};
  wire [1:0] _27335 = {_0, _9342} + {_0, _10527};
  wire [3:0] _27336 = {_0, _27334} + {_0, _0, _27335};
  wire _27337 = _12301 < _27336;
  wire _27338 = r377 ^ _27337;
  wire _27339 = _12298 ? coded_block[377] : r377;
  wire _27340 = _12296 ? _27338 : _27339;
  always @ (posedge reset or posedge clock) if (reset) r377 <= 1'd0; else if (_12300) r377 <= _27340;
  wire [1:0] _27341 = {_0, _1439} + {_0, _3198};
  wire [1:0] _27342 = {_0, _4926} + {_0, _7132};
  wire [2:0] _27343 = {_0, _27341} + {_0, _27342};
  wire [1:0] _27344 = {_0, _8991} + {_0, _11422};
  wire [3:0] _27345 = {_0, _27343} + {_0, _0, _27344};
  wire _27346 = _12301 < _27345;
  wire _27347 = r376 ^ _27346;
  wire _27348 = _12298 ? coded_block[376] : r376;
  wire _27349 = _12296 ? _27347 : _27348;
  always @ (posedge reset or posedge clock) if (reset) r376 <= 1'd0; else if (_12300) r376 <= _27349;
  wire [1:0] _27350 = {_0, _1470} + {_0, _3933};
  wire [1:0] _27351 = {_0, _5279} + {_0, _7005};
  wire [2:0] _27352 = {_0, _27350} + {_0, _27351};
  wire [1:0] _27353 = {_0, _9212} + {_0, _11069};
  wire [3:0] _27354 = {_0, _27352} + {_0, _0, _27353};
  wire _27355 = _12301 < _27354;
  wire _27356 = r375 ^ _27355;
  wire _27357 = _12298 ? coded_block[375] : r375;
  wire _27358 = _12296 ? _27356 : _27357;
  always @ (posedge reset or posedge clock) if (reset) r375 <= 1'd0; else if (_12300) r375 <= _27358;
  wire [1:0] _27359 = {_0, _1502} + {_0, _2526};
  wire [1:0] _27360 = {_0, _6012} + {_0, _7357};
  wire [2:0] _27361 = {_0, _27359} + {_0, _27360};
  wire [1:0] _27362 = {_0, _9085} + {_0, _11295};
  wire [3:0] _27363 = {_0, _27361} + {_0, _0, _27362};
  wire _27364 = _12301 < _27363;
  wire _27365 = r374 ^ _27364;
  wire _27366 = _12298 ? coded_block[374] : r374;
  wire _27367 = _12296 ? _27365 : _27366;
  always @ (posedge reset or posedge clock) if (reset) r374 <= 1'd0; else if (_12300) r374 <= _27367;
  wire [1:0] _27368 = {_0, _1533} + {_0, _4091};
  wire [1:0] _27369 = {_0, _4605} + {_0, _8092};
  wire [2:0] _27370 = {_0, _27368} + {_0, _27369};
  wire [1:0] _27371 = {_0, _9438} + {_0, _11165};
  wire [3:0] _27372 = {_0, _27370} + {_0, _0, _27371};
  wire _27373 = _12301 < _27372;
  wire _27374 = r373 ^ _27373;
  wire _27375 = _12298 ? coded_block[373] : r373;
  wire _27376 = _12296 ? _27374 : _27375;
  always @ (posedge reset or posedge clock) if (reset) r373 <= 1'd0; else if (_12300) r373 <= _27376;
  wire [1:0] _27377 = {_0, _1568} + {_0, _3709};
  wire [1:0] _27378 = {_0, _4160} + {_0, _6687};
  wire [2:0] _27379 = {_0, _27377} + {_0, _27378};
  wire [1:0] _27380 = {_0, _10172} + {_0, _11516};
  wire [3:0] _27381 = {_0, _27379} + {_0, _0, _27380};
  wire _27382 = _12301 < _27381;
  wire _27383 = r372 ^ _27382;
  wire _27384 = _12298 ? coded_block[372] : r372;
  wire _27385 = _12296 ? _27383 : _27384;
  always @ (posedge reset or posedge clock) if (reset) r372 <= 1'd0; else if (_12300) r372 <= _27385;
  wire [1:0] _27386 = {_0, _1599} + {_0, _2719};
  wire [1:0] _27387 = {_0, _5790} + {_0, _6239};
  wire [2:0] _27388 = {_0, _27386} + {_0, _27387};
  wire [1:0] _27389 = {_0, _8767} + {_0, _12251};
  wire [3:0] _27390 = {_0, _27388} + {_0, _0, _27389};
  wire _27391 = _12301 < _27390;
  wire _27392 = r371 ^ _27391;
  wire _27393 = _12298 ? coded_block[371] : r371;
  wire _27394 = _12296 ? _27392 : _27393;
  always @ (posedge reset or posedge clock) if (reset) r371 <= 1'd0; else if (_12300) r371 <= _27394;
  wire [1:0] _27395 = {_0, _1631} + {_0, _3135};
  wire [1:0] _27396 = {_0, _4798} + {_0, _7868};
  wire [2:0] _27397 = {_0, _27395} + {_0, _27396};
  wire [1:0] _27398 = {_0, _8319} + {_0, _10846};
  wire [3:0] _27399 = {_0, _27397} + {_0, _0, _27398};
  wire _27400 = _12301 < _27399;
  wire _27401 = r370 ^ _27400;
  wire _27402 = _12298 ? coded_block[370] : r370;
  wire _27403 = _12296 ? _27401 : _27402;
  always @ (posedge reset or posedge clock) if (reset) r370 <= 1'd0; else if (_12300) r370 <= _27403;
  wire [1:0] _27404 = {_0, _1662} + {_0, _3615};
  wire [1:0] _27405 = {_0, _5215} + {_0, _6877};
  wire [2:0] _27406 = {_0, _27404} + {_0, _27405};
  wire [1:0] _27407 = {_0, _9949} + {_0, _10399};
  wire [3:0] _27408 = {_0, _27406} + {_0, _0, _27407};
  wire _27409 = _12301 < _27408;
  wire _27410 = r369 ^ _27409;
  wire _27411 = _12298 ? coded_block[369] : r369;
  wire _27412 = _12296 ? _27410 : _27411;
  always @ (posedge reset or posedge clock) if (reset) r369 <= 1'd0; else if (_12300) r369 <= _27412;
  wire [1:0] _27413 = {_0, _1695} + {_0, _3037};
  wire [1:0] _27414 = {_0, _5694} + {_0, _7293};
  wire [2:0] _27415 = {_0, _27413} + {_0, _27414};
  wire [1:0] _27416 = {_0, _8957} + {_0, _12027};
  wire [3:0] _27417 = {_0, _27415} + {_0, _0, _27416};
  wire _27418 = _12301 < _27417;
  wire _27419 = r368 ^ _27418;
  wire _27420 = _12298 ? coded_block[368] : r368;
  wire _27421 = _12296 ? _27419 : _27420;
  always @ (posedge reset or posedge clock) if (reset) r368 <= 1'd0; else if (_12300) r368 <= _27421;
  wire [1:0] _27422 = {_0, _1726} + {_0, _2336};
  wire [1:0] _27423 = {_0, _5116} + {_0, _7773};
  wire [2:0] _27424 = {_0, _27422} + {_0, _27423};
  wire [1:0] _27425 = {_0, _9375} + {_0, _11038};
  wire [3:0] _27426 = {_0, _27424} + {_0, _0, _27425};
  wire _27427 = _12301 < _27426;
  wire _27428 = r367 ^ _27427;
  wire _27429 = _12298 ? coded_block[367] : r367;
  wire _27430 = _12296 ? _27428 : _27429;
  always @ (posedge reset or posedge clock) if (reset) r367 <= 1'd0; else if (_12300) r367 <= _27430;
  wire [1:0] _27431 = {_0, _1758} + {_0, _4028};
  wire [1:0] _27432 = {_0, _4415} + {_0, _7199};
  wire [2:0] _27433 = {_0, _27431} + {_0, _27432};
  wire [1:0] _27434 = {_0, _9853} + {_0, _11453};
  wire [3:0] _27435 = {_0, _27433} + {_0, _0, _27434};
  wire _27436 = _12301 < _27435;
  wire _27437 = r366 ^ _27436;
  wire _27438 = _12298 ? coded_block[366] : r366;
  wire _27439 = _12296 ? _27437 : _27438;
  always @ (posedge reset or posedge clock) if (reset) r366 <= 1'd0; else if (_12300) r366 <= _27439;
  wire [1:0] _27440 = {_0, _1789} + {_0, _2175};
  wire [1:0] _27441 = {_0, _6108} + {_0, _6494};
  wire [2:0] _27442 = {_0, _27440} + {_0, _27441};
  wire [1:0] _27443 = {_0, _9279} + {_0, _11933};
  wire [3:0] _27444 = {_0, _27442} + {_0, _0, _27443};
  wire _27445 = _12301 < _27444;
  wire _27446 = r365 ^ _27445;
  wire _27447 = _12298 ? coded_block[365] : r365;
  wire _27448 = _12296 ? _27446 : _27447;
  always @ (posedge reset or posedge clock) if (reset) r365 <= 1'd0; else if (_12300) r365 <= _27448;
  wire [1:0] _27449 = {_0, _1823} + {_0, _3997};
  wire [1:0] _27450 = {_0, _4256} + {_0, _8186};
  wire [2:0] _27451 = {_0, _27449} + {_0, _27450};
  wire [1:0] _27452 = {_0, _8574} + {_0, _11358};
  wire [3:0] _27453 = {_0, _27451} + {_0, _0, _27452};
  wire _27454 = _12301 < _27453;
  wire _27455 = r364 ^ _27454;
  wire _27456 = _12298 ? coded_block[364] : r364;
  wire _27457 = _12296 ? _27455 : _27456;
  always @ (posedge reset or posedge clock) if (reset) r364 <= 1'd0; else if (_12300) r364 <= _27457;
  wire [1:0] _27458 = {_0, _1854} + {_0, _2367};
  wire [1:0] _27459 = {_0, _6076} + {_0, _6334};
  wire [2:0] _27460 = {_0, _27458} + {_0, _27459};
  wire [1:0] _27461 = {_0, _8256} + {_0, _10654};
  wire [3:0] _27462 = {_0, _27460} + {_0, _0, _27461};
  wire _27463 = _12301 < _27462;
  wire _27464 = r363 ^ _27463;
  wire _27465 = _12298 ? coded_block[363] : r363;
  wire _27466 = _12296 ? _27464 : _27465;
  always @ (posedge reset or posedge clock) if (reset) r363 <= 1'd0; else if (_12300) r363 <= _27466;
  wire [1:0] _27467 = {_0, _1886} + {_0, _3517};
  wire [1:0] _27468 = {_0, _4447} + {_0, _8155};
  wire [2:0] _27469 = {_0, _27467} + {_0, _27468};
  wire [1:0] _27470 = {_0, _8415} + {_0, _10335};
  wire [3:0] _27471 = {_0, _27469} + {_0, _0, _27470};
  wire _27472 = _12301 < _27471;
  wire _27473 = r362 ^ _27472;
  wire _27474 = _12298 ? coded_block[362] : r362;
  wire _27475 = _12296 ? _27473 : _27474;
  always @ (posedge reset or posedge clock) if (reset) r362 <= 1'd0; else if (_12300) r362 <= _27475;
  wire [1:0] _27476 = {_0, _1917} + {_0, _3294};
  wire [1:0] _27477 = {_0, _5597} + {_0, _6525};
  wire [2:0] _27478 = {_0, _27476} + {_0, _27477};
  wire [1:0] _27479 = {_0, _10235} + {_0, _10493};
  wire [3:0] _27480 = {_0, _27478} + {_0, _0, _27479};
  wire _27481 = _12301 < _27480;
  wire _27482 = r361 ^ _27481;
  wire _27483 = _12298 ? coded_block[361] : r361;
  wire _27484 = _12296 ? _27482 : _27483;
  always @ (posedge reset or posedge clock) if (reset) r361 <= 1'd0; else if (_12300) r361 <= _27484;
  wire [1:0] _27485 = {_0, _1950} + {_0, _3870};
  wire [1:0] _27486 = {_0, _5373} + {_0, _7675};
  wire [2:0] _27487 = {_0, _27485} + {_0, _27486};
  wire [1:0] _27488 = {_0, _8607} + {_0, _10303};
  wire [3:0] _27489 = {_0, _27487} + {_0, _0, _27488};
  wire _27490 = _12301 < _27489;
  wire _27491 = r360 ^ _27490;
  wire _27492 = _12298 ? coded_block[360] : r360;
  wire _27493 = _12296 ? _27491 : _27492;
  always @ (posedge reset or posedge clock) if (reset) r360 <= 1'd0; else if (_12300) r360 <= _27493;
  wire [1:0] _27494 = {_0, _1981} + {_0, _3805};
  wire [1:0] _27495 = {_0, _5949} + {_0, _7454};
  wire [2:0] _27496 = {_0, _27494} + {_0, _27495};
  wire [1:0] _27497 = {_0, _9759} + {_0, _10685};
  wire [3:0] _27498 = {_0, _27496} + {_0, _0, _27497};
  wire _27499 = _12301 < _27498;
  wire _27500 = r359 ^ _27499;
  wire _27501 = _12298 ? coded_block[359] : r359;
  wire _27502 = _12296 ? _27500 : _27501;
  always @ (posedge reset or posedge clock) if (reset) r359 <= 1'd0; else if (_12300) r359 <= _27502;
  wire [1:0] _27503 = {_0, _2013} + {_0, _2910};
  wire [1:0] _27504 = {_0, _5884} + {_0, _8028};
  wire [2:0] _27505 = {_0, _27503} + {_0, _27504};
  wire [1:0] _27506 = {_0, _9534} + {_0, _11837};
  wire [3:0] _27507 = {_0, _27505} + {_0, _0, _27506};
  wire _27508 = _12301 < _27507;
  wire _27509 = r358 ^ _27508;
  wire _27510 = _12298 ? coded_block[358] : r358;
  wire _27511 = _12296 ? _27509 : _27510;
  always @ (posedge reset or posedge clock) if (reset) r358 <= 1'd0; else if (_12300) r358 <= _27511;
  wire [1:0] _27512 = {_0, _2044} + {_0, _3580};
  wire [1:0] _27513 = {_0, _4989} + {_0, _7965};
  wire [2:0] _27514 = {_0, _27512} + {_0, _27513};
  wire [1:0] _27515 = {_0, _10108} + {_0, _11613};
  wire [3:0] _27516 = {_0, _27514} + {_0, _0, _27515};
  wire _27517 = _12301 < _27516;
  wire _27518 = r357 ^ _27517;
  wire _27519 = _12298 ? coded_block[357] : r357;
  wire _27520 = _12296 ? _27518 : _27519;
  always @ (posedge reset or posedge clock) if (reset) r357 <= 1'd0; else if (_12300) r357 <= _27520;
  wire [1:0] _27521 = {_0, _65} + {_0, _3167};
  wire [1:0] _27522 = {_0, _5663} + {_0, _7069};
  wire [2:0] _27523 = {_0, _27521} + {_0, _27522};
  wire [1:0] _27524 = {_0, _10045} + {_0, _12188};
  wire [3:0] _27525 = {_0, _27523} + {_0, _0, _27524};
  wire _27526 = _12301 < _27525;
  wire _27527 = r356 ^ _27526;
  wire _27528 = _12298 ? coded_block[356] : r356;
  wire _27529 = _12296 ? _27527 : _27528;
  always @ (posedge reset or posedge clock) if (reset) r356 <= 1'd0; else if (_12300) r356 <= _27529;
  wire [1:0] _27530 = {_0, _97} + {_0, _2878};
  wire [1:0] _27531 = {_0, _5246} + {_0, _7741};
  wire [2:0] _27532 = {_0, _27530} + {_0, _27531};
  wire [1:0] _27533 = {_0, _9149} + {_0, _12124};
  wire [3:0] _27534 = {_0, _27532} + {_0, _0, _27533};
  wire _27535 = _12301 < _27534;
  wire _27536 = r355 ^ _27535;
  wire _27537 = _12298 ? coded_block[355] : r355;
  wire _27538 = _12296 ? _27536 : _27537;
  always @ (posedge reset or posedge clock) if (reset) r355 <= 1'd0; else if (_12300) r355 <= _27538;
  wire [1:0] _27539 = {_0, _161} + {_0, _3325};
  wire [1:0] _27540 = {_0, _5918} + {_0, _7036};
  wire [2:0] _27541 = {_0, _27539} + {_0, _27540};
  wire [1:0] _27542 = {_0, _9406} + {_0, _11900};
  wire [3:0] _27543 = {_0, _27541} + {_0, _0, _27542};
  wire _27544 = _12301 < _27543;
  wire _27545 = r354 ^ _27544;
  wire _27546 = _12298 ? coded_block[354] : r354;
  wire _27547 = _12296 ? _27545 : _27546;
  always @ (posedge reset or posedge clock) if (reset) r354 <= 1'd0; else if (_12300) r354 <= _27547;
  wire [1:0] _27548 = {_0, _192} + {_0, _2302};
  wire [1:0] _27549 = {_0, _5407} + {_0, _7996};
  wire [2:0] _27550 = {_0, _27548} + {_0, _27549};
  wire [1:0] _27551 = {_0, _9118} + {_0, _11485};
  wire [3:0] _27552 = {_0, _27550} + {_0, _0, _27551};
  wire _27553 = _12301 < _27552;
  wire _27554 = r353 ^ _27553;
  wire _27555 = _12298 ? coded_block[353] : r353;
  wire _27556 = _12296 ? _27554 : _27555;
  always @ (posedge reset or posedge clock) if (reset) r353 <= 1'd0; else if (_12300) r353 <= _27556;
  wire [1:0] _27557 = {_0, _224} + {_0, _3068};
  wire [1:0] _27558 = {_0, _4384} + {_0, _7485};
  wire [2:0] _27559 = {_0, _27557} + {_0, _27558};
  wire [1:0] _27560 = {_0, _10077} + {_0, _11196};
  wire [3:0] _27561 = {_0, _27559} + {_0, _0, _27560};
  wire _27562 = _12301 < _27561;
  wire _27563 = r352 ^ _27562;
  wire _27564 = _12298 ? coded_block[352] : r352;
  wire _27565 = _12296 ? _27563 : _27564;
  always @ (posedge reset or posedge clock) if (reset) r352 <= 1'd0; else if (_12300) r352 <= _27565;
  wire [1:0] _27566 = {_0, _255} + {_0, _2239};
  wire [1:0] _27567 = {_0, _5152} + {_0, _6462};
  wire [2:0] _27568 = {_0, _27566} + {_0, _27567};
  wire [1:0] _27569 = {_0, _9566} + {_0, _12155};
  wire [3:0] _27570 = {_0, _27568} + {_0, _0, _27569};
  wire _27571 = _12301 < _27570;
  wire _27572 = r351 ^ _27571;
  wire _27573 = _12298 ? coded_block[351] : r351;
  wire _27574 = _12296 ? _27572 : _27573;
  always @ (posedge reset or posedge clock) if (reset) r351 <= 1'd0; else if (_12300) r351 <= _27574;
  wire [1:0] _27575 = {_0, _320} + {_0, _3901};
  wire [1:0] _27576 = {_0, _5853} + {_0, _6397};
  wire [2:0] _27577 = {_0, _27575} + {_0, _27576};
  wire [1:0] _27578 = {_0, _9311} + {_0, _10621};
  wire [3:0] _27579 = {_0, _27577} + {_0, _0, _27578};
  wire _27580 = _12301 < _27579;
  wire _27581 = r350 ^ _27580;
  wire _27582 = _12298 ? coded_block[350] : r350;
  wire _27583 = _12296 ? _27581 : _27582;
  always @ (posedge reset or posedge clock) if (reset) r350 <= 1'd0; else if (_12300) r350 <= _27583;
  wire [1:0] _27584 = {_0, _352} + {_0, _3231};
  wire [1:0] _27585 = {_0, _5981} + {_0, _7931};
  wire [2:0] _27586 = {_0, _27584} + {_0, _27585};
  wire [1:0] _27587 = {_0, _8480} + {_0, _11389};
  wire [3:0] _27588 = {_0, _27586} + {_0, _0, _27587};
  wire _27589 = _12301 < _27588;
  wire _27590 = r349 ^ _27589;
  wire _27591 = _12298 ? coded_block[349] : r349;
  wire _27592 = _12296 ? _27590 : _27591;
  always @ (posedge reset or posedge clock) if (reset) r349 <= 1'd0; else if (_12300) r349 <= _27592;
  wire [1:0] _27593 = {_0, _383} + {_0, _2463};
  wire [1:0] _27594 = {_0, _5310} + {_0, _8059};
  wire [2:0] _27595 = {_0, _27593} + {_0, _27594};
  wire [1:0] _27596 = {_0, _10014} + {_0, _10558};
  wire [3:0] _27597 = {_0, _27595} + {_0, _0, _27596};
  wire _27598 = _12301 < _27597;
  wire _27599 = r348 ^ _27598;
  wire _27600 = _12298 ? coded_block[348] : r348;
  wire _27601 = _12296 ? _27599 : _27600;
  always @ (posedge reset or posedge clock) if (reset) r348 <= 1'd0; else if (_12300) r348 <= _27601;
  wire [1:0] _27602 = {_0, _416} + {_0, _2430};
  wire [1:0] _27603 = {_0, _4542} + {_0, _7389};
  wire [2:0] _27604 = {_0, _27602} + {_0, _27603};
  wire [1:0] _27605 = {_0, _10141} + {_0, _12092};
  wire [3:0] _27606 = {_0, _27604} + {_0, _0, _27605};
  wire _27607 = _12301 < _27606;
  wire _27608 = r347 ^ _27607;
  wire _27609 = _12298 ? coded_block[347] : r347;
  wire _27610 = _12296 ? _27608 : _27609;
  always @ (posedge reset or posedge clock) if (reset) r347 <= 1'd0; else if (_12300) r347 <= _27610;
  wire [1:0] _27611 = {_0, _447} + {_0, _3262};
  wire [1:0] _27612 = {_0, _4511} + {_0, _6621};
  wire [2:0] _27613 = {_0, _27611} + {_0, _27612};
  wire [1:0] _27614 = {_0, _9469} + {_0, _12219};
  wire [3:0] _27615 = {_0, _27613} + {_0, _0, _27614};
  wire _27616 = _12301 < _27615;
  wire _27617 = r346 ^ _27616;
  wire _27618 = _12298 ? coded_block[346] : r346;
  wire _27619 = _12296 ? _27617 : _27618;
  always @ (posedge reset or posedge clock) if (reset) r346 <= 1'd0; else if (_12300) r346 <= _27619;
  wire [1:0] _27620 = {_0, _479} + {_0, _3549};
  wire [1:0] _27621 = {_0, _5342} + {_0, _6589};
  wire [2:0] _27622 = {_0, _27620} + {_0, _27621};
  wire [1:0] _27623 = {_0, _8701} + {_0, _11550};
  wire [3:0] _27624 = {_0, _27622} + {_0, _0, _27623};
  wire _27625 = _12301 < _27624;
  wire _27626 = r345 ^ _27625;
  wire _27627 = _12298 ? coded_block[345] : r345;
  wire _27628 = _12296 ? _27626 : _27627;
  always @ (posedge reset or posedge clock) if (reset) r345 <= 1'd0; else if (_12300) r345 <= _27628;
  wire [1:0] _27629 = {_0, _510} + {_0, _2941};
  wire [1:0] _27630 = {_0, _5628} + {_0, _7420};
  wire [2:0] _27631 = {_0, _27629} + {_0, _27630};
  wire [1:0] _27632 = {_0, _8670} + {_0, _10783};
  wire [3:0] _27633 = {_0, _27631} + {_0, _0, _27632};
  wire _27634 = _12301 < _27633;
  wire _27635 = r344 ^ _27634;
  wire _27636 = _12298 ? coded_block[344] : r344;
  wire _27637 = _12296 ? _27635 : _27636;
  always @ (posedge reset or posedge clock) if (reset) r344 <= 1'd0; else if (_12300) r344 <= _27637;
  wire [1:0] _27638 = {_0, _545} + {_0, _2782};
  wire [1:0] _27639 = {_0, _5022} + {_0, _7710};
  wire [2:0] _27640 = {_0, _27638} + {_0, _27639};
  wire [1:0] _27641 = {_0, _9503} + {_0, _10748};
  wire [3:0] _27642 = {_0, _27640} + {_0, _0, _27641};
  wire _27643 = _12301 < _27642;
  wire _27644 = r343 ^ _27643;
  wire _27645 = _12298 ? coded_block[343] : r343;
  wire _27646 = _12296 ? _27644 : _27645;
  always @ (posedge reset or posedge clock) if (reset) r343 <= 1'd0; else if (_12300) r343 <= _27646;
  wire [1:0] _27647 = {_0, _576} + {_0, _2081};
  wire [1:0] _27648 = {_0, _4861} + {_0, _7100};
  wire [2:0] _27649 = {_0, _27647} + {_0, _27648};
  wire [1:0] _27650 = {_0, _9790} + {_0, _11581};
  wire [3:0] _27651 = {_0, _27649} + {_0, _0, _27650};
  wire _27652 = _12301 < _27651;
  wire _27653 = r342 ^ _27652;
  wire _27654 = _12298 ? coded_block[342] : r342;
  wire _27655 = _12296 ? _27653 : _27654;
  always @ (posedge reset or posedge clock) if (reset) r342 <= 1'd0; else if (_12300) r342 <= _27655;
  wire [1:0] _27656 = {_0, _608} + {_0, _2813};
  wire [1:0] _27657 = {_0, _4129} + {_0, _6942};
  wire [2:0] _27658 = {_0, _27656} + {_0, _27657};
  wire [1:0] _27659 = {_0, _9181} + {_0, _11869};
  wire [3:0] _27660 = {_0, _27658} + {_0, _0, _27659};
  wire _27661 = _12301 < _27660;
  wire _27662 = r341 ^ _27661;
  wire _27663 = _12298 ? coded_block[341] : r341;
  wire _27664 = _12296 ? _27662 : _27663;
  always @ (posedge reset or posedge clock) if (reset) r341 <= 1'd0; else if (_12300) r341 <= _27664;
  wire [1:0] _27665 = {_0, _639} + {_0, _3005};
  wire [1:0] _27666 = {_0, _4895} + {_0, _6176};
  wire [2:0] _27667 = {_0, _27665} + {_0, _27666};
  wire [1:0] _27668 = {_0, _9022} + {_0, _11259};
  wire [3:0] _27669 = {_0, _27667} + {_0, _0, _27668};
  wire _27670 = _12301 < _27669;
  wire _27671 = r340 ^ _27670;
  wire _27672 = _12298 ? coded_block[340] : r340;
  wire _27673 = _12296 ? _27671 : _27672;
  always @ (posedge reset or posedge clock) if (reset) r340 <= 1'd0; else if (_12300) r340 <= _27673;
  wire [1:0] _27674 = {_0, _672} + {_0, _3646};
  wire [1:0] _27675 = {_0, _5085} + {_0, _6973};
  wire [2:0] _27676 = {_0, _27674} + {_0, _27675};
  wire [1:0] _27677 = {_0, _8225} + {_0, _11101};
  wire [3:0] _27678 = {_0, _27676} + {_0, _0, _27677};
  wire _27679 = _12301 < _27678;
  wire _27680 = r339 ^ _27679;
  wire _27681 = _12298 ? coded_block[339] : r339;
  wire _27682 = _12296 ? _27680 : _27681;
  always @ (posedge reset or posedge clock) if (reset) r339 <= 1'd0; else if (_12300) r339 <= _27682;
  wire [1:0] _27683 = {_0, _703} + {_0, _3390};
  wire [1:0] _27684 = {_0, _5726} + {_0, _7163};
  wire [2:0] _27685 = {_0, _27683} + {_0, _27684};
  wire [1:0] _27686 = {_0, _9054} + {_0, _10272};
  wire [3:0] _27687 = {_0, _27685} + {_0, _0, _27686};
  wire _27688 = _12301 < _27687;
  wire _27689 = r338 ^ _27688;
  wire _27690 = _12298 ? coded_block[338] : r338;
  wire _27691 = _12296 ? _27689 : _27690;
  always @ (posedge reset or posedge clock) if (reset) r338 <= 1'd0; else if (_12300) r338 <= _27691;
  wire [1:0] _27692 = {_0, _735} + {_0, _2592};
  wire [1:0] _27693 = {_0, _5470} + {_0, _7804};
  wire [2:0] _27694 = {_0, _27692} + {_0, _27693};
  wire [1:0] _27695 = {_0, _9248} + {_0, _11132};
  wire [3:0] _27696 = {_0, _27694} + {_0, _0, _27695};
  wire _27697 = _12301 < _27696;
  wire _27698 = r337 ^ _27697;
  wire _27699 = _12298 ? coded_block[337] : r337;
  wire _27700 = _12296 ? _27698 : _27699;
  always @ (posedge reset or posedge clock) if (reset) r337 <= 1'd0; else if (_12300) r337 <= _27700;
  wire [1:0] _27701 = {_0, _766} + {_0, _2655};
  wire [1:0] _27702 = {_0, _4671} + {_0, _7548};
  wire [2:0] _27703 = {_0, _27701} + {_0, _27702};
  wire [1:0] _27704 = {_0, _9886} + {_0, _11326};
  wire [3:0] _27705 = {_0, _27703} + {_0, _0, _27704};
  wire _27706 = _12301 < _27705;
  wire _27707 = r336 ^ _27706;
  wire _27708 = _12298 ? coded_block[336] : r336;
  wire _27709 = _12296 ? _27707 : _27708;
  always @ (posedge reset or posedge clock) if (reset) r336 <= 1'd0; else if (_12300) r336 <= _27709;
  wire [1:0] _27710 = {_0, _800} + {_0, _3453};
  wire [1:0] _27711 = {_0, _4734} + {_0, _6750};
  wire [2:0] _27712 = {_0, _27710} + {_0, _27711};
  wire [1:0] _27713 = {_0, _9630} + {_0, _11964};
  wire [3:0] _27714 = {_0, _27712} + {_0, _0, _27713};
  wire _27715 = _12301 < _27714;
  wire _27716 = r335 ^ _27715;
  wire _27717 = _12298 ? coded_block[335] : r335;
  wire _27718 = _12296 ? _27716 : _27717;
  always @ (posedge reset or posedge clock) if (reset) r335 <= 1'd0; else if (_12300) r335 <= _27718;
  wire [1:0] _27719 = {_0, _863} + {_0, _4060};
  wire [1:0] _27720 = {_0, _4223} + {_0, _7612};
  wire [2:0] _27721 = {_0, _27719} + {_0, _27720};
  wire [1:0] _27722 = {_0, _8894} + {_0, _10910};
  wire [3:0] _27723 = {_0, _27721} + {_0, _0, _27722};
  wire _27724 = _12301 < _27723;
  wire _27725 = r334 ^ _27724;
  wire _27726 = _12298 ? coded_block[334] : r334;
  wire _27727 = _12296 ? _27725 : _27726;
  always @ (posedge reset or posedge clock) if (reset) r334 <= 1'd0; else if (_12300) r334 <= _27727;
  wire [1:0] _27728 = {_0, _927} + {_0, _3422};
  wire [1:0] _27729 = {_0, _4640} + {_0, _6207};
  wire [2:0] _27730 = {_0, _27728} + {_0, _27729};
  wire [1:0] _27731 = {_0, _8383} + {_0, _11771};
  wire [3:0] _27732 = {_0, _27730} + {_0, _0, _27731};
  wire _27733 = _12301 < _27732;
  wire _27734 = r333 ^ _27733;
  wire _27735 = _12298 ? coded_block[333] : r333;
  wire _27736 = _12296 ? _27734 : _27735;
  always @ (posedge reset or posedge clock) if (reset) r333 <= 1'd0; else if (_12300) r333 <= _27736;
  wire [1:0] _27737 = {_0, _34} + {_0, _2463};
  wire [1:0] _27738 = {_0, _4542} + {_0, _6621};
  wire [2:0] _27739 = {_0, _27737} + {_0, _27738};
  wire [1:0] _27740 = {_0, _8701} + {_0, _10783};
  wire [3:0] _27741 = {_0, _27739} + {_0, _0, _27740};
  wire _27742 = _12301 < _27741;
  wire _27743 = r332 ^ _27742;
  wire _27744 = _12298 ? coded_block[332] : r332;
  wire _27745 = _12296 ? _27743 : _27744;
  always @ (posedge reset or posedge clock) if (reset) r332 <= 1'd0; else if (_12300) r332 <= _27745;
  wire [1:0] _27746 = {_0, _1215} + {_0, _2813};
  wire [1:0] _27747 = {_0, _4671} + {_0, _7100};
  wire [2:0] _27748 = {_0, _27746} + {_0, _27747};
  wire [1:0] _27749 = {_0, _8288} + {_0, _12124};
  wire [3:0] _27750 = {_0, _27748} + {_0, _0, _27749};
  wire _27751 = _12301 < _27750;
  wire _27752 = r331 ^ _27751;
  wire _27753 = _12298 ? coded_block[331] : r331;
  wire _27754 = _12296 ? _27752 : _27753;
  always @ (posedge reset or posedge clock) if (reset) r331 <= 1'd0; else if (_12300) r331 <= _27754;
  wire [1:0] _27755 = {_0, _1247} + {_0, _2686};
  wire [1:0] _27756 = {_0, _4895} + {_0, _6750};
  wire [2:0] _27757 = {_0, _27755} + {_0, _27756};
  wire [1:0] _27758 = {_0, _9181} + {_0, _10366};
  wire [3:0] _27759 = {_0, _27757} + {_0, _0, _27758};
  wire _27760 = _12301 < _27759;
  wire _27761 = r330 ^ _27760;
  wire _27762 = _12298 ? coded_block[330] : r330;
  wire _27763 = _12296 ? _27761 : _27762;
  always @ (posedge reset or posedge clock) if (reset) r330 <= 1'd0; else if (_12300) r330 <= _27763;
  wire [1:0] _27764 = {_0, _1278} + {_0, _3037};
  wire [1:0] _27765 = {_0, _4767} + {_0, _6973};
  wire [2:0] _27766 = {_0, _27764} + {_0, _27765};
  wire [1:0] _27767 = {_0, _8830} + {_0, _11259};
  wire [3:0] _27768 = {_0, _27766} + {_0, _0, _27767};
  wire _27769 = _12301 < _27768;
  wire _27770 = r329 ^ _27769;
  wire _27771 = _12298 ? coded_block[329] : r329;
  wire _27772 = _12296 ? _27770 : _27771;
  always @ (posedge reset or posedge clock) if (reset) r329 <= 1'd0; else if (_12300) r329 <= _27772;
  wire [1:0] _27773 = {_0, _1343} + {_0, _2367};
  wire [1:0] _27774 = {_0, _5853} + {_0, _7199};
  wire [2:0] _27775 = {_0, _27773} + {_0, _27774};
  wire [1:0] _27776 = {_0, _8926} + {_0, _11132};
  wire [3:0] _27777 = {_0, _27775} + {_0, _0, _27776};
  wire _27778 = _12301 < _27777;
  wire _27779 = r328 ^ _27778;
  wire _27780 = _12298 ? coded_block[328] : r328;
  wire _27781 = _12296 ? _27779 : _27780;
  always @ (posedge reset or posedge clock) if (reset) r328 <= 1'd0; else if (_12300) r328 <= _27781;
  wire [1:0] _27782 = {_0, _1375} + {_0, _3933};
  wire [1:0] _27783 = {_0, _4447} + {_0, _7931};
  wire [2:0] _27784 = {_0, _27782} + {_0, _27783};
  wire [1:0] _27785 = {_0, _9279} + {_0, _11004};
  wire [3:0] _27786 = {_0, _27784} + {_0, _0, _27785};
  wire _27787 = _12301 < _27786;
  wire _27788 = r327 ^ _27787;
  wire _27789 = _12298 ? coded_block[327] : r327;
  wire _27790 = _12296 ? _27788 : _27789;
  always @ (posedge reset or posedge clock) if (reset) r327 <= 1'd0; else if (_12300) r327 <= _27790;
  wire [1:0] _27791 = {_0, _1406} + {_0, _3549};
  wire [1:0] _27792 = {_0, _6012} + {_0, _6525};
  wire [2:0] _27793 = {_0, _27791} + {_0, _27792};
  wire [1:0] _27794 = {_0, _10014} + {_0, _11358};
  wire [3:0] _27795 = {_0, _27793} + {_0, _0, _27794};
  wire _27796 = _12301 < _27795;
  wire _27797 = r326 ^ _27796;
  wire _27798 = _12298 ? coded_block[326] : r326;
  wire _27799 = _12296 ? _27797 : _27798;
  always @ (posedge reset or posedge clock) if (reset) r326 <= 1'd0; else if (_12300) r326 <= _27799;
  wire [1:0] _27800 = {_0, _1439} + {_0, _2557};
  wire [1:0] _27801 = {_0, _5628} + {_0, _8092};
  wire [2:0] _27802 = {_0, _27800} + {_0, _27801};
  wire [1:0] _27803 = {_0, _8607} + {_0, _12092};
  wire [3:0] _27804 = {_0, _27802} + {_0, _0, _27803};
  wire _27805 = _12301 < _27804;
  wire _27806 = r325 ^ _27805;
  wire _27807 = _12298 ? coded_block[325] : r325;
  wire _27808 = _12296 ? _27806 : _27807;
  always @ (posedge reset or posedge clock) if (reset) r325 <= 1'd0; else if (_12300) r325 <= _27808;
  wire [1:0] _27809 = {_0, _1470} + {_0, _2974};
  wire [1:0] _27810 = {_0, _4640} + {_0, _7710};
  wire [2:0] _27811 = {_0, _27809} + {_0, _27810};
  wire [1:0] _27812 = {_0, _10172} + {_0, _10685};
  wire [3:0] _27813 = {_0, _27811} + {_0, _0, _27812};
  wire _27814 = _12301 < _27813;
  wire _27815 = r324 ^ _27814;
  wire _27816 = _12298 ? coded_block[324] : r324;
  wire _27817 = _12296 ? _27815 : _27816;
  always @ (posedge reset or posedge clock) if (reset) r324 <= 1'd0; else if (_12300) r324 <= _27817;
  wire [1:0] _27818 = {_0, _1502} + {_0, _3453};
  wire [1:0] _27819 = {_0, _5053} + {_0, _6718};
  wire [2:0] _27820 = {_0, _27818} + {_0, _27819};
  wire [1:0] _27821 = {_0, _9790} + {_0, _12251};
  wire [3:0] _27822 = {_0, _27820} + {_0, _0, _27821};
  wire _27823 = _12301 < _27822;
  wire _27824 = r323 ^ _27823;
  wire _27825 = _12298 ? coded_block[323] : r323;
  wire _27826 = _12296 ? _27824 : _27825;
  always @ (posedge reset or posedge clock) if (reset) r323 <= 1'd0; else if (_12300) r323 <= _27826;
  wire [1:0] _27827 = {_0, _1568} + {_0, _2175};
  wire [1:0] _27828 = {_0, _4958} + {_0, _7612};
  wire [2:0] _27829 = {_0, _27827} + {_0, _27828};
  wire [1:0] _27830 = {_0, _9212} + {_0, _10877};
  wire [3:0] _27831 = {_0, _27829} + {_0, _0, _27830};
  wire _27832 = _12301 < _27831;
  wire _27833 = r322 ^ _27832;
  wire _27834 = _12298 ? coded_block[322] : r322;
  wire _27835 = _12296 ? _27833 : _27834;
  always @ (posedge reset or posedge clock) if (reset) r322 <= 1'd0; else if (_12300) r322 <= _27835;
  wire [1:0] _27836 = {_0, _1599} + {_0, _3870};
  wire [1:0] _27837 = {_0, _4256} + {_0, _7036};
  wire [2:0] _27838 = {_0, _27836} + {_0, _27837};
  wire [1:0] _27839 = {_0, _9693} + {_0, _11295};
  wire [3:0] _27840 = {_0, _27838} + {_0, _0, _27839};
  wire _27841 = _12301 < _27840;
  wire _27842 = r321 ^ _27841;
  wire _27843 = _12298 ? coded_block[321] : r321;
  wire _27844 = _12296 ? _27842 : _27843;
  always @ (posedge reset or posedge clock) if (reset) r321 <= 1'd0; else if (_12300) r321 <= _27844;
  wire [1:0] _27845 = {_0, _1631} + {_0, _4028};
  wire [1:0] _27846 = {_0, _5949} + {_0, _6334};
  wire [2:0] _27847 = {_0, _27845} + {_0, _27846};
  wire [1:0] _27848 = {_0, _9118} + {_0, _11771};
  wire [3:0] _27849 = {_0, _27847} + {_0, _0, _27848};
  wire _27850 = _12301 < _27849;
  wire _27851 = r320 ^ _27850;
  wire _27852 = _12298 ? coded_block[320] : r320;
  wire _27853 = _12296 ? _27851 : _27852;
  always @ (posedge reset or posedge clock) if (reset) r320 <= 1'd0; else if (_12300) r320 <= _27853;
  wire [1:0] _27854 = {_0, _1662} + {_0, _3836};
  wire [1:0] _27855 = {_0, _6108} + {_0, _8028};
  wire [2:0] _27856 = {_0, _27854} + {_0, _27855};
  wire [1:0] _27857 = {_0, _8415} + {_0, _11196};
  wire [3:0] _27858 = {_0, _27856} + {_0, _0, _27857};
  wire _27859 = _12301 < _27858;
  wire _27860 = r319 ^ _27859;
  wire _27861 = _12298 ? coded_block[319] : r319;
  wire _27862 = _12296 ? _27860 : _27861;
  always @ (posedge reset or posedge clock) if (reset) r319 <= 1'd0; else if (_12300) r319 <= _27862;
  wire [1:0] _27863 = {_0, _1695} + {_0, _2208};
  wire [1:0] _27864 = {_0, _5918} + {_0, _8186};
  wire [2:0] _27865 = {_0, _27863} + {_0, _27864};
  wire [1:0] _27866 = {_0, _10108} + {_0, _10493};
  wire [3:0] _27867 = {_0, _27865} + {_0, _0, _27866};
  wire _27868 = _12301 < _27867;
  wire _27869 = r318 ^ _27868;
  wire _27870 = _12298 ? coded_block[318] : r318;
  wire _27871 = _12296 ? _27869 : _27870;
  always @ (posedge reset or posedge clock) if (reset) r318 <= 1'd0; else if (_12300) r318 <= _27871;
  wire [1:0] _27872 = {_0, _1726} + {_0, _3359};
  wire [1:0] _27873 = {_0, _4287} + {_0, _7996};
  wire [2:0] _27874 = {_0, _27872} + {_0, _27873};
  wire [1:0] _27875 = {_0, _8256} + {_0, _12188};
  wire [3:0] _27876 = {_0, _27874} + {_0, _0, _27875};
  wire _27877 = _12301 < _27876;
  wire _27878 = r317 ^ _27877;
  wire _27879 = _12298 ? coded_block[317] : r317;
  wire _27880 = _12296 ? _27878 : _27879;
  always @ (posedge reset or posedge clock) if (reset) r317 <= 1'd0; else if (_12300) r317 <= _27880;
  wire [1:0] _27881 = {_0, _1758} + {_0, _3135};
  wire [1:0] _27882 = {_0, _5438} + {_0, _6366};
  wire [2:0] _27883 = {_0, _27881} + {_0, _27882};
  wire [1:0] _27884 = {_0, _10077} + {_0, _10335};
  wire [3:0] _27885 = {_0, _27883} + {_0, _0, _27884};
  wire _27886 = _12301 < _27885;
  wire _27887 = r316 ^ _27886;
  wire _27888 = _12298 ? coded_block[316] : r316;
  wire _27889 = _12296 ? _27887 : _27888;
  always @ (posedge reset or posedge clock) if (reset) r316 <= 1'd0; else if (_12300) r316 <= _27889;
  wire [1:0] _27890 = {_0, _1789} + {_0, _3709};
  wire [1:0] _27891 = {_0, _5215} + {_0, _7517};
  wire [2:0] _27892 = {_0, _27890} + {_0, _27891};
  wire [1:0] _27893 = {_0, _8446} + {_0, _12155};
  wire [3:0] _27894 = {_0, _27892} + {_0, _0, _27893};
  wire _27895 = _12301 < _27894;
  wire _27896 = r315 ^ _27895;
  wire _27897 = _12298 ? coded_block[315] : r315;
  wire _27898 = _12296 ? _27896 : _27897;
  always @ (posedge reset or posedge clock) if (reset) r315 <= 1'd0; else if (_12300) r315 <= _27898;
  wire [1:0] _27899 = {_0, _1823} + {_0, _3646};
  wire [1:0] _27900 = {_0, _5790} + {_0, _7293};
  wire [2:0] _27901 = {_0, _27899} + {_0, _27900};
  wire [1:0] _27902 = {_0, _9597} + {_0, _10527};
  wire [3:0] _27903 = {_0, _27901} + {_0, _0, _27902};
  wire _27904 = _12301 < _27903;
  wire _27905 = r314 ^ _27904;
  wire _27906 = _12298 ? coded_block[314] : r314;
  wire _27907 = _12296 ? _27905 : _27906;
  always @ (posedge reset or posedge clock) if (reset) r314 <= 1'd0; else if (_12300) r314 <= _27907;
  wire [1:0] _27908 = {_0, _1854} + {_0, _2750};
  wire [1:0] _27909 = {_0, _5726} + {_0, _7868};
  wire [2:0] _27910 = {_0, _27908} + {_0, _27909};
  wire [1:0] _27911 = {_0, _9375} + {_0, _11677};
  wire [3:0] _27912 = {_0, _27910} + {_0, _0, _27911};
  wire _27913 = _12301 < _27912;
  wire _27914 = r313 ^ _27913;
  wire _27915 = _12298 ? coded_block[313] : r313;
  wire _27916 = _12296 ? _27914 : _27915;
  always @ (posedge reset or posedge clock) if (reset) r313 <= 1'd0; else if (_12300) r313 <= _27916;
  wire [1:0] _27917 = {_0, _1886} + {_0, _3422};
  wire [1:0] _27918 = {_0, _4830} + {_0, _7804};
  wire [2:0] _27919 = {_0, _27917} + {_0, _27918};
  wire [1:0] _27920 = {_0, _9949} + {_0, _11453};
  wire [3:0] _27921 = {_0, _27919} + {_0, _0, _27920};
  wire _27922 = _12301 < _27921;
  wire _27923 = r312 ^ _27922;
  wire _27924 = _12298 ? coded_block[312] : r312;
  wire _27925 = _12296 ? _27923 : _27924;
  always @ (posedge reset or posedge clock) if (reset) r312 <= 1'd0; else if (_12300) r312 <= _27925;
  wire [1:0] _27926 = {_0, _1917} + {_0, _3005};
  wire [1:0] _27927 = {_0, _5501} + {_0, _6908};
  wire [2:0] _27928 = {_0, _27926} + {_0, _27927};
  wire [1:0] _27929 = {_0, _9886} + {_0, _12027};
  wire [3:0] _27930 = {_0, _27928} + {_0, _0, _27929};
  wire _27931 = _12301 < _27930;
  wire _27932 = r311 ^ _27931;
  wire _27933 = _12298 ? coded_block[311] : r311;
  wire _27934 = _12296 ? _27932 : _27933;
  always @ (posedge reset or posedge clock) if (reset) r311 <= 1'd0; else if (_12300) r311 <= _27934;
  wire [1:0] _27935 = {_0, _1950} + {_0, _2719};
  wire [1:0] _27936 = {_0, _5085} + {_0, _7581};
  wire [2:0] _27937 = {_0, _27935} + {_0, _27936};
  wire [1:0] _27938 = {_0, _8991} + {_0, _11964};
  wire [3:0] _27939 = {_0, _27937} + {_0, _0, _27938};
  wire _27940 = _12301 < _27939;
  wire _27941 = r310 ^ _27940;
  wire _27942 = _12298 ? coded_block[310] : r310;
  wire _27943 = _12296 ? _27941 : _27942;
  always @ (posedge reset or posedge clock) if (reset) r310 <= 1'd0; else if (_12300) r310 <= _27943;
  wire [1:0] _27944 = {_0, _1981} + {_0, _3678};
  wire [1:0] _27945 = {_0, _4798} + {_0, _7163};
  wire [2:0] _27946 = {_0, _27944} + {_0, _27945};
  wire [1:0] _27947 = {_0, _9661} + {_0, _11069};
  wire [3:0] _27948 = {_0, _27946} + {_0, _0, _27947};
  wire _27949 = _12301 < _27948;
  wire _27950 = r309 ^ _27949;
  wire _27951 = _12298 ? coded_block[309] : r309;
  wire _27952 = _12296 ? _27950 : _27951;
  always @ (posedge reset or posedge clock) if (reset) r309 <= 1'd0; else if (_12300) r309 <= _27952;
  wire [1:0] _27953 = {_0, _2013} + {_0, _3167};
  wire [1:0] _27954 = {_0, _5757} + {_0, _6877};
  wire [2:0] _27955 = {_0, _27953} + {_0, _27954};
  wire [1:0] _27956 = {_0, _9248} + {_0, _11740};
  wire [3:0] _27957 = {_0, _27955} + {_0, _0, _27956};
  wire _27958 = _12301 < _27957;
  wire _27959 = r308 ^ _27958;
  wire _27960 = _12298 ? coded_block[308] : r308;
  wire _27961 = _12296 ? _27959 : _27960;
  always @ (posedge reset or posedge clock) if (reset) r308 <= 1'd0; else if (_12300) r308 <= _27961;
  wire [1:0] _27962 = {_0, _65} + {_0, _2910};
  wire [1:0] _27963 = {_0, _4223} + {_0, _7326};
  wire [2:0] _27964 = {_0, _27962} + {_0, _27963};
  wire [1:0] _27965 = {_0, _9917} + {_0, _11038};
  wire [3:0] _27966 = {_0, _27964} + {_0, _0, _27965};
  wire _27967 = _12301 < _27966;
  wire _27968 = r307 ^ _27967;
  wire _27969 = _12298 ? coded_block[307] : r307;
  wire _27970 = _12296 ? _27968 : _27969;
  always @ (posedge reset or posedge clock) if (reset) r307 <= 1'd0; else if (_12300) r307 <= _27970;
  wire [1:0] _27971 = {_0, _97} + {_0, _4091};
  wire [1:0] _27972 = {_0, _4989} + {_0, _6303};
  wire [2:0] _27973 = {_0, _27971} + {_0, _27972};
  wire [1:0] _27974 = {_0, _9406} + {_0, _11996};
  wire [3:0] _27975 = {_0, _27973} + {_0, _0, _27974};
  wire _27976 = _12301 < _27975;
  wire _27977 = r306 ^ _27976;
  wire _27978 = _12298 ? coded_block[306] : r306;
  wire _27979 = _12296 ? _27977 : _27978;
  always @ (posedge reset or posedge clock) if (reset) r306 <= 1'd0; else if (_12300) r306 <= _27979;
  wire [1:0] _27980 = {_0, _128} + {_0, _3615};
  wire [1:0] _27981 = {_0, _4160} + {_0, _7069};
  wire [2:0] _27982 = {_0, _27980} + {_0, _27981};
  wire [1:0] _27983 = {_0, _8383} + {_0, _11485};
  wire [3:0] _27984 = {_0, _27982} + {_0, _0, _27983};
  wire _27985 = _12301 < _27984;
  wire _27986 = r305 ^ _27985;
  wire _27987 = _12298 ? coded_block[305] : r305;
  wire _27988 = _12296 ? _27986 : _27987;
  always @ (posedge reset or posedge clock) if (reset) r305 <= 1'd0; else if (_12300) r305 <= _27988;
  wire [1:0] _27989 = {_0, _161} + {_0, _3742};
  wire [1:0] _27990 = {_0, _5694} + {_0, _6239};
  wire [2:0] _27991 = {_0, _27989} + {_0, _27990};
  wire [1:0] _27992 = {_0, _9149} + {_0, _10462};
  wire [3:0] _27993 = {_0, _27991} + {_0, _0, _27992};
  wire _27994 = _12301 < _27993;
  wire _27995 = r304 ^ _27994;
  wire _27996 = _12298 ? coded_block[304] : r304;
  wire _27997 = _12296 ? _27995 : _27996;
  always @ (posedge reset or posedge clock) if (reset) r304 <= 1'd0; else if (_12300) r304 <= _27997;
  wire [1:0] _27998 = {_0, _192} + {_0, _3068};
  wire [1:0] _27999 = {_0, _5821} + {_0, _7773};
  wire [2:0] _28000 = {_0, _27998} + {_0, _27999};
  wire [1:0] _28001 = {_0, _8319} + {_0, _11228};
  wire [3:0] _28002 = {_0, _28000} + {_0, _0, _28001};
  wire _28003 = _12301 < _28002;
  wire _28004 = r303 ^ _28003;
  wire _28005 = _12298 ? coded_block[303] : r303;
  wire _28006 = _12296 ? _28004 : _28005;
  always @ (posedge reset or posedge clock) if (reset) r303 <= 1'd0; else if (_12300) r303 <= _28006;
  wire [1:0] _28007 = {_0, _224} + {_0, _2302};
  wire [1:0] _28008 = {_0, _5152} + {_0, _7900};
  wire [2:0] _28009 = {_0, _28007} + {_0, _28008};
  wire [1:0] _28010 = {_0, _9853} + {_0, _10399};
  wire [3:0] _28011 = {_0, _28009} + {_0, _0, _28010};
  wire _28012 = _12301 < _28011;
  wire _28013 = r302 ^ _28012;
  wire _28014 = _12298 ? coded_block[302] : r302;
  wire _28015 = _12296 ? _28013 : _28014;
  always @ (posedge reset or posedge clock) if (reset) r302 <= 1'd0; else if (_12300) r302 <= _28015;
  wire [1:0] _28016 = {_0, _255} + {_0, _2271};
  wire [1:0] _28017 = {_0, _4384} + {_0, _7230};
  wire [2:0] _28018 = {_0, _28016} + {_0, _28017};
  wire [1:0] _28019 = {_0, _9980} + {_0, _11933};
  wire [3:0] _28020 = {_0, _28018} + {_0, _0, _28019};
  wire _28021 = _12301 < _28020;
  wire _28022 = r301 ^ _28021;
  wire _28023 = _12298 ? coded_block[301] : r301;
  wire _28024 = _12296 ? _28022 : _28023;
  always @ (posedge reset or posedge clock) if (reset) r301 <= 1'd0; else if (_12300) r301 <= _28024;
  wire [1:0] _28025 = {_0, _320} + {_0, _3390};
  wire [1:0] _28026 = {_0, _5183} + {_0, _6431};
  wire [2:0] _28027 = {_0, _28025} + {_0, _28026};
  wire [1:0] _28028 = {_0, _8543} + {_0, _11389};
  wire [3:0] _28029 = {_0, _28027} + {_0, _0, _28028};
  wire _28030 = _12301 < _28029;
  wire _28031 = r300 ^ _28030;
  wire _28032 = _12298 ? coded_block[300] : r300;
  wire _28033 = _12296 ? _28031 : _28032;
  always @ (posedge reset or posedge clock) if (reset) r300 <= 1'd0; else if (_12300) r300 <= _28033;
  wire [1:0] _28034 = {_0, _416} + {_0, _2081};
  wire [1:0] _28035 = {_0, _4703} + {_0, _6942};
  wire [2:0] _28036 = {_0, _28034} + {_0, _28035};
  wire [1:0] _28037 = {_0, _9630} + {_0, _11422};
  wire [3:0] _28038 = {_0, _28036} + {_0, _0, _28037};
  wire _28039 = _12301 < _28038;
  wire _28040 = r299 ^ _28039;
  wire _28041 = _12298 ? coded_block[299] : r299;
  wire _28042 = _12296 ? _28040 : _28041;
  always @ (posedge reset or posedge clock) if (reset) r299 <= 1'd0; else if (_12300) r299 <= _28042;
  wire [1:0] _28043 = {_0, _447} + {_0, _2655};
  wire [1:0] _28044 = {_0, _4129} + {_0, _6781};
  wire [2:0] _28045 = {_0, _28043} + {_0, _28044};
  wire [1:0] _28046 = {_0, _9022} + {_0, _11708};
  wire [3:0] _28047 = {_0, _28045} + {_0, _0, _28046};
  wire _28048 = _12301 < _28047;
  wire _28049 = r298 ^ _28048;
  wire _28050 = _12298 ? coded_block[298] : r298;
  wire _28051 = _12296 ? _28049 : _28050;
  always @ (posedge reset or posedge clock) if (reset) r298 <= 1'd0; else if (_12300) r298 <= _28051;
  wire [1:0] _28052 = {_0, _479} + {_0, _2847};
  wire [1:0] _28053 = {_0, _4734} + {_0, _6176};
  wire [2:0] _28054 = {_0, _28052} + {_0, _28053};
  wire [1:0] _28055 = {_0, _8863} + {_0, _11101};
  wire [3:0] _28056 = {_0, _28054} + {_0, _0, _28055};
  wire _28057 = _12301 < _28056;
  wire _28058 = r297 ^ _28057;
  wire _28059 = _12298 ? coded_block[297] : r297;
  wire _28060 = _12296 ? _28058 : _28059;
  always @ (posedge reset or posedge clock) if (reset) r297 <= 1'd0; else if (_12300) r297 <= _28060;
  wire [1:0] _28061 = {_0, _510} + {_0, _3486};
  wire [1:0] _28062 = {_0, _4926} + {_0, _6814};
  wire [2:0] _28063 = {_0, _28061} + {_0, _28062};
  wire [1:0] _28064 = {_0, _8225} + {_0, _10941};
  wire [3:0] _28065 = {_0, _28063} + {_0, _0, _28064};
  wire _28066 = _12301 < _28065;
  wire _28067 = r296 ^ _28066;
  wire _28068 = _12298 ? coded_block[296] : r296;
  wire _28069 = _12296 ? _28067 : _28068;
  always @ (posedge reset or posedge clock) if (reset) r296 <= 1'd0; else if (_12300) r296 <= _28069;
  wire [1:0] _28070 = {_0, _545} + {_0, _3231};
  wire [1:0] _28071 = {_0, _5565} + {_0, _7005};
  wire [2:0] _28072 = {_0, _28070} + {_0, _28071};
  wire [1:0] _28073 = {_0, _8894} + {_0, _10272};
  wire [3:0] _28074 = {_0, _28072} + {_0, _0, _28073};
  wire _28075 = _12301 < _28074;
  wire _28076 = r295 ^ _28075;
  wire _28077 = _12298 ? coded_block[295] : r295;
  wire _28078 = _12296 ? _28076 : _28077;
  always @ (posedge reset or posedge clock) if (reset) r295 <= 1'd0; else if (_12300) r295 <= _28078;
  wire [1:0] _28079 = {_0, _576} + {_0, _2430};
  wire [1:0] _28080 = {_0, _5310} + {_0, _7644};
  wire [2:0] _28081 = {_0, _28079} + {_0, _28080};
  wire [1:0] _28082 = {_0, _9085} + {_0, _10973};
  wire [3:0] _28083 = {_0, _28081} + {_0, _0, _28082};
  wire _28084 = _12301 < _28083;
  wire _28085 = r294 ^ _28084;
  wire _28086 = _12298 ? coded_block[294] : r294;
  wire _28087 = _12296 ? _28085 : _28086;
  always @ (posedge reset or posedge clock) if (reset) r294 <= 1'd0; else if (_12300) r294 <= _28087;
  wire [1:0] _28088 = {_0, _608} + {_0, _2494};
  wire [1:0] _28089 = {_0, _4511} + {_0, _7389};
  wire [2:0] _28090 = {_0, _28088} + {_0, _28089};
  wire [1:0] _28091 = {_0, _9724} + {_0, _11165};
  wire [3:0] _28092 = {_0, _28090} + {_0, _0, _28091};
  wire _28093 = _12301 < _28092;
  wire _28094 = r293 ^ _28093;
  wire _28095 = _12298 ? coded_block[293] : r293;
  wire _28096 = _12296 ? _28094 : _28095;
  always @ (posedge reset or posedge clock) if (reset) r293 <= 1'd0; else if (_12300) r293 <= _28096;
  wire [1:0] _28097 = {_0, _672} + {_0, _3997};
  wire [1:0] _28098 = {_0, _5373} + {_0, _6652};
  wire [2:0] _28099 = {_0, _28097} + {_0, _28098};
  wire [1:0] _28100 = {_0, _8670} + {_0, _11550};
  wire [3:0] _28101 = {_0, _28099} + {_0, _0, _28100};
  wire _28102 = _12301 < _28101;
  wire _28103 = r292 ^ _28102;
  wire _28104 = _12298 ? coded_block[292] : r292;
  wire _28105 = _12296 ? _28103 : _28104;
  always @ (posedge reset or posedge clock) if (reset) r292 <= 1'd0; else if (_12300) r292 <= _28105;
  wire [1:0] _28106 = {_0, _703} + {_0, _3901};
  wire [1:0] _28107 = {_0, _6076} + {_0, _7454};
  wire [2:0] _28108 = {_0, _28106} + {_0, _28107};
  wire [1:0] _28109 = {_0, _8736} + {_0, _10748};
  wire [3:0] _28110 = {_0, _28108} + {_0, _0, _28109};
  wire _28111 = _12301 < _28110;
  wire _28112 = r291 ^ _28111;
  wire _28113 = _12298 ? coded_block[291] : r291;
  wire _28114 = _12296 ? _28112 : _28113;
  always @ (posedge reset or posedge clock) if (reset) r291 <= 1'd0; else if (_12300) r291 <= _28114;
  wire [1:0] _28115 = {_0, _735} + {_0, _2399};
  wire [1:0] _28116 = {_0, _5981} + {_0, _8155};
  wire [2:0] _28117 = {_0, _28115} + {_0, _28116};
  wire [1:0] _28118 = {_0, _9534} + {_0, _10814};
  wire [3:0] _28119 = {_0, _28117} + {_0, _0, _28118};
  wire _28120 = _12301 < _28119;
  wire _28121 = r290 ^ _28120;
  wire _28122 = _12298 ? coded_block[290] : r290;
  wire _28123 = _12296 ? _28121 : _28122;
  always @ (posedge reset or posedge clock) if (reset) r290 <= 1'd0; else if (_12300) r290 <= _28123;
  wire [1:0] _28124 = {_0, _766} + {_0, _3262};
  wire [1:0] _28125 = {_0, _4478} + {_0, _8059};
  wire [2:0] _28126 = {_0, _28124} + {_0, _28125};
  wire [1:0] _28127 = {_0, _10235} + {_0, _11613};
  wire [3:0] _28128 = {_0, _28126} + {_0, _0, _28127};
  wire _28129 = _12301 < _28128;
  wire _28130 = r289 ^ _28129;
  wire _28131 = _12298 ? coded_block[289] : r289;
  wire _28132 = _12296 ? _28130 : _28131;
  always @ (posedge reset or posedge clock) if (reset) r289 <= 1'd0; else if (_12300) r289 <= _28132;
  wire [1:0] _28133 = {_0, _800} + {_0, _2526};
  wire [1:0] _28134 = {_0, _5342} + {_0, _6558};
  wire [2:0] _28135 = {_0, _28133} + {_0, _28134};
  wire [1:0] _28136 = {_0, _10141} + {_0, _10303};
  wire [3:0] _28137 = {_0, _28135} + {_0, _0, _28136};
  wire _28138 = _12301 < _28137;
  wire _28139 = r288 ^ _28138;
  wire _28140 = _12298 ? coded_block[288] : r288;
  wire _28141 = _12296 ? _28139 : _28140;
  always @ (posedge reset or posedge clock) if (reset) r288 <= 1'd0; else if (_12300) r288 <= _28141;
  wire [1:0] _28142 = {_0, _831} + {_0, _3580};
  wire [1:0] _28143 = {_0, _4605} + {_0, _7420};
  wire [2:0] _28144 = {_0, _28142} + {_0, _28143};
  wire [1:0] _28145 = {_0, _8638} + {_0, _12219};
  wire [3:0] _28146 = {_0, _28144} + {_0, _0, _28145};
  wire _28147 = _12301 < _28146;
  wire _28148 = r287 ^ _28147;
  wire _28149 = _12298 ? coded_block[287] : r287;
  wire _28150 = _12296 ? _28148 : _28149;
  always @ (posedge reset or posedge clock) if (reset) r287 <= 1'd0; else if (_12300) r287 <= _28150;
  wire [1:0] _28151 = {_0, _863} + {_0, _2112};
  wire [1:0] _28152 = {_0, _5663} + {_0, _6687};
  wire [2:0] _28153 = {_0, _28151} + {_0, _28152};
  wire [1:0] _28154 = {_0, _9503} + {_0, _10717};
  wire [3:0] _28155 = {_0, _28153} + {_0, _0, _28154};
  wire _28156 = _12301 < _28155;
  wire _28157 = r286 ^ _28156;
  wire _28158 = _12298 ? coded_block[286] : r286;
  wire _28159 = _12296 ? _28157 : _28158;
  always @ (posedge reset or posedge clock) if (reset) r286 <= 1'd0; else if (_12300) r286 <= _28159;
  wire [1:0] _28160 = {_0, _894} + {_0, _3198};
  wire [1:0] _28161 = {_0, _4192} + {_0, _7741};
  wire [2:0] _28162 = {_0, _28160} + {_0, _28161};
  wire [1:0] _28163 = {_0, _8767} + {_0, _11581};
  wire [3:0] _28164 = {_0, _28162} + {_0, _0, _28163};
  wire _28165 = _12301 < _28164;
  wire _28166 = r285 ^ _28165;
  wire _28167 = _12298 ? coded_block[285] : r285;
  wire _28168 = _12296 ? _28166 : _28167;
  always @ (posedge reset or posedge clock) if (reset) r285 <= 1'd0; else if (_12300) r285 <= _28168;
  wire [1:0] _28169 = {_0, _990} + {_0, _3325};
  wire [1:0] _28170 = {_0, _6045} + {_0, _7675};
  wire [2:0] _28171 = {_0, _28169} + {_0, _28170};
  wire [1:0] _28172 = {_0, _9438} + {_0, _10430};
  wire [3:0] _28173 = {_0, _28171} + {_0, _0, _28172};
  wire _28174 = _12301 < _28173;
  wire _28175 = r284 ^ _28174;
  wire _28176 = _12298 ? coded_block[284] : r284;
  wire _28177 = _12296 ? _28175 : _28176;
  always @ (posedge reset or posedge clock) if (reset) r284 <= 1'd0; else if (_12300) r284 <= _28177;
  wire [1:0] _28178 = {_0, _1021} + {_0, _2239};
  wire [1:0] _28179 = {_0, _5407} + {_0, _8123};
  wire [2:0] _28180 = {_0, _28178} + {_0, _28179};
  wire [1:0] _28181 = {_0, _9759} + {_0, _11516};
  wire [3:0] _28182 = {_0, _28180} + {_0, _0, _28181};
  wire _28183 = _12301 < _28182;
  wire _28184 = r283 ^ _28183;
  wire _28185 = _12298 ? coded_block[283] : r283;
  wire _28186 = _12296 ? _28184 : _28185;
  always @ (posedge reset or posedge clock) if (reset) r283 <= 1'd0; else if (_12300) r283 <= _28186;
  wire [1:0] _28187 = {_0, _1088} + {_0, _3805};
  wire [1:0] _28188 = {_0, _4415} + {_0, _6397};
  wire [2:0] _28189 = {_0, _28187} + {_0, _28188};
  wire [1:0] _28190 = {_0, _9566} + {_0, _12282};
  wire [3:0] _28191 = {_0, _28189} + {_0, _0, _28190};
  wire _28192 = _12301 < _28191;
  wire _28193 = r282 ^ _28192;
  wire _28194 = _12298 ? coded_block[282] : r282;
  wire _28195 = _12296 ? _28193 : _28194;
  always @ (posedge reset or posedge clock) if (reset) r282 <= 1'd0; else if (_12300) r282 <= _28195;
  wire [1:0] _28196 = {_0, _1120} + {_0, _4060};
  wire [1:0] _28197 = {_0, _5884} + {_0, _6494};
  wire [2:0] _28198 = {_0, _28196} + {_0, _28197};
  wire [1:0] _28199 = {_0, _8480} + {_0, _11644};
  wire [3:0] _28200 = {_0, _28198} + {_0, _0, _28199};
  wire _28201 = _12301 < _28200;
  wire _28202 = r281 ^ _28201;
  wire _28203 = _12298 ? coded_block[281] : r281;
  wire _28204 = _12296 ? _28202 : _28203;
  always @ (posedge reset or posedge clock) if (reset) r281 <= 1'd0; else if (_12300) r281 <= _28204;
  wire [1:0] _28205 = {_0, _1151} + {_0, _2941};
  wire [1:0] _28206 = {_0, _6139} + {_0, _7965};
  wire [2:0] _28207 = {_0, _28205} + {_0, _28206};
  wire [1:0] _28208 = {_0, _8574} + {_0, _10558};
  wire [3:0] _28209 = {_0, _28207} + {_0, _0, _28208};
  wire _28210 = _12301 < _28209;
  wire _28211 = r280 ^ _28210;
  wire _28212 = _12298 ? coded_block[280] : r280;
  wire _28213 = _12296 ? _28211 : _28212;
  always @ (posedge reset or posedge clock) if (reset) r280 <= 1'd0; else if (_12300) r280 <= _28213;
  wire [1:0] _28214 = {_0, _34} + {_0, _3964};
  wire [1:0] _28215 = {_0, _6045} + {_0, _8123};
  wire [2:0] _28216 = {_0, _28214} + {_0, _28215};
  wire [1:0] _28217 = {_0, _10204} + {_0, _12282};
  wire [3:0] _28218 = {_0, _28216} + {_0, _0, _28217};
  wire _28219 = _12301 < _28218;
  wire _28220 = r279 ^ _28219;
  wire _28221 = _12298 ? coded_block[279] : r279;
  wire _28222 = _12296 ? _28220 : _28221;
  always @ (posedge reset or posedge clock) if (reset) r279 <= 1'd0; else if (_12300) r279 <= _28222;
  wire [1:0] _28223 = {_0, _639} + {_0, _2430};
  wire [1:0] _28224 = {_0, _5628} + {_0, _7454};
  wire [2:0] _28225 = {_0, _28223} + {_0, _28224};
  wire [1:0] _28226 = {_0, _10077} + {_0, _12061};
  wire [3:0] _28227 = {_0, _28225} + {_0, _0, _28226};
  wire _28228 = _12301 < _28227;
  wire _28229 = r278 ^ _28228;
  wire _28230 = _12298 ? coded_block[278] : r278;
  wire _28231 = _12296 ? _28229 : _28230;
  always @ (posedge reset or posedge clock) if (reset) r278 <= 1'd0; else if (_12300) r278 <= _28231;
  wire [1:0] _28232 = {_0, _672} + {_0, _4091};
  wire [1:0] _28233 = {_0, _4511} + {_0, _7710};
  wire [2:0] _28234 = {_0, _28232} + {_0, _28233};
  wire [1:0] _28235 = {_0, _9534} + {_0, _12155};
  wire [3:0] _28236 = {_0, _28234} + {_0, _0, _28235};
  wire _28237 = _12301 < _28236;
  wire _28238 = r277 ^ _28237;
  wire _28239 = _12298 ? coded_block[277] : r277;
  wire _28240 = _12296 ? _28238 : _28239;
  always @ (posedge reset or posedge clock) if (reset) r277 <= 1'd0; else if (_12300) r277 <= _28240;
  wire [1:0] _28241 = {_0, _703} + {_0, _2302};
  wire [1:0] _28242 = {_0, _4160} + {_0, _6589};
  wire [2:0] _28243 = {_0, _28241} + {_0, _28242};
  wire [1:0] _28244 = {_0, _9790} + {_0, _11613};
  wire [3:0] _28245 = {_0, _28243} + {_0, _0, _28244};
  wire _28246 = _12301 < _28245;
  wire _28247 = r276 ^ _28246;
  wire _28248 = _12298 ? coded_block[276] : r276;
  wire _28249 = _12296 ? _28247 : _28248;
  always @ (posedge reset or posedge clock) if (reset) r276 <= 1'd0; else if (_12300) r276 <= _28249;
  wire [1:0] _28250 = {_0, _735} + {_0, _2175};
  wire [1:0] _28251 = {_0, _4384} + {_0, _6239};
  wire [2:0] _28252 = {_0, _28250} + {_0, _28251};
  wire [1:0] _28253 = {_0, _8670} + {_0, _11869};
  wire [3:0] _28254 = {_0, _28252} + {_0, _0, _28253};
  wire _28255 = _12301 < _28254;
  wire _28256 = r275 ^ _28255;
  wire _28257 = _12298 ? coded_block[275] : r275;
  wire _28258 = _12296 ? _28256 : _28257;
  always @ (posedge reset or posedge clock) if (reset) r275 <= 1'd0; else if (_12300) r275 <= _28258;
  wire [1:0] _28259 = {_0, _766} + {_0, _2526};
  wire [1:0] _28260 = {_0, _4256} + {_0, _6462};
  wire [2:0] _28261 = {_0, _28259} + {_0, _28260};
  wire [1:0] _28262 = {_0, _8319} + {_0, _10748};
  wire [3:0] _28263 = {_0, _28261} + {_0, _0, _28262};
  wire _28264 = _12301 < _28263;
  wire _28265 = r274 ^ _28264;
  wire _28266 = _12298 ? coded_block[274] : r274;
  wire _28267 = _12296 ? _28265 : _28266;
  always @ (posedge reset or posedge clock) if (reset) r274 <= 1'd0; else if (_12300) r274 <= _28267;
  wire [1:0] _28268 = {_0, _800} + {_0, _3262};
  wire [1:0] _28269 = {_0, _4605} + {_0, _6334};
  wire [2:0] _28270 = {_0, _28268} + {_0, _28269};
  wire [1:0] _28271 = {_0, _8543} + {_0, _10399};
  wire [3:0] _28272 = {_0, _28270} + {_0, _0, _28271};
  wire _28273 = _12301 < _28272;
  wire _28274 = r273 ^ _28273;
  wire _28275 = _12298 ? coded_block[273] : r273;
  wire _28276 = _12296 ? _28274 : _28275;
  always @ (posedge reset or posedge clock) if (reset) r273 <= 1'd0; else if (_12300) r273 <= _28276;
  wire [1:0] _28277 = {_0, _863} + {_0, _3422};
  wire [1:0] _28278 = {_0, _5949} + {_0, _7420};
  wire [2:0] _28279 = {_0, _28277} + {_0, _28278};
  wire [1:0] _28280 = {_0, _8767} + {_0, _10493};
  wire [3:0] _28281 = {_0, _28279} + {_0, _0, _28280};
  wire _28282 = _12301 < _28281;
  wire _28283 = r272 ^ _28282;
  wire _28284 = _12298 ? coded_block[272] : r272;
  wire _28285 = _12296 ? _28283 : _28284;
  always @ (posedge reset or posedge clock) if (reset) r272 <= 1'd0; else if (_12300) r272 <= _28285;
  wire [1:0] _28286 = {_0, _927} + {_0, _4060};
  wire [1:0] _28287 = {_0, _5116} + {_0, _7581};
  wire [2:0] _28288 = {_0, _28286} + {_0, _28287};
  wire [1:0] _28289 = {_0, _10108} + {_0, _11581};
  wire [3:0] _28290 = {_0, _28288} + {_0, _0, _28289};
  wire _28291 = _12301 < _28290;
  wire _28292 = r271 ^ _28291;
  wire _28293 = _12298 ? coded_block[271] : r271;
  wire _28294 = _12296 ? _28292 : _28293;
  always @ (posedge reset or posedge clock) if (reset) r271 <= 1'd0; else if (_12300) r271 <= _28294;
  wire [1:0] _28295 = {_0, _958} + {_0, _2463};
  wire [1:0] _28296 = {_0, _6139} + {_0, _7199};
  wire [2:0] _28297 = {_0, _28295} + {_0, _28296};
  wire [1:0] _28298 = {_0, _9661} + {_0, _12188};
  wire [3:0] _28299 = {_0, _28297} + {_0, _0, _28298};
  wire _28300 = _12301 < _28299;
  wire _28301 = r270 ^ _28300;
  wire _28302 = _12298 ? coded_block[270] : r270;
  wire _28303 = _12296 ? _28301 : _28302;
  always @ (posedge reset or posedge clock) if (reset) r270 <= 1'd0; else if (_12300) r270 <= _28303;
  wire [1:0] _28304 = {_0, _990} + {_0, _2941};
  wire [1:0] _28305 = {_0, _4542} + {_0, _6207};
  wire [2:0] _28306 = {_0, _28304} + {_0, _28305};
  wire [1:0] _28307 = {_0, _9279} + {_0, _11740};
  wire [3:0] _28308 = {_0, _28306} + {_0, _0, _28307};
  wire _28309 = _12301 < _28308;
  wire _28310 = r269 ^ _28309;
  wire _28311 = _12298 ? coded_block[269] : r269;
  wire _28312 = _12296 ? _28310 : _28311;
  always @ (posedge reset or posedge clock) if (reset) r269 <= 1'd0; else if (_12300) r269 <= _28312;
  wire [1:0] _28313 = {_0, _1057} + {_0, _3678};
  wire [1:0] _28314 = {_0, _4447} + {_0, _7100};
  wire [2:0] _28315 = {_0, _28313} + {_0, _28314};
  wire [1:0] _28316 = {_0, _8701} + {_0, _10366};
  wire [3:0] _28317 = {_0, _28315} + {_0, _0, _28316};
  wire _28318 = _12301 < _28317;
  wire _28319 = r268 ^ _28318;
  wire _28320 = _12298 ? coded_block[268] : r268;
  wire _28321 = _12296 ? _28319 : _28320;
  always @ (posedge reset or posedge clock) if (reset) r268 <= 1'd0; else if (_12300) r268 <= _28321;
  wire [1:0] _28322 = {_0, _1088} + {_0, _3359};
  wire [1:0] _28323 = {_0, _5757} + {_0, _6525};
  wire [2:0] _28324 = {_0, _28322} + {_0, _28323};
  wire [1:0] _28325 = {_0, _9181} + {_0, _10783};
  wire [3:0] _28326 = {_0, _28324} + {_0, _0, _28325};
  wire _28327 = _12301 < _28326;
  wire _28328 = r267 ^ _28327;
  wire _28329 = _12298 ? coded_block[267] : r267;
  wire _28330 = _12296 ? _28328 : _28329;
  always @ (posedge reset or posedge clock) if (reset) r267 <= 1'd0; else if (_12300) r267 <= _28330;
  wire [1:0] _28331 = {_0, _1120} + {_0, _3517};
  wire [1:0] _28332 = {_0, _5438} + {_0, _7837};
  wire [2:0] _28333 = {_0, _28331} + {_0, _28332};
  wire [1:0] _28334 = {_0, _8607} + {_0, _11259};
  wire [3:0] _28335 = {_0, _28333} + {_0, _0, _28334};
  wire _28336 = _12301 < _28335;
  wire _28337 = r266 ^ _28336;
  wire _28338 = _12298 ? coded_block[266] : r266;
  wire _28339 = _12296 ? _28337 : _28338;
  always @ (posedge reset or posedge clock) if (reset) r266 <= 1'd0; else if (_12300) r266 <= _28339;
  wire [1:0] _28340 = {_0, _1151} + {_0, _3325};
  wire [1:0] _28341 = {_0, _5597} + {_0, _7517};
  wire [2:0] _28342 = {_0, _28340} + {_0, _28341};
  wire [1:0] _28343 = {_0, _9917} + {_0, _10685};
  wire [3:0] _28344 = {_0, _28342} + {_0, _0, _28343};
  wire _28345 = _12301 < _28344;
  wire _28346 = r265 ^ _28345;
  wire _28347 = _12298 ? coded_block[265] : r265;
  wire _28348 = _12296 ? _28346 : _28347;
  always @ (posedge reset or posedge clock) if (reset) r265 <= 1'd0; else if (_12300) r265 <= _28348;
  wire [1:0] _28349 = {_0, _1184} + {_0, _3709};
  wire [1:0] _28350 = {_0, _5407} + {_0, _7675};
  wire [2:0] _28351 = {_0, _28349} + {_0, _28350};
  wire [1:0] _28352 = {_0, _9597} + {_0, _11996};
  wire [3:0] _28353 = {_0, _28351} + {_0, _0, _28352};
  wire _28354 = _12301 < _28353;
  wire _28355 = r264 ^ _28354;
  wire _28356 = _12298 ? coded_block[264] : r264;
  wire _28357 = _12296 ? _28355 : _28356;
  always @ (posedge reset or posedge clock) if (reset) r264 <= 1'd0; else if (_12300) r264 <= _28357;
  wire [1:0] _28358 = {_0, _1215} + {_0, _2847};
  wire [1:0] _28359 = {_0, _5790} + {_0, _7485};
  wire [2:0] _28360 = {_0, _28358} + {_0, _28359};
  wire [1:0] _28361 = {_0, _9759} + {_0, _11677};
  wire [3:0] _28362 = {_0, _28360} + {_0, _0, _28361};
  wire _28363 = _12301 < _28362;
  wire _28364 = r263 ^ _28363;
  wire _28365 = _12298 ? coded_block[263] : r263;
  wire _28366 = _12296 ? _28364 : _28365;
  always @ (posedge reset or posedge clock) if (reset) r263 <= 1'd0; else if (_12300) r263 <= _28366;
  wire [1:0] _28367 = {_0, _1247} + {_0, _2623};
  wire [1:0] _28368 = {_0, _4926} + {_0, _7868};
  wire [2:0] _28369 = {_0, _28367} + {_0, _28368};
  wire [1:0] _28370 = {_0, _9566} + {_0, _11837};
  wire [3:0] _28371 = {_0, _28369} + {_0, _0, _28370};
  wire _28372 = _12301 < _28371;
  wire _28373 = r262 ^ _28372;
  wire _28374 = _12298 ? coded_block[262] : r262;
  wire _28375 = _12296 ? _28373 : _28374;
  always @ (posedge reset or posedge clock) if (reset) r262 <= 1'd0; else if (_12300) r262 <= _28375;
  wire [1:0] _28376 = {_0, _1278} + {_0, _3198};
  wire [1:0] _28377 = {_0, _4703} + {_0, _7005};
  wire [2:0] _28378 = {_0, _28376} + {_0, _28377};
  wire [1:0] _28379 = {_0, _9949} + {_0, _11644};
  wire [3:0] _28380 = {_0, _28378} + {_0, _0, _28379};
  wire _28381 = _12301 < _28380;
  wire _28382 = r261 ^ _28381;
  wire _28383 = _12298 ? coded_block[261] : r261;
  wire _28384 = _12296 ? _28382 : _28383;
  always @ (posedge reset or posedge clock) if (reset) r261 <= 1'd0; else if (_12300) r261 <= _28384;
  wire [1:0] _28385 = {_0, _1312} + {_0, _3135};
  wire [1:0] _28386 = {_0, _5279} + {_0, _6781};
  wire [2:0] _28387 = {_0, _28385} + {_0, _28386};
  wire [1:0] _28388 = {_0, _9085} + {_0, _12027};
  wire [3:0] _28389 = {_0, _28387} + {_0, _0, _28388};
  wire _28390 = _12301 < _28389;
  wire _28391 = r260 ^ _28390;
  wire _28392 = _12298 ? coded_block[260] : r260;
  wire _28393 = _12296 ? _28391 : _28392;
  always @ (posedge reset or posedge clock) if (reset) r260 <= 1'd0; else if (_12300) r260 <= _28393;
  wire [1:0] _28394 = {_0, _1343} + {_0, _2239};
  wire [1:0] _28395 = {_0, _5215} + {_0, _7357};
  wire [2:0] _28396 = {_0, _28394} + {_0, _28395};
  wire [1:0] _28397 = {_0, _8863} + {_0, _11165};
  wire [3:0] _28398 = {_0, _28396} + {_0, _0, _28397};
  wire _28399 = _12301 < _28398;
  wire _28400 = r259 ^ _28399;
  wire _28401 = _12298 ? coded_block[259] : r259;
  wire _28402 = _12296 ? _28400 : _28401;
  always @ (posedge reset or posedge clock) if (reset) r259 <= 1'd0; else if (_12300) r259 <= _28402;
  wire [1:0] _28403 = {_0, _1375} + {_0, _2910};
  wire [1:0] _28404 = {_0, _4319} + {_0, _7293};
  wire [2:0] _28405 = {_0, _28403} + {_0, _28404};
  wire [1:0] _28406 = {_0, _9438} + {_0, _10941};
  wire [3:0] _28407 = {_0, _28405} + {_0, _0, _28406};
  wire _28408 = _12301 < _28407;
  wire _28409 = r258 ^ _28408;
  wire _28410 = _12298 ? coded_block[258] : r258;
  wire _28411 = _12296 ? _28409 : _28410;
  always @ (posedge reset or posedge clock) if (reset) r258 <= 1'd0; else if (_12300) r258 <= _28411;
  wire [1:0] _28412 = {_0, _1406} + {_0, _2494};
  wire [1:0] _28413 = {_0, _4989} + {_0, _6397};
  wire [2:0] _28414 = {_0, _28412} + {_0, _28413};
  wire [1:0] _28415 = {_0, _9375} + {_0, _11516};
  wire [3:0] _28416 = {_0, _28414} + {_0, _0, _28415};
  wire _28417 = _12301 < _28416;
  wire _28418 = r257 ^ _28417;
  wire _28419 = _12298 ? coded_block[257] : r257;
  wire _28420 = _12296 ? _28418 : _28419;
  always @ (posedge reset or posedge clock) if (reset) r257 <= 1'd0; else if (_12300) r257 <= _28420;
  wire [1:0] _28421 = {_0, _1439} + {_0, _2208};
  wire [1:0] _28422 = {_0, _4574} + {_0, _7069};
  wire [2:0] _28423 = {_0, _28421} + {_0, _28422};
  wire [1:0] _28424 = {_0, _8480} + {_0, _11453};
  wire [3:0] _28425 = {_0, _28423} + {_0, _0, _28424};
  wire _28426 = _12301 < _28425;
  wire _28427 = r256 ^ _28426;
  wire _28428 = _12298 ? coded_block[256] : r256;
  wire _28429 = _12296 ? _28427 : _28428;
  always @ (posedge reset or posedge clock) if (reset) r256 <= 1'd0; else if (_12300) r256 <= _28429;
  wire [1:0] _28430 = {_0, _1470} + {_0, _3167};
  wire [1:0] _28431 = {_0, _4287} + {_0, _6652};
  wire [2:0] _28432 = {_0, _28430} + {_0, _28431};
  wire [1:0] _28433 = {_0, _9149} + {_0, _10558};
  wire [3:0] _28434 = {_0, _28432} + {_0, _0, _28433};
  wire _28435 = _12301 < _28434;
  wire _28436 = r255 ^ _28435;
  wire _28437 = _12298 ? coded_block[255] : r255;
  wire _28438 = _12296 ? _28436 : _28437;
  always @ (posedge reset or posedge clock) if (reset) r255 <= 1'd0; else if (_12300) r255 <= _28438;
  wire [1:0] _28439 = {_0, _1502} + {_0, _2655};
  wire [1:0] _28440 = {_0, _5246} + {_0, _6366};
  wire [2:0] _28441 = {_0, _28439} + {_0, _28440};
  wire [1:0] _28442 = {_0, _8736} + {_0, _11228};
  wire [3:0] _28443 = {_0, _28441} + {_0, _0, _28442};
  wire _28444 = _12301 < _28443;
  wire _28445 = r254 ^ _28444;
  wire _28446 = _12298 ? coded_block[254] : r254;
  wire _28447 = _12296 ? _28445 : _28446;
  always @ (posedge reset or posedge clock) if (reset) r254 <= 1'd0; else if (_12300) r254 <= _28447;
  wire [1:0] _28448 = {_0, _1533} + {_0, _3646};
  wire [1:0] _28449 = {_0, _4734} + {_0, _7326};
  wire [2:0] _28450 = {_0, _28448} + {_0, _28449};
  wire [1:0] _28451 = {_0, _8446} + {_0, _10814};
  wire [3:0] _28452 = {_0, _28450} + {_0, _0, _28451};
  wire _28453 = _12301 < _28452;
  wire _28454 = r253 ^ _28453;
  wire _28455 = _12298 ? coded_block[253] : r253;
  wire _28456 = _12296 ? _28454 : _28455;
  always @ (posedge reset or posedge clock) if (reset) r253 <= 1'd0; else if (_12300) r253 <= _28456;
  wire [1:0] _28457 = {_0, _1599} + {_0, _3580};
  wire [1:0] _28458 = {_0, _4478} + {_0, _7804};
  wire [2:0] _28459 = {_0, _28457} + {_0, _28458};
  wire [1:0] _28460 = {_0, _8894} + {_0, _11485};
  wire [3:0] _28461 = {_0, _28459} + {_0, _0, _28460};
  wire _28462 = _12301 < _28461;
  wire _28463 = r252 ^ _28462;
  wire _28464 = _12298 ? coded_block[252] : r252;
  wire _28465 = _12296 ? _28463 : _28464;
  always @ (posedge reset or posedge clock) if (reset) r252 <= 1'd0; else if (_12300) r252 <= _28465;
  wire [1:0] _28466 = {_0, _1631} + {_0, _3104};
  wire [1:0] _28467 = {_0, _5663} + {_0, _6558};
  wire [2:0] _28468 = {_0, _28466} + {_0, _28467};
  wire [1:0] _28469 = {_0, _9886} + {_0, _10973};
  wire [3:0] _28470 = {_0, _28468} + {_0, _0, _28469};
  wire _28471 = _12301 < _28470;
  wire _28472 = r251 ^ _28471;
  wire _28473 = _12298 ? coded_block[251] : r251;
  wire _28474 = _12296 ? _28472 : _28473;
  always @ (posedge reset or posedge clock) if (reset) r251 <= 1'd0; else if (_12300) r251 <= _28474;
  wire [1:0] _28475 = {_0, _1662} + {_0, _3231};
  wire [1:0] _28476 = {_0, _5183} + {_0, _7741};
  wire [2:0] _28477 = {_0, _28475} + {_0, _28476};
  wire [1:0] _28478 = {_0, _8638} + {_0, _11964};
  wire [3:0] _28479 = {_0, _28477} + {_0, _0, _28478};
  wire _28480 = _12301 < _28479;
  wire _28481 = r250 ^ _28480;
  wire _28482 = _12298 ? coded_block[250] : r250;
  wire _28483 = _12296 ? _28481 : _28482;
  always @ (posedge reset or posedge clock) if (reset) r250 <= 1'd0; else if (_12300) r250 <= _28483;
  wire [1:0] _28484 = {_0, _1726} + {_0, _3805};
  wire [1:0] _28485 = {_0, _4640} + {_0, _7389};
  wire [2:0] _28486 = {_0, _28484} + {_0, _28485};
  wire [1:0] _28487 = {_0, _9342} + {_0, _11900};
  wire [3:0] _28488 = {_0, _28486} + {_0, _0, _28487};
  wire _28489 = _12301 < _28488;
  wire _28490 = r249 ^ _28489;
  wire _28491 = _12298 ? coded_block[249] : r249;
  wire _28492 = _12296 ? _28490 : _28491;
  always @ (posedge reset or posedge clock) if (reset) r249 <= 1'd0; else if (_12300) r249 <= _28492;
  wire [1:0] _28493 = {_0, _1789} + {_0, _2592};
  wire [1:0] _28494 = {_0, _5853} + {_0, _7965};
  wire [2:0] _28495 = {_0, _28493} + {_0, _28494};
  wire [1:0] _28496 = {_0, _8799} + {_0, _11550};
  wire [3:0] _28497 = {_0, _28495} + {_0, _0, _28496};
  wire _28498 = _12301 < _28497;
  wire _28499 = r248 ^ _28498;
  wire _28500 = _12298 ? coded_block[248] : r248;
  wire _28501 = _12296 ? _28499 : _28500;
  always @ (posedge reset or posedge clock) if (reset) r248 <= 1'd0; else if (_12300) r248 <= _28501;
  wire [1:0] _28502 = {_0, _1823} + {_0, _2878};
  wire [1:0] _28503 = {_0, _4671} + {_0, _7931};
  wire [2:0] _28504 = {_0, _28502} + {_0, _28503};
  wire [1:0] _28505 = {_0, _10045} + {_0, _10877};
  wire [3:0] _28506 = {_0, _28504} + {_0, _0, _28505};
  wire _28507 = _12301 < _28506;
  wire _28508 = r247 ^ _28507;
  wire _28509 = _12298 ? coded_block[247] : r247;
  wire _28510 = _12296 ? _28508 : _28509;
  always @ (posedge reset or posedge clock) if (reset) r247 <= 1'd0; else if (_12300) r247 <= _28510;
  wire [1:0] _28511 = {_0, _1854} + {_0, _2271};
  wire [1:0] _28512 = {_0, _4958} + {_0, _6750};
  wire [2:0] _28513 = {_0, _28511} + {_0, _28512};
  wire [1:0] _28514 = {_0, _10014} + {_0, _12124};
  wire [3:0] _28515 = {_0, _28513} + {_0, _0, _28514};
  wire _28516 = _12301 < _28515;
  wire _28517 = r246 ^ _28516;
  wire _28518 = _12298 ? coded_block[246] : r246;
  wire _28519 = _12296 ? _28517 : _28518;
  always @ (posedge reset or posedge clock) if (reset) r246 <= 1'd0; else if (_12300) r246 <= _28519;
  wire [1:0] _28520 = {_0, _1917} + {_0, _2081};
  wire [1:0] _28521 = {_0, _4192} + {_0, _6431};
  wire [2:0] _28522 = {_0, _28520} + {_0, _28521};
  wire [1:0] _28523 = {_0, _9118} + {_0, _10910};
  wire [3:0] _28524 = {_0, _28522} + {_0, _0, _28523};
  wire _28525 = _12301 < _28524;
  wire _28526 = r245 ^ _28525;
  wire _28527 = _12298 ? coded_block[245] : r245;
  wire _28528 = _12296 ? _28526 : _28527;
  always @ (posedge reset or posedge clock) if (reset) r245 <= 1'd0; else if (_12300) r245 <= _28528;
  wire [1:0] _28529 = {_0, _1950} + {_0, _2144};
  wire [1:0] _28530 = {_0, _4129} + {_0, _6270};
  wire [2:0] _28531 = {_0, _28529} + {_0, _28530};
  wire [1:0] _28532 = {_0, _8511} + {_0, _11196};
  wire [3:0] _28533 = {_0, _28531} + {_0, _0, _28532};
  wire _28534 = _12301 < _28533;
  wire _28535 = r244 ^ _28534;
  wire _28536 = _12298 ? coded_block[244] : r244;
  wire _28537 = _12296 ? _28535 : _28536;
  always @ (posedge reset or posedge clock) if (reset) r244 <= 1'd0; else if (_12300) r244 <= _28537;
  wire [1:0] _28538 = {_0, _1981} + {_0, _2336};
  wire [1:0] _28539 = {_0, _4223} + {_0, _6176};
  wire [2:0] _28540 = {_0, _28538} + {_0, _28539};
  wire [1:0] _28541 = {_0, _8352} + {_0, _10590};
  wire [3:0] _28542 = {_0, _28540} + {_0, _0, _28541};
  wire _28543 = _12301 < _28542;
  wire _28544 = r243 ^ _28543;
  wire _28545 = _12298 ? coded_block[243] : r243;
  wire _28546 = _12296 ? _28544 : _28545;
  always @ (posedge reset or posedge clock) if (reset) r243 <= 1'd0; else if (_12300) r243 <= _28546;
  wire [1:0] _28547 = {_0, _2013} + {_0, _2974};
  wire [1:0] _28548 = {_0, _4415} + {_0, _6303};
  wire [2:0] _28549 = {_0, _28547} + {_0, _28548};
  wire [1:0] _28550 = {_0, _8225} + {_0, _10430};
  wire [3:0] _28551 = {_0, _28549} + {_0, _0, _28550};
  wire _28552 = _12301 < _28551;
  wire _28553 = r242 ^ _28552;
  wire _28554 = _12298 ? coded_block[242] : r242;
  wire _28555 = _12296 ? _28553 : _28554;
  always @ (posedge reset or posedge clock) if (reset) r242 <= 1'd0; else if (_12300) r242 <= _28555;
  wire [1:0] _28556 = {_0, _65} + {_0, _3933};
  wire [1:0] _28557 = {_0, _4798} + {_0, _7132};
  wire [2:0] _28558 = {_0, _28556} + {_0, _28557};
  wire [1:0] _28559 = {_0, _8574} + {_0, _10462};
  wire [3:0] _28560 = {_0, _28558} + {_0, _0, _28559};
  wire _28561 = _12301 < _28560;
  wire _28562 = r241 ^ _28561;
  wire _28563 = _12298 ? coded_block[241] : r241;
  wire _28564 = _12296 ? _28562 : _28563;
  always @ (posedge reset or posedge clock) if (reset) r241 <= 1'd0; else if (_12300) r241 <= _28564;
  wire [1:0] _28565 = {_0, _97} + {_0, _3997};
  wire [1:0] _28566 = {_0, _6012} + {_0, _6877};
  wire [2:0] _28567 = {_0, _28565} + {_0, _28566};
  wire [1:0] _28568 = {_0, _9212} + {_0, _10654};
  wire [3:0] _28569 = {_0, _28567} + {_0, _0, _28568};
  wire _28570 = _12301 < _28569;
  wire _28571 = r240 ^ _28570;
  wire _28572 = _12298 ? coded_block[240] : r240;
  wire _28573 = _12296 ? _28571 : _28572;
  always @ (posedge reset or posedge clock) if (reset) r240 <= 1'd0; else if (_12300) r240 <= _28573;
  wire [1:0] _28574 = {_0, _128} + {_0, _2782};
  wire [1:0] _28575 = {_0, _6076} + {_0, _8092};
  wire [2:0] _28576 = {_0, _28574} + {_0, _28575};
  wire [1:0] _28577 = {_0, _8957} + {_0, _11295};
  wire [3:0] _28578 = {_0, _28576} + {_0, _0, _28577};
  wire _28579 = _12301 < _28578;
  wire _28580 = r239 ^ _28579;
  wire _28581 = _12298 ? coded_block[239] : r239;
  wire _28582 = _12296 ? _28580 : _28581;
  always @ (posedge reset or posedge clock) if (reset) r239 <= 1'd0; else if (_12300) r239 <= _28582;
  wire [1:0] _28583 = {_0, _161} + {_0, _3486};
  wire [1:0] _28584 = {_0, _4861} + {_0, _8155};
  wire [2:0] _28585 = {_0, _28583} + {_0, _28584};
  wire [1:0] _28586 = {_0, _10172} + {_0, _11038};
  wire [3:0] _28587 = {_0, _28585} + {_0, _0, _28586};
  wire _28588 = _12301 < _28587;
  wire _28589 = r238 ^ _28588;
  wire _28590 = _12298 ? coded_block[238] : r238;
  wire _28591 = _12296 ? _28589 : _28590;
  always @ (posedge reset or posedge clock) if (reset) r238 <= 1'd0; else if (_12300) r238 <= _28591;
  wire [1:0] _28592 = {_0, _192} + {_0, _3390};
  wire [1:0] _28593 = {_0, _5565} + {_0, _6942};
  wire [2:0] _28594 = {_0, _28592} + {_0, _28593};
  wire [1:0] _28595 = {_0, _10235} + {_0, _12251};
  wire [3:0] _28596 = {_0, _28594} + {_0, _0, _28595};
  wire _28597 = _12301 < _28596;
  wire _28598 = r237 ^ _28597;
  wire _28599 = _12298 ? coded_block[237] : r237;
  wire _28600 = _12296 ? _28598 : _28599;
  always @ (posedge reset or posedge clock) if (reset) r237 <= 1'd0; else if (_12300) r237 <= _28600;
  wire [1:0] _28601 = {_0, _224} + {_0, _3901};
  wire [1:0] _28602 = {_0, _5470} + {_0, _7644};
  wire [2:0] _28603 = {_0, _28601} + {_0, _28602};
  wire [1:0] _28604 = {_0, _9022} + {_0, _10303};
  wire [3:0] _28605 = {_0, _28603} + {_0, _0, _28604};
  wire _28606 = _12301 < _28605;
  wire _28607 = r236 ^ _28606;
  wire _28608 = _12298 ? coded_block[236] : r236;
  wire _28609 = _12296 ? _28607 : _28608;
  always @ (posedge reset or posedge clock) if (reset) r236 <= 1'd0; else if (_12300) r236 <= _28609;
  wire [1:0] _28610 = {_0, _255} + {_0, _2750};
  wire [1:0] _28611 = {_0, _5981} + {_0, _7548};
  wire [2:0] _28612 = {_0, _28610} + {_0, _28611};
  wire [1:0] _28613 = {_0, _9724} + {_0, _11101};
  wire [3:0] _28614 = {_0, _28612} + {_0, _0, _28613};
  wire _28615 = _12301 < _28614;
  wire _28616 = r235 ^ _28615;
  wire _28617 = _12298 ? coded_block[235] : r235;
  wire _28618 = _12296 ? _28616 : _28617;
  always @ (posedge reset or posedge clock) if (reset) r235 <= 1'd0; else if (_12300) r235 <= _28618;
  wire [1:0] _28619 = {_0, _320} + {_0, _3068};
  wire [1:0] _28620 = {_0, _6108} + {_0, _6908};
  wire [2:0] _28621 = {_0, _28619} + {_0, _28620};
  wire [1:0] _28622 = {_0, _10141} + {_0, _11708};
  wire [3:0] _28623 = {_0, _28621} + {_0, _0, _28622};
  wire _28624 = _12301 < _28623;
  wire _28625 = r234 ^ _28624;
  wire _28626 = _12298 ? coded_block[234] : r234;
  wire _28627 = _12296 ? _28625 : _28626;
  always @ (posedge reset or posedge clock) if (reset) r234 <= 1'd0; else if (_12300) r234 <= _28627;
  wire [1:0] _28628 = {_0, _352} + {_0, _3615};
  wire [1:0] _28629 = {_0, _5152} + {_0, _8186};
  wire [2:0] _28630 = {_0, _28628} + {_0, _28629};
  wire [1:0] _28631 = {_0, _8991} + {_0, _12219};
  wire [3:0] _28632 = {_0, _28630} + {_0, _0, _28631};
  wire _28633 = _12301 < _28632;
  wire _28634 = r233 ^ _28633;
  wire _28635 = _12298 ? coded_block[233] : r233;
  wire _28636 = _12296 ? _28634 : _28635;
  always @ (posedge reset or posedge clock) if (reset) r233 <= 1'd0; else if (_12300) r233 <= _28636;
  wire [1:0] _28637 = {_0, _383} + {_0, _2686};
  wire [1:0] _28638 = {_0, _5694} + {_0, _7230};
  wire [2:0] _28639 = {_0, _28637} + {_0, _28638};
  wire [1:0] _28640 = {_0, _8256} + {_0, _11069};
  wire [3:0] _28641 = {_0, _28639} + {_0, _0, _28640};
  wire _28642 = _12301 < _28641;
  wire _28643 = r232 ^ _28642;
  wire _28644 = _12298 ? coded_block[232] : r232;
  wire _28645 = _12296 ? _28643 : _28644;
  always @ (posedge reset or posedge clock) if (reset) r232 <= 1'd0; else if (_12300) r232 <= _28645;
  wire [1:0] _28646 = {_0, _416} + {_0, _3005};
  wire [1:0] _28647 = {_0, _4767} + {_0, _7773};
  wire [2:0] _28648 = {_0, _28646} + {_0, _28647};
  wire [1:0] _28649 = {_0, _9311} + {_0, _10335};
  wire [3:0] _28650 = {_0, _28648} + {_0, _0, _28649};
  wire _28651 = _12301 < _28650;
  wire _28652 = r231 ^ _28651;
  wire _28653 = _12298 ? coded_block[231] : r231;
  wire _28654 = _12296 ? _28652 : _28653;
  always @ (posedge reset or posedge clock) if (reset) r231 <= 1'd0; else if (_12300) r231 <= _28654;
  wire [1:0] _28655 = {_0, _447} + {_0, _3453};
  wire [1:0] _28656 = {_0, _5085} + {_0, _6845};
  wire [2:0] _28657 = {_0, _28655} + {_0, _28656};
  wire [1:0] _28658 = {_0, _9853} + {_0, _11389};
  wire [3:0] _28659 = {_0, _28657} + {_0, _0, _28658};
  wire _28660 = _12301 < _28659;
  wire _28661 = r230 ^ _28660;
  wire _28662 = _12298 ? coded_block[230] : r230;
  wire _28663 = _12296 ? _28661 : _28662;
  always @ (posedge reset or posedge clock) if (reset) r230 <= 1'd0; else if (_12300) r230 <= _28663;
  wire [1:0] _28664 = {_0, _479} + {_0, _2813};
  wire [1:0] _28665 = {_0, _5534} + {_0, _7163};
  wire [2:0] _28666 = {_0, _28664} + {_0, _28665};
  wire [1:0] _28667 = {_0, _8926} + {_0, _11933};
  wire [3:0] _28668 = {_0, _28666} + {_0, _0, _28667};
  wire _28669 = _12301 < _28668;
  wire _28670 = r229 ^ _28669;
  wire _28671 = _12298 ? coded_block[229] : r229;
  wire _28672 = _12296 ? _28670 : _28671;
  always @ (posedge reset or posedge clock) if (reset) r229 <= 1'd0; else if (_12300) r229 <= _28672;
  wire [1:0] _28673 = {_0, _510} + {_0, _3742};
  wire [1:0] _28674 = {_0, _4895} + {_0, _7612};
  wire [2:0] _28675 = {_0, _28673} + {_0, _28674};
  wire [1:0] _28676 = {_0, _9248} + {_0, _11004};
  wire [3:0] _28677 = {_0, _28675} + {_0, _0, _28676};
  wire _28678 = _12301 < _28677;
  wire _28679 = r228 ^ _28678;
  wire _28680 = _12298 ? coded_block[228] : r228;
  wire _28681 = _12296 ? _28679 : _28680;
  always @ (posedge reset or posedge clock) if (reset) r228 <= 1'd0; else if (_12300) r228 <= _28681;
  wire [1:0] _28682 = {_0, _545} + {_0, _3836};
  wire [1:0] _28683 = {_0, _5821} + {_0, _6973};
  wire [2:0] _28684 = {_0, _28682} + {_0, _28683};
  wire [1:0] _28685 = {_0, _9693} + {_0, _11326};
  wire [3:0] _28686 = {_0, _28684} + {_0, _0, _28685};
  wire _28687 = _12301 < _28686;
  wire _28688 = r227 ^ _28687;
  wire _28689 = _12298 ? coded_block[227] : r227;
  wire _28690 = _12296 ? _28688 : _28689;
  always @ (posedge reset or posedge clock) if (reset) r227 <= 1'd0; else if (_12300) r227 <= _28690;
  wire [1:0] _28691 = {_0, _576} + {_0, _3294};
  wire [1:0] _28692 = {_0, _5918} + {_0, _7900};
  wire [2:0] _28693 = {_0, _28691} + {_0, _28692};
  wire [1:0] _28694 = {_0, _9054} + {_0, _11771};
  wire [3:0] _28695 = {_0, _28693} + {_0, _0, _28694};
  wire _28696 = _12301 < _28695;
  wire _28697 = r226 ^ _28696;
  wire _28698 = _12298 ? coded_block[226] : r226;
  wire _28699 = _12296 ? _28697 : _28698;
  always @ (posedge reset or posedge clock) if (reset) r226 <= 1'd0; else if (_12300) r226 <= _28699;
  wire [1:0] _28700 = {_0, _608} + {_0, _3549};
  wire [1:0] _28701 = {_0, _5373} + {_0, _7996};
  wire [2:0] _28702 = {_0, _28700} + {_0, _28701};
  wire [1:0] _28703 = {_0, _9980} + {_0, _11132};
  wire [3:0] _28704 = {_0, _28702} + {_0, _0, _28703};
  wire _28705 = _12301 < _28704;
  wire _28706 = r225 ^ _28705;
  wire _28707 = _12298 ? coded_block[225] : r225;
  wire _28708 = _12296 ? _28706 : _28707;
  always @ (posedge reset or posedge clock) if (reset) r225 <= 1'd0; else if (_12300) r225 <= _28708;
  wire [1:0] _28709 = {_0, _34} + {_0, _3005};
  wire [1:0] _28710 = {_0, _5085} + {_0, _7163};
  wire [2:0] _28711 = {_0, _28709} + {_0, _28710};
  wire [1:0] _28712 = {_0, _9248} + {_0, _11326};
  wire [3:0] _28713 = {_0, _28711} + {_0, _0, _28712};
  wire _28714 = _12301 < _28713;
  wire _28715 = r224 ^ _28714;
  wire _28716 = _12298 ? coded_block[224] : r224;
  wire _28717 = _12296 ? _28715 : _28716;
  always @ (posedge reset or posedge clock) if (reset) r224 <= 1'd0; else if (_12300) r224 <= _28717;
  wire [1:0] _28718 = {_0, _65} + {_0, _3422};
  wire [1:0] _28719 = {_0, _6076} + {_0, _7675};
  wire [2:0] _28720 = {_0, _28718} + {_0, _28719};
  wire [1:0] _28721 = {_0, _9342} + {_0, _10399};
  wire [3:0] _28722 = {_0, _28720} + {_0, _0, _28721};
  wire _28723 = _12301 < _28722;
  wire _28724 = r223 ^ _28723;
  wire _28725 = _12298 ? coded_block[223] : r223;
  wire _28726 = _12296 ? _28724 : _28725;
  always @ (posedge reset or posedge clock) if (reset) r223 <= 1'd0; else if (_12300) r223 <= _28726;
  wire [1:0] _28727 = {_0, _97} + {_0, _2719};
  wire [1:0] _28728 = {_0, _5501} + {_0, _8155};
  wire [2:0] _28729 = {_0, _28727} + {_0, _28728};
  wire [1:0] _28730 = {_0, _9759} + {_0, _11422};
  wire [3:0] _28731 = {_0, _28729} + {_0, _0, _28730};
  wire _28732 = _12301 < _28731;
  wire _28733 = r222 ^ _28732;
  wire _28734 = _12298 ? coded_block[222] : r222;
  wire _28735 = _12296 ? _28733 : _28734;
  always @ (posedge reset or posedge clock) if (reset) r222 <= 1'd0; else if (_12300) r222 <= _28735;
  wire [1:0] _28736 = {_0, _128} + {_0, _2399};
  wire [1:0] _28737 = {_0, _4798} + {_0, _7581};
  wire [2:0] _28738 = {_0, _28736} + {_0, _28737};
  wire [1:0] _28739 = {_0, _10235} + {_0, _11837};
  wire [3:0] _28740 = {_0, _28738} + {_0, _0, _28739};
  wire _28741 = _12301 < _28740;
  wire _28742 = r221 ^ _28741;
  wire _28743 = _12298 ? coded_block[221] : r221;
  wire _28744 = _12296 ? _28742 : _28743;
  always @ (posedge reset or posedge clock) if (reset) r221 <= 1'd0; else if (_12300) r221 <= _28744;
  wire [1:0] _28745 = {_0, _161} + {_0, _2557};
  wire [1:0] _28746 = {_0, _4478} + {_0, _6877};
  wire [2:0] _28747 = {_0, _28745} + {_0, _28746};
  wire [1:0] _28748 = {_0, _9661} + {_0, _10303};
  wire [3:0] _28749 = {_0, _28747} + {_0, _0, _28748};
  wire _28750 = _12301 < _28749;
  wire _28751 = r220 ^ _28750;
  wire _28752 = _12298 ? coded_block[220] : r220;
  wire _28753 = _12296 ? _28751 : _28752;
  always @ (posedge reset or posedge clock) if (reset) r220 <= 1'd0; else if (_12300) r220 <= _28753;
  wire [1:0] _28754 = {_0, _192} + {_0, _2367};
  wire [1:0] _28755 = {_0, _4640} + {_0, _6558};
  wire [2:0] _28756 = {_0, _28754} + {_0, _28755};
  wire [1:0] _28757 = {_0, _8957} + {_0, _11740};
  wire [3:0] _28758 = {_0, _28756} + {_0, _0, _28757};
  wire _28759 = _12301 < _28758;
  wire _28760 = r219 ^ _28759;
  wire _28761 = _12298 ? coded_block[219] : r219;
  wire _28762 = _12296 ? _28760 : _28761;
  always @ (posedge reset or posedge clock) if (reset) r219 <= 1'd0; else if (_12300) r219 <= _28762;
  wire [1:0] _28763 = {_0, _224} + {_0, _2750};
  wire [1:0] _28764 = {_0, _4447} + {_0, _6718};
  wire [2:0] _28765 = {_0, _28763} + {_0, _28764};
  wire [1:0] _28766 = {_0, _8638} + {_0, _11038};
  wire [3:0] _28767 = {_0, _28765} + {_0, _0, _28766};
  wire _28768 = _12301 < _28767;
  wire _28769 = r218 ^ _28768;
  wire _28770 = _12298 ? coded_block[218] : r218;
  wire _28771 = _12296 ? _28769 : _28770;
  always @ (posedge reset or posedge clock) if (reset) r218 <= 1'd0; else if (_12300) r218 <= _28771;
  wire [1:0] _28772 = {_0, _255} + {_0, _3901};
  wire [1:0] _28773 = {_0, _4830} + {_0, _6525};
  wire [2:0] _28774 = {_0, _28772} + {_0, _28773};
  wire [1:0] _28775 = {_0, _8799} + {_0, _10717};
  wire [3:0] _28776 = {_0, _28774} + {_0, _0, _28775};
  wire _28777 = _12301 < _28776;
  wire _28778 = r217 ^ _28777;
  wire _28779 = _12298 ? coded_block[217] : r217;
  wire _28780 = _12296 ? _28778 : _28779;
  always @ (posedge reset or posedge clock) if (reset) r217 <= 1'd0; else if (_12300) r217 <= _28780;
  wire [1:0] _28781 = {_0, _289} + {_0, _3678};
  wire [1:0] _28782 = {_0, _5981} + {_0, _6908};
  wire [2:0] _28783 = {_0, _28781} + {_0, _28782};
  wire [1:0] _28784 = {_0, _8607} + {_0, _10877};
  wire [3:0] _28785 = {_0, _28783} + {_0, _0, _28784};
  wire _28786 = _12301 < _28785;
  wire _28787 = r216 ^ _28786;
  wire _28788 = _12298 ? coded_block[216] : r216;
  wire _28789 = _12296 ? _28787 : _28788;
  always @ (posedge reset or posedge clock) if (reset) r216 <= 1'd0; else if (_12300) r216 <= _28789;
  wire [1:0] _28790 = {_0, _320} + {_0, _2239};
  wire [1:0] _28791 = {_0, _5757} + {_0, _8059};
  wire [2:0] _28792 = {_0, _28790} + {_0, _28791};
  wire [1:0] _28793 = {_0, _8991} + {_0, _10685};
  wire [3:0] _28794 = {_0, _28792} + {_0, _0, _28793};
  wire _28795 = _12301 < _28794;
  wire _28796 = r215 ^ _28795;
  wire _28797 = _12298 ? coded_block[215] : r215;
  wire _28798 = _12296 ? _28796 : _28797;
  always @ (posedge reset or posedge clock) if (reset) r215 <= 1'd0; else if (_12300) r215 <= _28798;
  wire [1:0] _28799 = {_0, _383} + {_0, _3294};
  wire [1:0] _28800 = {_0, _4256} + {_0, _6397};
  wire [2:0] _28801 = {_0, _28799} + {_0, _28800};
  wire [1:0] _28802 = {_0, _9917} + {_0, _12219};
  wire [3:0] _28803 = {_0, _28801} + {_0, _0, _28802};
  wire _28804 = _12301 < _28803;
  wire _28805 = r214 ^ _28804;
  wire _28806 = _12298 ? coded_block[214] : r214;
  wire _28807 = _12296 ? _28805 : _28806;
  always @ (posedge reset or posedge clock) if (reset) r214 <= 1'd0; else if (_12300) r214 <= _28807;
  wire [1:0] _28808 = {_0, _416} + {_0, _3964};
  wire [1:0] _28809 = {_0, _5373} + {_0, _6334};
  wire [2:0] _28810 = {_0, _28808} + {_0, _28809};
  wire [1:0] _28811 = {_0, _8480} + {_0, _11996};
  wire [3:0] _28812 = {_0, _28810} + {_0, _0, _28811};
  wire _28813 = _12301 < _28812;
  wire _28814 = r213 ^ _28813;
  wire _28815 = _12298 ? coded_block[213] : r213;
  wire _28816 = _12296 ? _28814 : _28815;
  always @ (posedge reset or posedge clock) if (reset) r213 <= 1'd0; else if (_12300) r213 <= _28816;
  wire [1:0] _28817 = {_0, _447} + {_0, _3549};
  wire [1:0] _28818 = {_0, _6045} + {_0, _7454};
  wire [2:0] _28819 = {_0, _28817} + {_0, _28818};
  wire [1:0] _28820 = {_0, _8415} + {_0, _10558};
  wire [3:0] _28821 = {_0, _28819} + {_0, _0, _28820};
  wire _28822 = _12301 < _28821;
  wire _28823 = r212 ^ _28822;
  wire _28824 = _12298 ? coded_block[212] : r212;
  wire _28825 = _12296 ? _28823 : _28824;
  always @ (posedge reset or posedge clock) if (reset) r212 <= 1'd0; else if (_12300) r212 <= _28825;
  wire [1:0] _28826 = {_0, _479} + {_0, _3262};
  wire [1:0] _28827 = {_0, _5628} + {_0, _8123};
  wire [2:0] _28828 = {_0, _28826} + {_0, _28827};
  wire [1:0] _28829 = {_0, _9534} + {_0, _10493};
  wire [3:0] _28830 = {_0, _28828} + {_0, _0, _28829};
  wire _28831 = _12301 < _28830;
  wire _28832 = r211 ^ _28831;
  wire _28833 = _12298 ? coded_block[211] : r211;
  wire _28834 = _12296 ? _28832 : _28833;
  always @ (posedge reset or posedge clock) if (reset) r211 <= 1'd0; else if (_12300) r211 <= _28834;
  wire [1:0] _28835 = {_0, _510} + {_0, _2208};
  wire [1:0] _28836 = {_0, _5342} + {_0, _7710};
  wire [2:0] _28837 = {_0, _28835} + {_0, _28836};
  wire [1:0] _28838 = {_0, _10204} + {_0, _11613};
  wire [3:0] _28839 = {_0, _28837} + {_0, _0, _28838};
  wire _28840 = _12301 < _28839;
  wire _28841 = r210 ^ _28840;
  wire _28842 = _12298 ? coded_block[210] : r210;
  wire _28843 = _12296 ? _28841 : _28842;
  always @ (posedge reset or posedge clock) if (reset) r210 <= 1'd0; else if (_12300) r210 <= _28843;
  wire [1:0] _28844 = {_0, _545} + {_0, _3709};
  wire [1:0] _28845 = {_0, _4287} + {_0, _7420};
  wire [2:0] _28846 = {_0, _28844} + {_0, _28845};
  wire [1:0] _28847 = {_0, _9790} + {_0, _12282};
  wire [3:0] _28848 = {_0, _28846} + {_0, _0, _28847};
  wire _28849 = _12301 < _28848;
  wire _28850 = r209 ^ _28849;
  wire _28851 = _12298 ? coded_block[209] : r209;
  wire _28852 = _12296 ? _28850 : _28851;
  always @ (posedge reset or posedge clock) if (reset) r209 <= 1'd0; else if (_12300) r209 <= _28852;
  wire [1:0] _28853 = {_0, _576} + {_0, _2686};
  wire [1:0] _28854 = {_0, _5790} + {_0, _6366};
  wire [2:0] _28855 = {_0, _28853} + {_0, _28854};
  wire [1:0] _28856 = {_0, _9503} + {_0, _11869};
  wire [3:0] _28857 = {_0, _28855} + {_0, _0, _28856};
  wire _28858 = _12301 < _28857;
  wire _28859 = r208 ^ _28858;
  wire _28860 = _12298 ? coded_block[208] : r208;
  wire _28861 = _12296 ? _28859 : _28860;
  always @ (posedge reset or posedge clock) if (reset) r208 <= 1'd0; else if (_12300) r208 <= _28861;
  wire [1:0] _28862 = {_0, _608} + {_0, _3453};
  wire [1:0] _28863 = {_0, _4767} + {_0, _7868};
  wire [2:0] _28864 = {_0, _28862} + {_0, _28863};
  wire [1:0] _28865 = {_0, _8446} + {_0, _11581};
  wire [3:0] _28866 = {_0, _28864} + {_0, _0, _28865};
  wire _28867 = _12301 < _28866;
  wire _28868 = r207 ^ _28867;
  wire _28869 = _12298 ? coded_block[207] : r207;
  wire _28870 = _12296 ? _28868 : _28869;
  always @ (posedge reset or posedge clock) if (reset) r207 <= 1'd0; else if (_12300) r207 <= _28870;
  wire [1:0] _28871 = {_0, _703} + {_0, _2271};
  wire [1:0] _28872 = {_0, _4223} + {_0, _6781};
  wire [2:0] _28873 = {_0, _28871} + {_0, _28872};
  wire [1:0] _28874 = {_0, _9693} + {_0, _11004};
  wire [3:0] _28875 = {_0, _28873} + {_0, _0, _28874};
  wire _28876 = _12301 < _28875;
  wire _28877 = r206 ^ _28876;
  wire _28878 = _12298 ? coded_block[206] : r206;
  wire _28879 = _12296 ? _28877 : _28878;
  always @ (posedge reset or posedge clock) if (reset) r206 <= 1'd0; else if (_12300) r206 <= _28879;
  wire [1:0] _28880 = {_0, _735} + {_0, _3615};
  wire [1:0] _28881 = {_0, _4350} + {_0, _6303};
  wire [2:0] _28882 = {_0, _28880} + {_0, _28881};
  wire [1:0] _28883 = {_0, _8863} + {_0, _11771};
  wire [3:0] _28884 = {_0, _28882} + {_0, _0, _28883};
  wire _28885 = _12301 < _28884;
  wire _28886 = r205 ^ _28885;
  wire _28887 = _12298 ? coded_block[205] : r205;
  wire _28888 = _12296 ? _28886 : _28887;
  always @ (posedge reset or posedge clock) if (reset) r205 <= 1'd0; else if (_12300) r205 <= _28888;
  wire [1:0] _28889 = {_0, _766} + {_0, _2847};
  wire [1:0] _28890 = {_0, _5694} + {_0, _6431};
  wire [2:0] _28891 = {_0, _28889} + {_0, _28890};
  wire [1:0] _28892 = {_0, _8383} + {_0, _10941};
  wire [3:0] _28893 = {_0, _28891} + {_0, _0, _28892};
  wire _28894 = _12301 < _28893;
  wire _28895 = r204 ^ _28894;
  wire _28896 = _12298 ? coded_block[204] : r204;
  wire _28897 = _12296 ? _28895 : _28896;
  always @ (posedge reset or posedge clock) if (reset) r204 <= 1'd0; else if (_12300) r204 <= _28897;
  wire [1:0] _28898 = {_0, _800} + {_0, _2813};
  wire [1:0] _28899 = {_0, _4926} + {_0, _7773};
  wire [2:0] _28900 = {_0, _28898} + {_0, _28899};
  wire [1:0] _28901 = {_0, _8511} + {_0, _10462};
  wire [3:0] _28902 = {_0, _28900} + {_0, _0, _28901};
  wire _28903 = _12301 < _28902;
  wire _28904 = r203 ^ _28903;
  wire _28905 = _12298 ? coded_block[203] : r203;
  wire _28906 = _12296 ? _28904 : _28905;
  always @ (posedge reset or posedge clock) if (reset) r203 <= 1'd0; else if (_12300) r203 <= _28906;
  wire [1:0] _28907 = {_0, _831} + {_0, _3646};
  wire [1:0] _28908 = {_0, _4895} + {_0, _7005};
  wire [2:0] _28909 = {_0, _28907} + {_0, _28908};
  wire [1:0] _28910 = {_0, _9853} + {_0, _10590};
  wire [3:0] _28911 = {_0, _28909} + {_0, _0, _28910};
  wire _28912 = _12301 < _28911;
  wire _28913 = r202 ^ _28912;
  wire _28914 = _12298 ? coded_block[202] : r202;
  wire _28915 = _12296 ? _28913 : _28914;
  always @ (posedge reset or posedge clock) if (reset) r202 <= 1'd0; else if (_12300) r202 <= _28915;
  wire [1:0] _28916 = {_0, _863} + {_0, _3933};
  wire [1:0] _28917 = {_0, _5726} + {_0, _6973};
  wire [2:0] _28918 = {_0, _28916} + {_0, _28917};
  wire [1:0] _28919 = {_0, _9085} + {_0, _11933};
  wire [3:0] _28920 = {_0, _28918} + {_0, _0, _28919};
  wire _28921 = _12301 < _28920;
  wire _28922 = r201 ^ _28921;
  wire _28923 = _12298 ? coded_block[201] : r201;
  wire _28924 = _12296 ? _28922 : _28923;
  always @ (posedge reset or posedge clock) if (reset) r201 <= 1'd0; else if (_12300) r201 <= _28924;
  wire [1:0] _28925 = {_0, _894} + {_0, _3325};
  wire [1:0] _28926 = {_0, _6012} + {_0, _7804};
  wire [2:0] _28927 = {_0, _28925} + {_0, _28926};
  wire [1:0] _28928 = {_0, _9054} + {_0, _11165};
  wire [3:0] _28929 = {_0, _28927} + {_0, _0, _28928};
  wire _28930 = _12301 < _28929;
  wire _28931 = r200 ^ _28930;
  wire _28932 = _12298 ? coded_block[200] : r200;
  wire _28933 = _12296 ? _28931 : _28932;
  always @ (posedge reset or posedge clock) if (reset) r200 <= 1'd0; else if (_12300) r200 <= _28933;
  wire [1:0] _28934 = {_0, _927} + {_0, _3167};
  wire [1:0] _28935 = {_0, _5407} + {_0, _8092};
  wire [2:0] _28936 = {_0, _28934} + {_0, _28935};
  wire [1:0] _28937 = {_0, _9886} + {_0, _11132};
  wire [3:0] _28938 = {_0, _28936} + {_0, _0, _28937};
  wire _28939 = _12301 < _28938;
  wire _28940 = r199 ^ _28939;
  wire _28941 = _12298 ? coded_block[199] : r199;
  wire _28942 = _12296 ? _28940 : _28941;
  always @ (posedge reset or posedge clock) if (reset) r199 <= 1'd0; else if (_12300) r199 <= _28942;
  wire [1:0] _28943 = {_0, _990} + {_0, _3198};
  wire [1:0] _28944 = {_0, _4129} + {_0, _7326};
  wire [2:0] _28945 = {_0, _28943} + {_0, _28944};
  wire [1:0] _28946 = {_0, _9566} + {_0, _12251};
  wire [3:0] _28947 = {_0, _28945} + {_0, _0, _28946};
  wire _28948 = _12301 < _28947;
  wire _28949 = r198 ^ _28948;
  wire _28950 = _12298 ? coded_block[198] : r198;
  wire _28951 = _12296 ? _28949 : _28950;
  always @ (posedge reset or posedge clock) if (reset) r198 <= 1'd0; else if (_12300) r198 <= _28951;
  wire [1:0] _28952 = {_0, _1021} + {_0, _3390};
  wire [1:0] _28953 = {_0, _5279} + {_0, _6176};
  wire [2:0] _28954 = {_0, _28952} + {_0, _28953};
  wire [1:0] _28955 = {_0, _9406} + {_0, _11644};
  wire [3:0] _28956 = {_0, _28954} + {_0, _0, _28955};
  wire _28957 = _12301 < _28956;
  wire _28958 = r197 ^ _28957;
  wire _28959 = _12298 ? coded_block[197] : r197;
  wire _28960 = _12296 ? _28958 : _28959;
  always @ (posedge reset or posedge clock) if (reset) r197 <= 1'd0; else if (_12300) r197 <= _28960;
  wire [1:0] _28961 = {_0, _1088} + {_0, _3773};
  wire [1:0] _28962 = {_0, _6108} + {_0, _7548};
  wire [2:0] _28963 = {_0, _28961} + {_0, _28962};
  wire [1:0] _28964 = {_0, _9438} + {_0, _10272};
  wire [3:0] _28965 = {_0, _28963} + {_0, _0, _28964};
  wire _28966 = _12301 < _28965;
  wire _28967 = r196 ^ _28966;
  wire _28968 = _12298 ? coded_block[196] : r196;
  wire _28969 = _12296 ? _28967 : _28968;
  always @ (posedge reset or posedge clock) if (reset) r196 <= 1'd0; else if (_12300) r196 <= _28969;
  wire [1:0] _28970 = {_0, _1120} + {_0, _2974};
  wire [1:0] _28971 = {_0, _5853} + {_0, _8186};
  wire [2:0] _28972 = {_0, _28970} + {_0, _28971};
  wire [1:0] _28973 = {_0, _9630} + {_0, _11516};
  wire [3:0] _28974 = {_0, _28972} + {_0, _0, _28973};
  wire _28975 = _12301 < _28974;
  wire _28976 = r195 ^ _28975;
  wire _28977 = _12298 ? coded_block[195] : r195;
  wire _28978 = _12296 ? _28976 : _28977;
  always @ (posedge reset or posedge clock) if (reset) r195 <= 1'd0; else if (_12300) r195 <= _28978;
  wire [1:0] _28979 = {_0, _1151} + {_0, _3037};
  wire [1:0] _28980 = {_0, _5053} + {_0, _7931};
  wire [2:0] _28981 = {_0, _28979} + {_0, _28980};
  wire [1:0] _28982 = {_0, _8256} + {_0, _11708};
  wire [3:0] _28983 = {_0, _28981} + {_0, _0, _28982};
  wire _28984 = _12301 < _28983;
  wire _28985 = r194 ^ _28984;
  wire _28986 = _12298 ? coded_block[194] : r194;
  wire _28987 = _12296 ? _28985 : _28986;
  always @ (posedge reset or posedge clock) if (reset) r194 <= 1'd0; else if (_12300) r194 <= _28987;
  wire [1:0] _28988 = {_0, _1215} + {_0, _2526};
  wire [1:0] _28989 = {_0, _5918} + {_0, _7199};
  wire [2:0] _28990 = {_0, _28988} + {_0, _28989};
  wire [1:0] _28991 = {_0, _9212} + {_0, _12092};
  wire [3:0] _28992 = {_0, _28990} + {_0, _0, _28991};
  wire _28993 = _12301 < _28992;
  wire _28994 = r193 ^ _28993;
  wire _28995 = _12298 ? coded_block[193] : r193;
  wire _28996 = _12296 ? _28994 : _28995;
  always @ (posedge reset or posedge clock) if (reset) r193 <= 1'd0; else if (_12300) r193 <= _28996;
  wire [1:0] _28997 = {_0, _1247} + {_0, _2430};
  wire [1:0] _28998 = {_0, _4605} + {_0, _7996};
  wire [2:0] _28999 = {_0, _28997} + {_0, _28998};
  wire [1:0] _29000 = {_0, _9279} + {_0, _11295};
  wire [3:0] _29001 = {_0, _28999} + {_0, _0, _29000};
  wire _29002 = _12301 < _29001;
  wire _29003 = r192 ^ _29002;
  wire _29004 = _12298 ? coded_block[192] : r192;
  wire _29005 = _12296 ? _29003 : _29004;
  always @ (posedge reset or posedge clock) if (reset) r192 <= 1'd0; else if (_12300) r192 <= _29005;
  wire [1:0] _29006 = {_0, _1278} + {_0, _2941};
  wire [1:0] _29007 = {_0, _4511} + {_0, _6687};
  wire [2:0] _29008 = {_0, _29006} + {_0, _29007};
  wire [1:0] _29009 = {_0, _10077} + {_0, _11358};
  wire [3:0] _29010 = {_0, _29008} + {_0, _0, _29009};
  wire _29011 = _12301 < _29010;
  wire _29012 = r191 ^ _29011;
  wire _29013 = _12298 ? coded_block[191] : r191;
  wire _29014 = _12296 ? _29012 : _29013;
  always @ (posedge reset or posedge clock) if (reset) r191 <= 1'd0; else if (_12300) r191 <= _29014;
  wire [1:0] _29015 = {_0, _1343} + {_0, _3068};
  wire [1:0] _29016 = {_0, _5884} + {_0, _7100};
  wire [2:0] _29017 = {_0, _29015} + {_0, _29016};
  wire [1:0] _29018 = {_0, _8670} + {_0, _10846};
  wire [3:0] _29019 = {_0, _29017} + {_0, _0, _29018};
  wire _29020 = _12301 < _29019;
  wire _29021 = r190 ^ _29020;
  wire _29022 = _12298 ? coded_block[190] : r190;
  wire _29023 = _12296 ? _29021 : _29022;
  always @ (posedge reset or posedge clock) if (reset) r190 <= 1'd0; else if (_12300) r190 <= _29023;
  wire [1:0] _29024 = {_0, _1375} + {_0, _2112};
  wire [1:0] _29025 = {_0, _5152} + {_0, _7965};
  wire [2:0] _29026 = {_0, _29024} + {_0, _29025};
  wire [1:0] _29027 = {_0, _9181} + {_0, _10748};
  wire [3:0] _29028 = {_0, _29026} + {_0, _0, _29027};
  wire _29029 = _12301 < _29028;
  wire _29030 = r189 ^ _29029;
  wire _29031 = _12298 ? coded_block[189] : r189;
  wire _29032 = _12296 ? _29030 : _29031;
  always @ (posedge reset or posedge clock) if (reset) r189 <= 1'd0; else if (_12300) r189 <= _29032;
  wire [1:0] _29033 = {_0, _1406} + {_0, _2655};
  wire [1:0] _29034 = {_0, _4192} + {_0, _7230};
  wire [2:0] _29035 = {_0, _29033} + {_0, _29034};
  wire [1:0] _29036 = {_0, _10045} + {_0, _11259};
  wire [3:0] _29037 = {_0, _29035} + {_0, _0, _29036};
  wire _29038 = _12301 < _29037;
  wire _29039 = r188 ^ _29038;
  wire _29040 = _12298 ? coded_block[188] : r188;
  wire _29041 = _12296 ? _29039 : _29040;
  always @ (posedge reset or posedge clock) if (reset) r188 <= 1'd0; else if (_12300) r188 <= _29041;
  wire [1:0] _29042 = {_0, _1439} + {_0, _3742};
  wire [1:0] _29043 = {_0, _4734} + {_0, _6270};
  wire [2:0] _29044 = {_0, _29042} + {_0, _29043};
  wire [1:0] _29045 = {_0, _9311} + {_0, _12124};
  wire [3:0] _29046 = {_0, _29044} + {_0, _0, _29045};
  wire _29047 = _12301 < _29046;
  wire _29048 = r187 ^ _29047;
  wire _29049 = _12298 ? coded_block[187] : r187;
  wire _29050 = _12296 ? _29048 : _29049;
  always @ (posedge reset or posedge clock) if (reset) r187 <= 1'd0; else if (_12300) r187 <= _29050;
  wire [1:0] _29051 = {_0, _1470} + {_0, _4060};
  wire [1:0] _29052 = {_0, _5821} + {_0, _6814};
  wire [2:0] _29053 = {_0, _29051} + {_0, _29052};
  wire [1:0] _29054 = {_0, _8352} + {_0, _11389};
  wire [3:0] _29055 = {_0, _29053} + {_0, _0, _29054};
  wire _29056 = _12301 < _29055;
  wire _29057 = r186 ^ _29056;
  wire _29058 = _12298 ? coded_block[186] : r186;
  wire _29059 = _12296 ? _29057 : _29058;
  always @ (posedge reset or posedge clock) if (reset) r186 <= 1'd0; else if (_12300) r186 <= _29059;
  wire [1:0] _29060 = {_0, _1502} + {_0, _2494};
  wire [1:0] _29061 = {_0, _6139} + {_0, _7900};
  wire [2:0] _29062 = {_0, _29060} + {_0, _29061};
  wire [1:0] _29063 = {_0, _8894} + {_0, _10430};
  wire [3:0] _29064 = {_0, _29062} + {_0, _0, _29063};
  wire _29065 = _12301 < _29064;
  wire _29066 = r185 ^ _29065;
  wire _29067 = _12298 ? coded_block[185] : r185;
  wire _29068 = _12296 ? _29066 : _29067;
  always @ (posedge reset or posedge clock) if (reset) r185 <= 1'd0; else if (_12300) r185 <= _29068;
  wire [1:0] _29069 = {_0, _1599} + {_0, _2878};
  wire [1:0] _29070 = {_0, _4861} + {_0, _8028};
  wire [2:0] _29071 = {_0, _29069} + {_0, _29070};
  wire [1:0] _29072 = {_0, _8736} + {_0, _10366};
  wire [3:0] _29073 = {_0, _29071} + {_0, _0, _29072};
  wire _29074 = _12301 < _29073;
  wire _29075 = r184 ^ _29074;
  wire _29076 = _12298 ? coded_block[184] : r184;
  wire _29077 = _12296 ? _29075 : _29076;
  always @ (posedge reset or posedge clock) if (reset) r184 <= 1'd0; else if (_12300) r184 <= _29077;
  wire [1:0] _29078 = {_0, _1631} + {_0, _2336};
  wire [1:0] _29079 = {_0, _4958} + {_0, _6942};
  wire [2:0] _29080 = {_0, _29078} + {_0, _29079};
  wire [1:0] _29081 = {_0, _10108} + {_0, _10814};
  wire [3:0] _29082 = {_0, _29080} + {_0, _0, _29081};
  wire _29083 = _12301 < _29082;
  wire _29084 = r183 ^ _29083;
  wire _29085 = _12298 ? coded_block[183] : r183;
  wire _29086 = _12296 ? _29084 : _29085;
  always @ (posedge reset or posedge clock) if (reset) r183 <= 1'd0; else if (_12300) r183 <= _29086;
  wire [1:0] _29087 = {_0, _1662} + {_0, _2592};
  wire [1:0] _29088 = {_0, _4415} + {_0, _7036};
  wire [2:0] _29089 = {_0, _29087} + {_0, _29088};
  wire [1:0] _29090 = {_0, _9022} + {_0, _12188};
  wire [3:0] _29091 = {_0, _29089} + {_0, _0, _29090};
  wire _29092 = _12301 < _29091;
  wire _29093 = r182 ^ _29092;
  wire _29094 = _12298 ? coded_block[182] : r182;
  wire _29095 = _12296 ? _29093 : _29094;
  always @ (posedge reset or posedge clock) if (reset) r182 <= 1'd0; else if (_12300) r182 <= _29095;
  wire [1:0] _29096 = {_0, _1695} + {_0, _3486};
  wire [1:0] _29097 = {_0, _4671} + {_0, _6494};
  wire [2:0] _29098 = {_0, _29096} + {_0, _29097};
  wire [1:0] _29099 = {_0, _9118} + {_0, _11101};
  wire [3:0] _29100 = {_0, _29098} + {_0, _0, _29099};
  wire _29101 = _12301 < _29100;
  wire _29102 = r181 ^ _29101;
  wire _29103 = _12298 ? coded_block[181] : r181;
  wire _29104 = _12296 ? _29102 : _29103;
  always @ (posedge reset or posedge clock) if (reset) r181 <= 1'd0; else if (_12300) r181 <= _29104;
  wire [1:0] _29105 = {_0, _1726} + {_0, _3135};
  wire [1:0] _29106 = {_0, _5565} + {_0, _6750};
  wire [2:0] _29107 = {_0, _29105} + {_0, _29106};
  wire [1:0] _29108 = {_0, _8574} + {_0, _11196};
  wire [3:0] _29109 = {_0, _29107} + {_0, _0, _29108};
  wire _29110 = _12301 < _29109;
  wire _29111 = r180 ^ _29110;
  wire _29112 = _12298 ? coded_block[180] : r180;
  wire _29113 = _12296 ? _29111 : _29112;
  always @ (posedge reset or posedge clock) if (reset) r180 <= 1'd0; else if (_12300) r180 <= _29113;
  wire [1:0] _29114 = {_0, _1758} + {_0, _3359};
  wire [1:0] _29115 = {_0, _5215} + {_0, _7644};
  wire [2:0] _29116 = {_0, _29114} + {_0, _29115};
  wire [1:0] _29117 = {_0, _8830} + {_0, _10654};
  wire [3:0] _29118 = {_0, _29116} + {_0, _0, _29117};
  wire _29119 = _12301 < _29118;
  wire _29120 = r179 ^ _29119;
  wire _29121 = _12298 ? coded_block[179] : r179;
  wire _29122 = _12296 ? _29120 : _29121;
  always @ (posedge reset or posedge clock) if (reset) r179 <= 1'd0; else if (_12300) r179 <= _29122;
  wire [1:0] _29123 = {_0, _1789} + {_0, _3231};
  wire [1:0] _29124 = {_0, _5438} + {_0, _7293};
  wire [2:0] _29125 = {_0, _29123} + {_0, _29124};
  wire [1:0] _29126 = {_0, _9724} + {_0, _10910};
  wire [3:0] _29127 = {_0, _29125} + {_0, _0, _29126};
  wire _29128 = _12301 < _29127;
  wire _29129 = r178 ^ _29128;
  wire _29130 = _12298 ? coded_block[178] : r178;
  wire _29131 = _12296 ? _29129 : _29130;
  always @ (posedge reset or posedge clock) if (reset) r178 <= 1'd0; else if (_12300) r178 <= _29131;
  wire [1:0] _29132 = {_0, _1823} + {_0, _3580};
  wire [1:0] _29133 = {_0, _5310} + {_0, _7517};
  wire [2:0] _29134 = {_0, _29132} + {_0, _29133};
  wire [1:0] _29135 = {_0, _9375} + {_0, _11806};
  wire [3:0] _29136 = {_0, _29134} + {_0, _0, _29135};
  wire _29137 = _12301 < _29136;
  wire _29138 = r177 ^ _29137;
  wire _29139 = _12298 ? coded_block[177] : r177;
  wire _29140 = _12296 ? _29138 : _29139;
  always @ (posedge reset or posedge clock) if (reset) r177 <= 1'd0; else if (_12300) r177 <= _29140;
  wire [1:0] _29141 = {_0, _1854} + {_0, _2302};
  wire [1:0] _29142 = {_0, _5663} + {_0, _7389};
  wire [2:0] _29143 = {_0, _29141} + {_0, _29142};
  wire [1:0] _29144 = {_0, _9597} + {_0, _11453};
  wire [3:0] _29145 = {_0, _29143} + {_0, _0, _29144};
  wire _29146 = _12301 < _29145;
  wire _29147 = r176 ^ _29146;
  wire _29148 = _12298 ? coded_block[176] : r176;
  wire _29149 = _12296 ? _29147 : _29148;
  always @ (posedge reset or posedge clock) if (reset) r176 <= 1'd0; else if (_12300) r176 <= _29149;
  wire [1:0] _29150 = {_0, _1886} + {_0, _2910};
  wire [1:0] _29151 = {_0, _4384} + {_0, _7741};
  wire [2:0] _29152 = {_0, _29150} + {_0, _29151};
  wire [1:0] _29153 = {_0, _9469} + {_0, _11677};
  wire [3:0] _29154 = {_0, _29152} + {_0, _0, _29153};
  wire _29155 = _12301 < _29154;
  wire _29156 = r175 ^ _29155;
  wire _29157 = _12298 ? coded_block[175] : r175;
  wire _29158 = _12296 ? _29156 : _29157;
  always @ (posedge reset or posedge clock) if (reset) r175 <= 1'd0; else if (_12300) r175 <= _29158;
  wire [1:0] _29159 = {_0, _1917} + {_0, _2463};
  wire [1:0] _29160 = {_0, _4989} + {_0, _6462};
  wire [2:0] _29161 = {_0, _29159} + {_0, _29160};
  wire [1:0] _29162 = {_0, _9822} + {_0, _11550};
  wire [3:0] _29163 = {_0, _29161} + {_0, _0, _29162};
  wire _29164 = _12301 < _29163;
  wire _29165 = r174 ^ _29164;
  wire _29166 = _12298 ? coded_block[174] : r174;
  wire _29167 = _12296 ? _29165 : _29166;
  always @ (posedge reset or posedge clock) if (reset) r174 <= 1'd0; else if (_12300) r174 <= _29167;
  wire [1:0] _29168 = {_0, _1950} + {_0, _4091};
  wire [1:0] _29169 = {_0, _4542} + {_0, _7069};
  wire [2:0] _29170 = {_0, _29168} + {_0, _29169};
  wire [1:0] _29171 = {_0, _8543} + {_0, _11900};
  wire [3:0] _29172 = {_0, _29170} + {_0, _0, _29171};
  wire _29173 = _12301 < _29172;
  wire _29174 = r173 ^ _29173;
  wire _29175 = _12298 ? coded_block[173] : r173;
  wire _29176 = _12296 ? _29174 : _29175;
  always @ (posedge reset or posedge clock) if (reset) r173 <= 1'd0; else if (_12300) r173 <= _29176;
  wire [1:0] _29177 = {_0, _1981} + {_0, _3104};
  wire [1:0] _29178 = {_0, _4160} + {_0, _6621};
  wire [2:0] _29179 = {_0, _29177} + {_0, _29178};
  wire [1:0] _29180 = {_0, _9149} + {_0, _10621};
  wire [3:0] _29181 = {_0, _29179} + {_0, _0, _29180};
  wire _29182 = _12301 < _29181;
  wire _29183 = r172 ^ _29182;
  wire _29184 = _12298 ? coded_block[172] : r172;
  wire _29185 = _12296 ? _29183 : _29184;
  always @ (posedge reset or posedge clock) if (reset) r172 <= 1'd0; else if (_12300) r172 <= _29185;
  wire [1:0] _29186 = {_0, _2013} + {_0, _3517};
  wire [1:0] _29187 = {_0, _5183} + {_0, _6239};
  wire [2:0] _29188 = {_0, _29186} + {_0, _29187};
  wire [1:0] _29189 = {_0, _8701} + {_0, _11228};
  wire [3:0] _29190 = {_0, _29188} + {_0, _0, _29189};
  wire _29191 = _12301 < _29190;
  wire _29192 = r171 ^ _29191;
  wire _29193 = _12298 ? coded_block[171] : r171;
  wire _29194 = _12296 ? _29192 : _29193;
  always @ (posedge reset or posedge clock) if (reset) r171 <= 1'd0; else if (_12300) r171 <= _29194;
  wire [1:0] _29195 = {_0, _34} + {_0, _2430};
  wire [1:0] _29196 = {_0, _4511} + {_0, _6589};
  wire [2:0] _29197 = {_0, _29195} + {_0, _29196};
  wire [1:0] _29198 = {_0, _8670} + {_0, _10748};
  wire [3:0] _29199 = {_0, _29197} + {_0, _0, _29198};
  wire _29200 = _12301 < _29199;
  wire _29201 = r170 ^ _29200;
  wire _29202 = _12298 ? coded_block[170] : r170;
  wire _29203 = _12296 ? _29201 : _29202;
  always @ (posedge reset or posedge clock) if (reset) r170 <= 1'd0; else if (_12300) r170 <= _29203;
  wire [1:0] _29204 = {_0, _1088} + {_0, _4028};
  wire [1:0] _29205 = {_0, _5853} + {_0, _6462};
  wire [2:0] _29206 = {_0, _29204} + {_0, _29205};
  wire [1:0] _29207 = {_0, _8446} + {_0, _11613};
  wire [3:0] _29208 = {_0, _29206} + {_0, _0, _29207};
  wire _29209 = _12301 < _29208;
  wire _29210 = r169 ^ _29209;
  wire _29211 = _12298 ? coded_block[169] : r169;
  wire _29212 = _12296 ? _29210 : _29211;
  always @ (posedge reset or posedge clock) if (reset) r169 <= 1'd0; else if (_12300) r169 <= _29212;
  wire [1:0] _29213 = {_0, _1120} + {_0, _2910};
  wire [1:0] _29214 = {_0, _6108} + {_0, _7931};
  wire [2:0] _29215 = {_0, _29213} + {_0, _29214};
  wire [1:0] _29216 = {_0, _8543} + {_0, _10527};
  wire [3:0] _29217 = {_0, _29215} + {_0, _0, _29216};
  wire _29218 = _12301 < _29217;
  wire _29219 = r168 ^ _29218;
  wire _29220 = _12298 ? coded_block[168] : r168;
  wire _29221 = _12296 ? _29219 : _29220;
  always @ (posedge reset or posedge clock) if (reset) r168 <= 1'd0; else if (_12300) r168 <= _29221;
  wire [1:0] _29222 = {_0, _1151} + {_0, _2557};
  wire [1:0] _29223 = {_0, _4989} + {_0, _8186};
  wire [2:0] _29224 = {_0, _29222} + {_0, _29223};
  wire [1:0] _29225 = {_0, _10014} + {_0, _10621};
  wire [3:0] _29226 = {_0, _29224} + {_0, _0, _29225};
  wire _29227 = _12301 < _29226;
  wire _29228 = r167 ^ _29227;
  wire _29229 = _12298 ? coded_block[167] : r167;
  wire _29230 = _12296 ? _29228 : _29229;
  always @ (posedge reset or posedge clock) if (reset) r167 <= 1'd0; else if (_12300) r167 <= _29230;
  wire [1:0] _29231 = {_0, _1184} + {_0, _2782};
  wire [1:0] _29232 = {_0, _4640} + {_0, _7069};
  wire [2:0] _29233 = {_0, _29231} + {_0, _29232};
  wire [1:0] _29234 = {_0, _8256} + {_0, _12092};
  wire [3:0] _29235 = {_0, _29233} + {_0, _0, _29234};
  wire _29236 = _12301 < _29235;
  wire _29237 = r166 ^ _29236;
  wire _29238 = _12298 ? coded_block[166] : r166;
  wire _29239 = _12296 ? _29237 : _29238;
  always @ (posedge reset or posedge clock) if (reset) r166 <= 1'd0; else if (_12300) r166 <= _29239;
  wire [1:0] _29240 = {_0, _1215} + {_0, _2655};
  wire [1:0] _29241 = {_0, _4861} + {_0, _6718};
  wire [2:0] _29242 = {_0, _29240} + {_0, _29241};
  wire [1:0] _29243 = {_0, _9149} + {_0, _10335};
  wire [3:0] _29244 = {_0, _29242} + {_0, _0, _29243};
  wire _29245 = _12301 < _29244;
  wire _29246 = r165 ^ _29245;
  wire _29247 = _12298 ? coded_block[165] : r165;
  wire _29248 = _12296 ? _29246 : _29247;
  always @ (posedge reset or posedge clock) if (reset) r165 <= 1'd0; else if (_12300) r165 <= _29248;
  wire [1:0] _29249 = {_0, _1247} + {_0, _3005};
  wire [1:0] _29250 = {_0, _4734} + {_0, _6942};
  wire [2:0] _29251 = {_0, _29249} + {_0, _29250};
  wire [1:0] _29252 = {_0, _8799} + {_0, _11228};
  wire [3:0] _29253 = {_0, _29251} + {_0, _0, _29252};
  wire _29254 = _12301 < _29253;
  wire _29255 = r164 ^ _29254;
  wire _29256 = _12298 ? coded_block[164] : r164;
  wire _29257 = _12296 ? _29255 : _29256;
  always @ (posedge reset or posedge clock) if (reset) r164 <= 1'd0; else if (_12300) r164 <= _29257;
  wire [1:0] _29258 = {_0, _1278} + {_0, _3742};
  wire [1:0] _29259 = {_0, _5085} + {_0, _6814};
  wire [2:0] _29260 = {_0, _29258} + {_0, _29259};
  wire [1:0] _29261 = {_0, _9022} + {_0, _10877};
  wire [3:0] _29262 = {_0, _29260} + {_0, _0, _29261};
  wire _29263 = _12301 < _29262;
  wire _29264 = r163 ^ _29263;
  wire _29265 = _12298 ? coded_block[163] : r163;
  wire _29266 = _12296 ? _29264 : _29265;
  always @ (posedge reset or posedge clock) if (reset) r163 <= 1'd0; else if (_12300) r163 <= _29266;
  wire [1:0] _29267 = {_0, _1312} + {_0, _2336};
  wire [1:0] _29268 = {_0, _5821} + {_0, _7163};
  wire [2:0] _29269 = {_0, _29267} + {_0, _29268};
  wire [1:0] _29270 = {_0, _8894} + {_0, _11101};
  wire [3:0] _29271 = {_0, _29269} + {_0, _0, _29270};
  wire _29272 = _12301 < _29271;
  wire _29273 = r162 ^ _29272;
  wire _29274 = _12298 ? coded_block[162] : r162;
  wire _29275 = _12296 ? _29273 : _29274;
  always @ (posedge reset or posedge clock) if (reset) r162 <= 1'd0; else if (_12300) r162 <= _29275;
  wire [1:0] _29276 = {_0, _1343} + {_0, _3901};
  wire [1:0] _29277 = {_0, _4415} + {_0, _7900};
  wire [2:0] _29278 = {_0, _29276} + {_0, _29277};
  wire [1:0] _29279 = {_0, _9248} + {_0, _10973};
  wire [3:0] _29280 = {_0, _29278} + {_0, _0, _29279};
  wire _29281 = _12301 < _29280;
  wire _29282 = r161 ^ _29281;
  wire _29283 = _12298 ? coded_block[161] : r161;
  wire _29284 = _12296 ? _29282 : _29283;
  always @ (posedge reset or posedge clock) if (reset) r161 <= 1'd0; else if (_12300) r161 <= _29284;
  wire [1:0] _29285 = {_0, _1375} + {_0, _3517};
  wire [1:0] _29286 = {_0, _5981} + {_0, _6494};
  wire [2:0] _29287 = {_0, _29285} + {_0, _29286};
  wire [1:0] _29288 = {_0, _9980} + {_0, _11326};
  wire [3:0] _29289 = {_0, _29287} + {_0, _0, _29288};
  wire _29290 = _12301 < _29289;
  wire _29291 = r160 ^ _29290;
  wire _29292 = _12298 ? coded_block[160] : r160;
  wire _29293 = _12296 ? _29291 : _29292;
  always @ (posedge reset or posedge clock) if (reset) r160 <= 1'd0; else if (_12300) r160 <= _29293;
  wire [1:0] _29294 = {_0, _1406} + {_0, _2526};
  wire [1:0] _29295 = {_0, _5597} + {_0, _8059};
  wire [2:0] _29296 = {_0, _29294} + {_0, _29295};
  wire [1:0] _29297 = {_0, _8574} + {_0, _12061};
  wire [3:0] _29298 = {_0, _29296} + {_0, _0, _29297};
  wire _29299 = _12301 < _29298;
  wire _29300 = r159 ^ _29299;
  wire _29301 = _12298 ? coded_block[159] : r159;
  wire _29302 = _12296 ? _29300 : _29301;
  always @ (posedge reset or posedge clock) if (reset) r159 <= 1'd0; else if (_12300) r159 <= _29302;
  wire [1:0] _29303 = {_0, _1439} + {_0, _2941};
  wire [1:0] _29304 = {_0, _4605} + {_0, _7675};
  wire [2:0] _29305 = {_0, _29303} + {_0, _29304};
  wire [1:0] _29306 = {_0, _10141} + {_0, _10654};
  wire [3:0] _29307 = {_0, _29305} + {_0, _0, _29306};
  wire _29308 = _12301 < _29307;
  wire _29309 = r158 ^ _29308;
  wire _29310 = _12298 ? coded_block[158] : r158;
  wire _29311 = _12296 ? _29309 : _29310;
  always @ (posedge reset or posedge clock) if (reset) r158 <= 1'd0; else if (_12300) r158 <= _29311;
  wire [1:0] _29312 = {_0, _1470} + {_0, _3422};
  wire [1:0] _29313 = {_0, _5022} + {_0, _6687};
  wire [2:0] _29314 = {_0, _29312} + {_0, _29313};
  wire [1:0] _29315 = {_0, _9759} + {_0, _12219};
  wire [3:0] _29316 = {_0, _29314} + {_0, _0, _29315};
  wire _29317 = _12301 < _29316;
  wire _29318 = r157 ^ _29317;
  wire _29319 = _12298 ? coded_block[157] : r157;
  wire _29320 = _12296 ? _29318 : _29319;
  always @ (posedge reset or posedge clock) if (reset) r157 <= 1'd0; else if (_12300) r157 <= _29320;
  wire [1:0] _29321 = {_0, _1502} + {_0, _2847};
  wire [1:0] _29322 = {_0, _5501} + {_0, _7100};
  wire [2:0] _29323 = {_0, _29321} + {_0, _29322};
  wire [1:0] _29324 = {_0, _8767} + {_0, _11837};
  wire [3:0] _29325 = {_0, _29323} + {_0, _0, _29324};
  wire _29326 = _12301 < _29325;
  wire _29327 = r156 ^ _29326;
  wire _29328 = _12298 ? coded_block[156] : r156;
  wire _29329 = _12296 ? _29327 : _29328;
  always @ (posedge reset or posedge clock) if (reset) r156 <= 1'd0; else if (_12300) r156 <= _29329;
  wire [1:0] _29330 = {_0, _1533} + {_0, _2144};
  wire [1:0] _29331 = {_0, _4926} + {_0, _7581};
  wire [2:0] _29332 = {_0, _29330} + {_0, _29331};
  wire [1:0] _29333 = {_0, _9181} + {_0, _10846};
  wire [3:0] _29334 = {_0, _29332} + {_0, _0, _29333};
  wire _29335 = _12301 < _29334;
  wire _29336 = r155 ^ _29335;
  wire _29337 = _12298 ? coded_block[155] : r155;
  wire _29338 = _12296 ? _29336 : _29337;
  always @ (posedge reset or posedge clock) if (reset) r155 <= 1'd0; else if (_12300) r155 <= _29338;
  wire [1:0] _29339 = {_0, _1568} + {_0, _3836};
  wire [1:0] _29340 = {_0, _4223} + {_0, _7005};
  wire [2:0] _29341 = {_0, _29339} + {_0, _29340};
  wire [1:0] _29342 = {_0, _9661} + {_0, _11259};
  wire [3:0] _29343 = {_0, _29341} + {_0, _0, _29342};
  wire _29344 = _12301 < _29343;
  wire _29345 = r154 ^ _29344;
  wire _29346 = _12298 ? coded_block[154] : r154;
  wire _29347 = _12296 ? _29345 : _29346;
  always @ (posedge reset or posedge clock) if (reset) r154 <= 1'd0; else if (_12300) r154 <= _29347;
  wire [1:0] _29348 = {_0, _1599} + {_0, _3997};
  wire [1:0] _29349 = {_0, _5918} + {_0, _6303};
  wire [2:0] _29350 = {_0, _29348} + {_0, _29349};
  wire [1:0] _29351 = {_0, _9085} + {_0, _11740};
  wire [3:0] _29352 = {_0, _29350} + {_0, _0, _29351};
  wire _29353 = _12301 < _29352;
  wire _29354 = r153 ^ _29353;
  wire _29355 = _12298 ? coded_block[153] : r153;
  wire _29356 = _12296 ? _29354 : _29355;
  always @ (posedge reset or posedge clock) if (reset) r153 <= 1'd0; else if (_12300) r153 <= _29356;
  wire [1:0] _29357 = {_0, _1631} + {_0, _3805};
  wire [1:0] _29358 = {_0, _6076} + {_0, _7996};
  wire [2:0] _29359 = {_0, _29357} + {_0, _29358};
  wire [1:0] _29360 = {_0, _8383} + {_0, _11165};
  wire [3:0] _29361 = {_0, _29359} + {_0, _0, _29360};
  wire _29362 = _12301 < _29361;
  wire _29363 = r152 ^ _29362;
  wire _29364 = _12298 ? coded_block[152] : r152;
  wire _29365 = _12296 ? _29363 : _29364;
  always @ (posedge reset or posedge clock) if (reset) r152 <= 1'd0; else if (_12300) r152 <= _29365;
  wire [1:0] _29366 = {_0, _1695} + {_0, _3325};
  wire [1:0] _29367 = {_0, _4256} + {_0, _7965};
  wire [2:0] _29368 = {_0, _29366} + {_0, _29367};
  wire [1:0] _29369 = {_0, _10235} + {_0, _12155};
  wire [3:0] _29370 = {_0, _29368} + {_0, _0, _29369};
  wire _29371 = _12301 < _29370;
  wire _29372 = r151 ^ _29371;
  wire _29373 = _12298 ? coded_block[151] : r151;
  wire _29374 = _12296 ? _29372 : _29373;
  always @ (posedge reset or posedge clock) if (reset) r151 <= 1'd0; else if (_12300) r151 <= _29374;
  wire [1:0] _29375 = {_0, _1726} + {_0, _3104};
  wire [1:0] _29376 = {_0, _5407} + {_0, _6334};
  wire [2:0] _29377 = {_0, _29375} + {_0, _29376};
  wire [1:0] _29378 = {_0, _10045} + {_0, _10303};
  wire [3:0] _29379 = {_0, _29377} + {_0, _0, _29378};
  wire _29380 = _12301 < _29379;
  wire _29381 = r150 ^ _29380;
  wire _29382 = _12298 ? coded_block[150] : r150;
  wire _29383 = _12296 ? _29381 : _29382;
  always @ (posedge reset or posedge clock) if (reset) r150 <= 1'd0; else if (_12300) r150 <= _29383;
  wire [1:0] _29384 = {_0, _1758} + {_0, _3678};
  wire [1:0] _29385 = {_0, _5183} + {_0, _7485};
  wire [2:0] _29386 = {_0, _29384} + {_0, _29385};
  wire [1:0] _29387 = {_0, _8415} + {_0, _12124};
  wire [3:0] _29388 = {_0, _29386} + {_0, _0, _29387};
  wire _29389 = _12301 < _29388;
  wire _29390 = r149 ^ _29389;
  wire _29391 = _12298 ? coded_block[149] : r149;
  wire _29392 = _12296 ? _29390 : _29391;
  always @ (posedge reset or posedge clock) if (reset) r149 <= 1'd0; else if (_12300) r149 <= _29392;
  wire [1:0] _29393 = {_0, _1789} + {_0, _3615};
  wire [1:0] _29394 = {_0, _5757} + {_0, _7262};
  wire [2:0] _29395 = {_0, _29393} + {_0, _29394};
  wire [1:0] _29396 = {_0, _9566} + {_0, _10493};
  wire [3:0] _29397 = {_0, _29395} + {_0, _0, _29396};
  wire _29398 = _12301 < _29397;
  wire _29399 = r148 ^ _29398;
  wire _29400 = _12298 ? coded_block[148] : r148;
  wire _29401 = _12296 ? _29399 : _29400;
  always @ (posedge reset or posedge clock) if (reset) r148 <= 1'd0; else if (_12300) r148 <= _29401;
  wire [1:0] _29402 = {_0, _1823} + {_0, _2719};
  wire [1:0] _29403 = {_0, _5694} + {_0, _7837};
  wire [2:0] _29404 = {_0, _29402} + {_0, _29403};
  wire [1:0] _29405 = {_0, _9342} + {_0, _11644};
  wire [3:0] _29406 = {_0, _29404} + {_0, _0, _29405};
  wire _29407 = _12301 < _29406;
  wire _29408 = r147 ^ _29407;
  wire _29409 = _12298 ? coded_block[147] : r147;
  wire _29410 = _12296 ? _29408 : _29409;
  always @ (posedge reset or posedge clock) if (reset) r147 <= 1'd0; else if (_12300) r147 <= _29410;
  wire [1:0] _29411 = {_0, _1854} + {_0, _3390};
  wire [1:0] _29412 = {_0, _4798} + {_0, _7773};
  wire [2:0] _29413 = {_0, _29411} + {_0, _29412};
  wire [1:0] _29414 = {_0, _9917} + {_0, _11422};
  wire [3:0] _29415 = {_0, _29413} + {_0, _0, _29414};
  wire _29416 = _12301 < _29415;
  wire _29417 = r146 ^ _29416;
  wire _29418 = _12298 ? coded_block[146] : r146;
  wire _29419 = _12296 ? _29417 : _29418;
  always @ (posedge reset or posedge clock) if (reset) r146 <= 1'd0; else if (_12300) r146 <= _29419;
  wire [1:0] _29420 = {_0, _1886} + {_0, _2974};
  wire [1:0] _29421 = {_0, _5470} + {_0, _6877};
  wire [2:0] _29422 = {_0, _29420} + {_0, _29421};
  wire [1:0] _29423 = {_0, _9853} + {_0, _11996};
  wire [3:0] _29424 = {_0, _29422} + {_0, _0, _29423};
  wire _29425 = _12301 < _29424;
  wire _29426 = r145 ^ _29425;
  wire _29427 = _12298 ? coded_block[145] : r145;
  wire _29428 = _12296 ? _29426 : _29427;
  always @ (posedge reset or posedge clock) if (reset) r145 <= 1'd0; else if (_12300) r145 <= _29428;
  wire [1:0] _29429 = {_0, _1917} + {_0, _2686};
  wire [1:0] _29430 = {_0, _5053} + {_0, _7548};
  wire [2:0] _29431 = {_0, _29429} + {_0, _29430};
  wire [1:0] _29432 = {_0, _8957} + {_0, _11933};
  wire [3:0] _29433 = {_0, _29431} + {_0, _0, _29432};
  wire _29434 = _12301 < _29433;
  wire _29435 = r144 ^ _29434;
  wire _29436 = _12298 ? coded_block[144] : r144;
  wire _29437 = _12296 ? _29435 : _29436;
  always @ (posedge reset or posedge clock) if (reset) r144 <= 1'd0; else if (_12300) r144 <= _29437;
  wire [1:0] _29438 = {_0, _1950} + {_0, _3646};
  wire [1:0] _29439 = {_0, _4767} + {_0, _7132};
  wire [2:0] _29440 = {_0, _29438} + {_0, _29439};
  wire [1:0] _29441 = {_0, _9630} + {_0, _11038};
  wire [3:0] _29442 = {_0, _29440} + {_0, _0, _29441};
  wire _29443 = _12301 < _29442;
  wire _29444 = r143 ^ _29443;
  wire _29445 = _12298 ? coded_block[143] : r143;
  wire _29446 = _12296 ? _29444 : _29445;
  always @ (posedge reset or posedge clock) if (reset) r143 <= 1'd0; else if (_12300) r143 <= _29446;
  wire [1:0] _29447 = {_0, _1981} + {_0, _3135};
  wire [1:0] _29448 = {_0, _5726} + {_0, _6845};
  wire [2:0] _29449 = {_0, _29447} + {_0, _29448};
  wire [1:0] _29450 = {_0, _9212} + {_0, _11708};
  wire [3:0] _29451 = {_0, _29449} + {_0, _0, _29450};
  wire _29452 = _12301 < _29451;
  wire _29453 = r142 ^ _29452;
  wire _29454 = _12298 ? coded_block[142] : r142;
  wire _29455 = _12296 ? _29453 : _29454;
  always @ (posedge reset or posedge clock) if (reset) r142 <= 1'd0; else if (_12300) r142 <= _29455;
  wire [1:0] _29456 = {_0, _2013} + {_0, _2112};
  wire [1:0] _29457 = {_0, _5215} + {_0, _7804};
  wire [2:0] _29458 = {_0, _29456} + {_0, _29457};
  wire [1:0] _29459 = {_0, _8926} + {_0, _11295};
  wire [3:0] _29460 = {_0, _29458} + {_0, _0, _29459};
  wire _29461 = _12301 < _29460;
  wire _29462 = r141 ^ _29461;
  wire _29463 = _12298 ? coded_block[141] : r141;
  wire _29464 = _12296 ? _29462 : _29463;
  always @ (posedge reset or posedge clock) if (reset) r141 <= 1'd0; else if (_12300) r141 <= _29464;
  wire [1:0] _29465 = {_0, _2044} + {_0, _2878};
  wire [1:0] _29466 = {_0, _4192} + {_0, _7293};
  wire [2:0] _29467 = {_0, _29465} + {_0, _29466};
  wire [1:0] _29468 = {_0, _9886} + {_0, _11004};
  wire [3:0] _29469 = {_0, _29467} + {_0, _0, _29468};
  wire _29470 = _12301 < _29469;
  wire _29471 = r140 ^ _29470;
  wire _29472 = _12298 ? coded_block[140] : r140;
  wire _29473 = _12296 ? _29471 : _29472;
  always @ (posedge reset or posedge clock) if (reset) r140 <= 1'd0; else if (_12300) r140 <= _29473;
  wire [1:0] _29474 = {_0, _65} + {_0, _4060};
  wire [1:0] _29475 = {_0, _4958} + {_0, _6270};
  wire [2:0] _29476 = {_0, _29474} + {_0, _29475};
  wire [1:0] _29477 = {_0, _9375} + {_0, _11964};
  wire [3:0] _29478 = {_0, _29476} + {_0, _0, _29477};
  wire _29479 = _12301 < _29478;
  wire _29480 = r139 ^ _29479;
  wire _29481 = _12298 ? coded_block[139] : r139;
  wire _29482 = _12296 ? _29480 : _29481;
  always @ (posedge reset or posedge clock) if (reset) r139 <= 1'd0; else if (_12300) r139 <= _29482;
  wire [1:0] _29483 = {_0, _97} + {_0, _3580};
  wire [1:0] _29484 = {_0, _6139} + {_0, _7036};
  wire [2:0] _29485 = {_0, _29483} + {_0, _29484};
  wire [1:0] _29486 = {_0, _8352} + {_0, _11453};
  wire [3:0] _29487 = {_0, _29485} + {_0, _0, _29486};
  wire _29488 = _12301 < _29487;
  wire _29489 = r138 ^ _29488;
  wire _29490 = _12298 ? coded_block[138] : r138;
  wire _29491 = _12296 ? _29489 : _29490;
  always @ (posedge reset or posedge clock) if (reset) r138 <= 1'd0; else if (_12300) r138 <= _29491;
  wire [1:0] _29492 = {_0, _128} + {_0, _3709};
  wire [1:0] _29493 = {_0, _5663} + {_0, _6207};
  wire [2:0] _29494 = {_0, _29492} + {_0, _29493};
  wire [1:0] _29495 = {_0, _9118} + {_0, _10430};
  wire [3:0] _29496 = {_0, _29494} + {_0, _0, _29495};
  wire _29497 = _12301 < _29496;
  wire _29498 = r137 ^ _29497;
  wire _29499 = _12298 ? coded_block[137] : r137;
  wire _29500 = _12296 ? _29498 : _29499;
  always @ (posedge reset or posedge clock) if (reset) r137 <= 1'd0; else if (_12300) r137 <= _29500;
  wire [1:0] _29501 = {_0, _192} + {_0, _2271};
  wire [1:0] _29502 = {_0, _5116} + {_0, _7868};
  wire [2:0] _29503 = {_0, _29501} + {_0, _29502};
  wire [1:0] _29504 = {_0, _9822} + {_0, _10366};
  wire [3:0] _29505 = {_0, _29503} + {_0, _0, _29504};
  wire _29506 = _12301 < _29505;
  wire _29507 = r136 ^ _29506;
  wire _29508 = _12298 ? coded_block[136] : r136;
  wire _29509 = _12296 ? _29507 : _29508;
  always @ (posedge reset or posedge clock) if (reset) r136 <= 1'd0; else if (_12300) r136 <= _29509;
  wire [1:0] _29510 = {_0, _224} + {_0, _2239};
  wire [1:0] _29511 = {_0, _4350} + {_0, _7199};
  wire [2:0] _29512 = {_0, _29510} + {_0, _29511};
  wire [1:0] _29513 = {_0, _9949} + {_0, _11900};
  wire [3:0] _29514 = {_0, _29512} + {_0, _0, _29513};
  wire _29515 = _12301 < _29514;
  wire _29516 = r135 ^ _29515;
  wire _29517 = _12298 ? coded_block[135] : r135;
  wire _29518 = _12296 ? _29516 : _29517;
  always @ (posedge reset or posedge clock) if (reset) r135 <= 1'd0; else if (_12300) r135 <= _29518;
  wire [1:0] _29519 = {_0, _255} + {_0, _3068};
  wire [1:0] _29520 = {_0, _4319} + {_0, _6431};
  wire [2:0] _29521 = {_0, _29519} + {_0, _29520};
  wire [1:0] _29522 = {_0, _9279} + {_0, _12027};
  wire [3:0] _29523 = {_0, _29521} + {_0, _0, _29522};
  wire _29524 = _12301 < _29523;
  wire _29525 = r134 ^ _29524;
  wire _29526 = _12298 ? coded_block[134] : r134;
  wire _29527 = _12296 ? _29525 : _29526;
  always @ (posedge reset or posedge clock) if (reset) r134 <= 1'd0; else if (_12300) r134 <= _29527;
  wire [1:0] _29528 = {_0, _289} + {_0, _3359};
  wire [1:0] _29529 = {_0, _5152} + {_0, _6397};
  wire [2:0] _29530 = {_0, _29528} + {_0, _29529};
  wire [1:0] _29531 = {_0, _8511} + {_0, _11358};
  wire [3:0] _29532 = {_0, _29530} + {_0, _0, _29531};
  wire _29533 = _12301 < _29532;
  wire _29534 = r133 ^ _29533;
  wire _29535 = _12298 ? coded_block[133] : r133;
  wire _29536 = _12296 ? _29534 : _29535;
  always @ (posedge reset or posedge clock) if (reset) r133 <= 1'd0; else if (_12300) r133 <= _29536;
  wire [1:0] _29537 = {_0, _320} + {_0, _2750};
  wire [1:0] _29538 = {_0, _5438} + {_0, _7230};
  wire [2:0] _29539 = {_0, _29537} + {_0, _29538};
  wire [1:0] _29540 = {_0, _8480} + {_0, _10590};
  wire [3:0] _29541 = {_0, _29539} + {_0, _0, _29540};
  wire _29542 = _12301 < _29541;
  wire _29543 = r132 ^ _29542;
  wire _29544 = _12298 ? coded_block[132] : r132;
  wire _29545 = _12296 ? _29543 : _29544;
  always @ (posedge reset or posedge clock) if (reset) r132 <= 1'd0; else if (_12300) r132 <= _29545;
  wire [1:0] _29546 = {_0, _352} + {_0, _2592};
  wire [1:0] _29547 = {_0, _4830} + {_0, _7517};
  wire [2:0] _29548 = {_0, _29546} + {_0, _29547};
  wire [1:0] _29549 = {_0, _9311} + {_0, _10558};
  wire [3:0] _29550 = {_0, _29548} + {_0, _0, _29549};
  wire _29551 = _12301 < _29550;
  wire _29552 = r131 ^ _29551;
  wire _29553 = _12298 ? coded_block[131] : r131;
  wire _29554 = _12296 ? _29552 : _29553;
  always @ (posedge reset or posedge clock) if (reset) r131 <= 1'd0; else if (_12300) r131 <= _29554;
  wire [1:0] _29555 = {_0, _383} + {_0, _2081};
  wire [1:0] _29556 = {_0, _4671} + {_0, _6908};
  wire [2:0] _29557 = {_0, _29555} + {_0, _29556};
  wire [1:0] _29558 = {_0, _9597} + {_0, _11389};
  wire [3:0] _29559 = {_0, _29557} + {_0, _0, _29558};
  wire _29560 = _12301 < _29559;
  wire _29561 = r130 ^ _29560;
  wire _29562 = _12298 ? coded_block[130] : r130;
  wire _29563 = _12296 ? _29561 : _29562;
  always @ (posedge reset or posedge clock) if (reset) r130 <= 1'd0; else if (_12300) r130 <= _29563;
  wire [1:0] _29564 = {_0, _416} + {_0, _2623};
  wire [1:0] _29565 = {_0, _4129} + {_0, _6750};
  wire [2:0] _29566 = {_0, _29564} + {_0, _29565};
  wire [1:0] _29567 = {_0, _8991} + {_0, _11677};
  wire [3:0] _29568 = {_0, _29566} + {_0, _0, _29567};
  wire _29569 = _12301 < _29568;
  wire _29570 = r129 ^ _29569;
  wire _29571 = _12298 ? coded_block[129] : r129;
  wire _29572 = _12296 ? _29570 : _29571;
  always @ (posedge reset or posedge clock) if (reset) r129 <= 1'd0; else if (_12300) r129 <= _29572;
  wire [1:0] _29573 = {_0, _447} + {_0, _2813};
  wire [1:0] _29574 = {_0, _4703} + {_0, _6176};
  wire [2:0] _29575 = {_0, _29573} + {_0, _29574};
  wire [1:0] _29576 = {_0, _8830} + {_0, _11069};
  wire [3:0] _29577 = {_0, _29575} + {_0, _0, _29576};
  wire _29578 = _12301 < _29577;
  wire _29579 = r128 ^ _29578;
  wire _29580 = _12298 ? coded_block[128] : r128;
  wire _29581 = _12296 ? _29579 : _29580;
  always @ (posedge reset or posedge clock) if (reset) r128 <= 1'd0; else if (_12300) r128 <= _29581;
  wire [1:0] _29582 = {_0, _479} + {_0, _3453};
  wire [1:0] _29583 = {_0, _4895} + {_0, _6781};
  wire [2:0] _29584 = {_0, _29582} + {_0, _29583};
  wire [1:0] _29585 = {_0, _8225} + {_0, _10910};
  wire [3:0] _29586 = {_0, _29584} + {_0, _0, _29585};
  wire _29587 = _12301 < _29586;
  wire _29588 = r127 ^ _29587;
  wire _29589 = _12298 ? coded_block[127] : r127;
  wire _29590 = _12296 ? _29588 : _29589;
  always @ (posedge reset or posedge clock) if (reset) r127 <= 1'd0; else if (_12300) r127 <= _29590;
  wire [1:0] _29591 = {_0, _510} + {_0, _3198};
  wire [1:0] _29592 = {_0, _5534} + {_0, _6973};
  wire [2:0] _29593 = {_0, _29591} + {_0, _29592};
  wire [1:0] _29594 = {_0, _8863} + {_0, _10272};
  wire [3:0] _29595 = {_0, _29593} + {_0, _0, _29594};
  wire _29596 = _12301 < _29595;
  wire _29597 = r126 ^ _29596;
  wire _29598 = _12298 ? coded_block[126] : r126;
  wire _29599 = _12296 ? _29597 : _29598;
  always @ (posedge reset or posedge clock) if (reset) r126 <= 1'd0; else if (_12300) r126 <= _29599;
  wire [1:0] _29600 = {_0, _545} + {_0, _2399};
  wire [1:0] _29601 = {_0, _5279} + {_0, _7612};
  wire [2:0] _29602 = {_0, _29600} + {_0, _29601};
  wire [1:0] _29603 = {_0, _9054} + {_0, _10941};
  wire [3:0] _29604 = {_0, _29602} + {_0, _0, _29603};
  wire _29605 = _12301 < _29604;
  wire _29606 = r125 ^ _29605;
  wire _29607 = _12298 ? coded_block[125] : r125;
  wire _29608 = _12296 ? _29606 : _29607;
  always @ (posedge reset or posedge clock) if (reset) r125 <= 1'd0; else if (_12300) r125 <= _29608;
  wire [1:0] _29609 = {_0, _576} + {_0, _2463};
  wire [1:0] _29610 = {_0, _4478} + {_0, _7357};
  wire [2:0] _29611 = {_0, _29609} + {_0, _29610};
  wire [1:0] _29612 = {_0, _9693} + {_0, _11132};
  wire [3:0] _29613 = {_0, _29611} + {_0, _0, _29612};
  wire _29614 = _12301 < _29613;
  wire _29615 = r124 ^ _29614;
  wire _29616 = _12298 ? coded_block[124] : r124;
  wire _29617 = _12296 ? _29615 : _29616;
  always @ (posedge reset or posedge clock) if (reset) r124 <= 1'd0; else if (_12300) r124 <= _29617;
  wire [1:0] _29618 = {_0, _608} + {_0, _3262};
  wire [1:0] _29619 = {_0, _4542} + {_0, _6558};
  wire [2:0] _29620 = {_0, _29618} + {_0, _29619};
  wire [1:0] _29621 = {_0, _9438} + {_0, _11771};
  wire [3:0] _29622 = {_0, _29620} + {_0, _0, _29621};
  wire _29623 = _12301 < _29622;
  wire _29624 = r123 ^ _29623;
  wire _29625 = _12298 ? coded_block[123] : r123;
  wire _29626 = _12296 ? _29624 : _29625;
  always @ (posedge reset or posedge clock) if (reset) r123 <= 1'd0; else if (_12300) r123 <= _29626;
  wire [1:0] _29627 = {_0, _639} + {_0, _3964};
  wire [1:0] _29628 = {_0, _5342} + {_0, _6621};
  wire [2:0] _29629 = {_0, _29627} + {_0, _29628};
  wire [1:0] _29630 = {_0, _8638} + {_0, _11516};
  wire [3:0] _29631 = {_0, _29629} + {_0, _0, _29630};
  wire _29632 = _12301 < _29631;
  wire _29633 = r122 ^ _29632;
  wire _29634 = _12298 ? coded_block[122] : r122;
  wire _29635 = _12296 ? _29633 : _29634;
  always @ (posedge reset or posedge clock) if (reset) r122 <= 1'd0; else if (_12300) r122 <= _29635;
  wire [1:0] _29636 = {_0, _703} + {_0, _2367};
  wire [1:0] _29637 = {_0, _5949} + {_0, _8123};
  wire [2:0] _29638 = {_0, _29636} + {_0, _29637};
  wire [1:0] _29639 = {_0, _9503} + {_0, _10783};
  wire [3:0] _29640 = {_0, _29638} + {_0, _0, _29639};
  wire _29641 = _12301 < _29640;
  wire _29642 = r121 ^ _29641;
  wire _29643 = _12298 ? coded_block[121] : r121;
  wire _29644 = _12296 ? _29642 : _29643;
  always @ (posedge reset or posedge clock) if (reset) r121 <= 1'd0; else if (_12300) r121 <= _29644;
  wire [1:0] _29645 = {_0, _735} + {_0, _3231};
  wire [1:0] _29646 = {_0, _4447} + {_0, _8028};
  wire [2:0] _29647 = {_0, _29645} + {_0, _29646};
  wire [1:0] _29648 = {_0, _10204} + {_0, _11581};
  wire [3:0] _29649 = {_0, _29647} + {_0, _0, _29648};
  wire _29650 = _12301 < _29649;
  wire _29651 = r120 ^ _29650;
  wire _29652 = _12298 ? coded_block[120] : r120;
  wire _29653 = _12296 ? _29651 : _29652;
  always @ (posedge reset or posedge clock) if (reset) r120 <= 1'd0; else if (_12300) r120 <= _29653;
  wire [1:0] _29654 = {_0, _766} + {_0, _2494};
  wire [1:0] _29655 = {_0, _5310} + {_0, _6525};
  wire [2:0] _29656 = {_0, _29654} + {_0, _29655};
  wire [1:0] _29657 = {_0, _10108} + {_0, _12282};
  wire [3:0] _29658 = {_0, _29656} + {_0, _0, _29657};
  wire _29659 = _12301 < _29658;
  wire _29660 = r119 ^ _29659;
  wire _29661 = _12298 ? coded_block[119] : r119;
  wire _29662 = _12296 ? _29660 : _29661;
  always @ (posedge reset or posedge clock) if (reset) r119 <= 1'd0; else if (_12300) r119 <= _29662;
  wire [1:0] _29663 = {_0, _800} + {_0, _3549};
  wire [1:0] _29664 = {_0, _4574} + {_0, _7389};
  wire [2:0] _29665 = {_0, _29663} + {_0, _29664};
  wire [1:0] _29666 = {_0, _8607} + {_0, _12188};
  wire [3:0] _29667 = {_0, _29665} + {_0, _0, _29666};
  wire _29668 = _12301 < _29667;
  wire _29669 = r118 ^ _29668;
  wire _29670 = _12298 ? coded_block[118] : r118;
  wire _29671 = _12296 ? _29669 : _29670;
  always @ (posedge reset or posedge clock) if (reset) r118 <= 1'd0; else if (_12300) r118 <= _29671;
  wire [1:0] _29672 = {_0, _831} + {_0, _4091};
  wire [1:0] _29673 = {_0, _5628} + {_0, _6652};
  wire [2:0] _29674 = {_0, _29672} + {_0, _29673};
  wire [1:0] _29675 = {_0, _9469} + {_0, _10685};
  wire [3:0] _29676 = {_0, _29674} + {_0, _0, _29675};
  wire _29677 = _12301 < _29676;
  wire _29678 = r117 ^ _29677;
  wire _29679 = _12298 ? coded_block[117] : r117;
  wire _29680 = _12296 ? _29678 : _29679;
  always @ (posedge reset or posedge clock) if (reset) r117 <= 1'd0; else if (_12300) r117 <= _29680;
  wire [1:0] _29681 = {_0, _863} + {_0, _3167};
  wire [1:0] _29682 = {_0, _4160} + {_0, _7710};
  wire [2:0] _29683 = {_0, _29681} + {_0, _29682};
  wire [1:0] _29684 = {_0, _8736} + {_0, _11550};
  wire [3:0] _29685 = {_0, _29683} + {_0, _0, _29684};
  wire _29686 = _12301 < _29685;
  wire _29687 = r116 ^ _29686;
  wire _29688 = _12298 ? coded_block[116] : r116;
  wire _29689 = _12296 ? _29687 : _29688;
  always @ (posedge reset or posedge clock) if (reset) r116 <= 1'd0; else if (_12300) r116 <= _29689;
  wire [1:0] _29690 = {_0, _894} + {_0, _3486};
  wire [1:0] _29691 = {_0, _5246} + {_0, _6239};
  wire [2:0] _29692 = {_0, _29690} + {_0, _29691};
  wire [1:0] _29693 = {_0, _9790} + {_0, _10814};
  wire [3:0] _29694 = {_0, _29692} + {_0, _0, _29693};
  wire _29695 = _12301 < _29694;
  wire _29696 = r115 ^ _29695;
  wire _29697 = _12298 ? coded_block[115] : r115;
  wire _29698 = _12296 ? _29696 : _29697;
  always @ (posedge reset or posedge clock) if (reset) r115 <= 1'd0; else if (_12300) r115 <= _29698;
  wire [1:0] _29699 = {_0, _927} + {_0, _3933};
  wire [1:0] _29700 = {_0, _5565} + {_0, _7326};
  wire [2:0] _29701 = {_0, _29699} + {_0, _29700};
  wire [1:0] _29702 = {_0, _8319} + {_0, _11869};
  wire [3:0] _29703 = {_0, _29701} + {_0, _0, _29702};
  wire _29704 = _12301 < _29703;
  wire _29705 = r114 ^ _29704;
  wire _29706 = _12298 ? coded_block[114] : r114;
  wire _29707 = _12296 ? _29705 : _29706;
  always @ (posedge reset or posedge clock) if (reset) r114 <= 1'd0; else if (_12300) r114 <= _29707;
  wire [1:0] _29708 = {_0, _958} + {_0, _3294};
  wire [1:0] _29709 = {_0, _6012} + {_0, _7644};
  wire [2:0] _29710 = {_0, _29708} + {_0, _29709};
  wire [1:0] _29711 = {_0, _9406} + {_0, _10399};
  wire [3:0] _29712 = {_0, _29710} + {_0, _0, _29711};
  wire _29713 = _12301 < _29712;
  wire _29714 = r113 ^ _29713;
  wire _29715 = _12298 ? coded_block[113] : r113;
  wire _29716 = _12296 ? _29714 : _29715;
  always @ (posedge reset or posedge clock) if (reset) r113 <= 1'd0; else if (_12300) r113 <= _29716;
  wire [1:0] _29717 = {_0, _990} + {_0, _2208};
  wire [1:0] _29718 = {_0, _5373} + {_0, _8092};
  wire [2:0] _29719 = {_0, _29717} + {_0, _29718};
  wire [1:0] _29720 = {_0, _9724} + {_0, _11485};
  wire [3:0] _29721 = {_0, _29719} + {_0, _0, _29720};
  wire _29722 = _12301 < _29721;
  wire _29723 = r112 ^ _29722;
  wire _29724 = _12298 ? coded_block[112] : r112;
  wire _29725 = _12296 ? _29723 : _29724;
  always @ (posedge reset or posedge clock) if (reset) r112 <= 1'd0; else if (_12300) r112 <= _29725;
  wire [1:0] _29726 = {_0, _1057} + {_0, _3773};
  wire [1:0] _29727 = {_0, _4384} + {_0, _6366};
  wire [2:0] _29728 = {_0, _29726} + {_0, _29727};
  wire [1:0] _29729 = {_0, _9534} + {_0, _12251};
  wire [3:0] _29730 = {_0, _29728} + {_0, _0, _29729};
  wire _29731 = _12301 < _29730;
  wire _29732 = r111 ^ _29731;
  wire _29733 = _12298 ? coded_block[111] : r111;
  wire _29734 = _12296 ? _29732 : _29733;
  always @ (posedge reset or posedge clock) if (reset) r111 <= 1'd0; else if (_12300) r111 <= _29734;
  wire [1:0] _29735 = {_0, _34} + {_0, _3453};
  wire [1:0] _29736 = {_0, _5534} + {_0, _7612};
  wire [2:0] _29737 = {_0, _29735} + {_0, _29736};
  wire [1:0] _29738 = {_0, _9693} + {_0, _11771};
  wire [3:0] _29739 = {_0, _29737} + {_0, _0, _29738};
  wire _29740 = _12301 < _29739;
  wire _29741 = r110 ^ _29740;
  wire _29742 = _12298 ? coded_block[110] : r110;
  wire _29743 = _12296 ? _29741 : _29742;
  always @ (posedge reset or posedge clock) if (reset) r110 <= 1'd0; else if (_12300) r110 <= _29743;
  wire [1:0] _29744 = {_0, _1406} + {_0, _2081};
  wire [1:0] _29745 = {_0, _5694} + {_0, _7931};
  wire [2:0] _29746 = {_0, _29744} + {_0, _29745};
  wire [1:0] _29747 = {_0, _8607} + {_0, _10399};
  wire [3:0] _29748 = {_0, _29746} + {_0, _0, _29747};
  wire _29749 = _12301 < _29748;
  wire _29750 = r109 ^ _29749;
  wire _29751 = _12298 ? coded_block[109] : r109;
  wire _29752 = _12296 ? _29750 : _29751;
  always @ (posedge reset or posedge clock) if (reset) r109 <= 1'd0; else if (_12300) r109 <= _29752;
  wire [1:0] _29753 = {_0, _1439} + {_0, _3646};
  wire [1:0] _29754 = {_0, _4129} + {_0, _7773};
  wire [2:0] _29755 = {_0, _29753} + {_0, _29754};
  wire [1:0] _29756 = {_0, _10014} + {_0, _10685};
  wire [3:0] _29757 = {_0, _29755} + {_0, _0, _29756};
  wire _29758 = _12301 < _29757;
  wire _29759 = r108 ^ _29758;
  wire _29760 = _12298 ? coded_block[108] : r108;
  wire _29761 = _12296 ? _29759 : _29760;
  always @ (posedge reset or posedge clock) if (reset) r108 <= 1'd0; else if (_12300) r108 <= _29761;
  wire [1:0] _29762 = {_0, _1470} + {_0, _3836};
  wire [1:0] _29763 = {_0, _5726} + {_0, _6176};
  wire [2:0] _29764 = {_0, _29762} + {_0, _29763};
  wire [1:0] _29765 = {_0, _9853} + {_0, _12092};
  wire [3:0] _29766 = {_0, _29764} + {_0, _0, _29765};
  wire _29767 = _12301 < _29766;
  wire _29768 = r107 ^ _29767;
  wire _29769 = _12298 ? coded_block[107] : r107;
  wire _29770 = _12296 ? _29768 : _29769;
  always @ (posedge reset or posedge clock) if (reset) r107 <= 1'd0; else if (_12300) r107 <= _29770;
  wire [1:0] _29771 = {_0, _1502} + {_0, _2463};
  wire [1:0] _29772 = {_0, _5918} + {_0, _7804};
  wire [2:0] _29773 = {_0, _29771} + {_0, _29772};
  wire [1:0] _29774 = {_0, _8225} + {_0, _11933};
  wire [3:0] _29775 = {_0, _29773} + {_0, _0, _29774};
  wire _29776 = _12301 < _29775;
  wire _29777 = r106 ^ _29776;
  wire _29778 = _12298 ? coded_block[106] : r106;
  wire _29779 = _12296 ? _29777 : _29778;
  always @ (posedge reset or posedge clock) if (reset) r106 <= 1'd0; else if (_12300) r106 <= _29779;
  wire [1:0] _29780 = {_0, _1599} + {_0, _3486};
  wire [1:0] _29781 = {_0, _5501} + {_0, _6366};
  wire [2:0] _29782 = {_0, _29780} + {_0, _29781};
  wire [1:0] _29783 = {_0, _8701} + {_0, _12155};
  wire [3:0] _29784 = {_0, _29782} + {_0, _0, _29783};
  wire _29785 = _12301 < _29784;
  wire _29786 = r105 ^ _29785;
  wire _29787 = _12298 ? coded_block[105] : r105;
  wire _29788 = _12296 ? _29786 : _29787;
  always @ (posedge reset or posedge clock) if (reset) r105 <= 1'd0; else if (_12300) r105 <= _29788;
  wire [1:0] _29789 = {_0, _1631} + {_0, _2271};
  wire [1:0] _29790 = {_0, _5565} + {_0, _7581};
  wire [2:0] _29791 = {_0, _29789} + {_0, _29790};
  wire [1:0] _29792 = {_0, _8446} + {_0, _10783};
  wire [3:0] _29793 = {_0, _29791} + {_0, _0, _29792};
  wire _29794 = _12301 < _29793;
  wire _29795 = r104 ^ _29794;
  wire _29796 = _12298 ? coded_block[104] : r104;
  wire _29797 = _12296 ? _29795 : _29796;
  always @ (posedge reset or posedge clock) if (reset) r104 <= 1'd0; else if (_12300) r104 <= _29797;
  wire [1:0] _29798 = {_0, _1662} + {_0, _2974};
  wire [1:0] _29799 = {_0, _4350} + {_0, _7644};
  wire [2:0] _29800 = {_0, _29798} + {_0, _29799};
  wire [1:0] _29801 = {_0, _9661} + {_0, _10527};
  wire [3:0] _29802 = {_0, _29800} + {_0, _0, _29801};
  wire _29803 = _12301 < _29802;
  wire _29804 = r103 ^ _29803;
  wire _29805 = _12298 ? coded_block[103] : r103;
  wire _29806 = _12296 ? _29804 : _29805;
  always @ (posedge reset or posedge clock) if (reset) r103 <= 1'd0; else if (_12300) r103 <= _29806;
  wire [1:0] _29807 = {_0, _1695} + {_0, _2878};
  wire [1:0] _29808 = {_0, _5053} + {_0, _6431};
  wire [2:0] _29809 = {_0, _29807} + {_0, _29808};
  wire [1:0] _29810 = {_0, _9724} + {_0, _11740};
  wire [3:0] _29811 = {_0, _29809} + {_0, _0, _29810};
  wire _29812 = _12301 < _29811;
  wire _29813 = r102 ^ _29812;
  wire _29814 = _12298 ? coded_block[102] : r102;
  wire _29815 = _12296 ? _29813 : _29814;
  always @ (posedge reset or posedge clock) if (reset) r102 <= 1'd0; else if (_12300) r102 <= _29815;
  wire [1:0] _29816 = {_0, _1758} + {_0, _2239};
  wire [1:0] _29817 = {_0, _5470} + {_0, _7036};
  wire [2:0] _29818 = {_0, _29816} + {_0, _29817};
  wire [1:0] _29819 = {_0, _9212} + {_0, _10590};
  wire [3:0] _29820 = {_0, _29818} + {_0, _0, _29819};
  wire _29821 = _12301 < _29820;
  wire _29822 = r101 ^ _29821;
  wire _29823 = _12298 ? coded_block[101] : r101;
  wire _29824 = _12296 ? _29822 : _29823;
  always @ (posedge reset or posedge clock) if (reset) r101 <= 1'd0; else if (_12300) r101 <= _29824;
  wire [1:0] _29825 = {_0, _1789} + {_0, _3517};
  wire [1:0] _29826 = {_0, _4319} + {_0, _7548};
  wire [2:0] _29827 = {_0, _29825} + {_0, _29826};
  wire [1:0] _29828 = {_0, _9118} + {_0, _11295};
  wire [3:0] _29829 = {_0, _29827} + {_0, _0, _29828};
  wire _29830 = _12301 < _29829;
  wire _29831 = r100 ^ _29830;
  wire _29832 = _12298 ? coded_block[100] : r100;
  wire _29833 = _12296 ? _29831 : _29832;
  always @ (posedge reset or posedge clock) if (reset) r100 <= 1'd0; else if (_12300) r100 <= _29833;
  wire [1:0] _29834 = {_0, _1823} + {_0, _2557};
  wire [1:0] _29835 = {_0, _5597} + {_0, _6397};
  wire [2:0] _29836 = {_0, _29834} + {_0, _29835};
  wire [1:0] _29837 = {_0, _9630} + {_0, _11196};
  wire [3:0] _29838 = {_0, _29836} + {_0, _0, _29837};
  wire _29839 = _12301 < _29838;
  wire _29840 = r99 ^ _29839;
  wire _29841 = _12298 ? coded_block[99] : r99;
  wire _29842 = _12296 ? _29840 : _29841;
  always @ (posedge reset or posedge clock) if (reset) r99 <= 1'd0; else if (_12300) r99 <= _29842;
  wire [1:0] _29843 = {_0, _1854} + {_0, _3104};
  wire [1:0] _29844 = {_0, _4640} + {_0, _7675};
  wire [2:0] _29845 = {_0, _29843} + {_0, _29844};
  wire [1:0] _29846 = {_0, _8480} + {_0, _11708};
  wire [3:0] _29847 = {_0, _29845} + {_0, _0, _29846};
  wire _29848 = _12301 < _29847;
  wire _29849 = r98 ^ _29848;
  wire _29850 = _12298 ? coded_block[98] : r98;
  wire _29851 = _12296 ? _29849 : _29850;
  always @ (posedge reset or posedge clock) if (reset) r98 <= 1'd0; else if (_12300) r98 <= _29851;
  wire [1:0] _29852 = {_0, _1886} + {_0, _2175};
  wire [1:0] _29853 = {_0, _5183} + {_0, _6718};
  wire [2:0] _29854 = {_0, _29852} + {_0, _29853};
  wire [1:0] _29855 = {_0, _9759} + {_0, _10558};
  wire [3:0] _29856 = {_0, _29854} + {_0, _0, _29855};
  wire _29857 = _12301 < _29856;
  wire _29858 = r97 ^ _29857;
  wire _29859 = _12298 ? coded_block[97] : r97;
  wire _29860 = _12296 ? _29858 : _29859;
  always @ (posedge reset or posedge clock) if (reset) r97 <= 1'd0; else if (_12300) r97 <= _29860;
  wire [1:0] _29861 = {_0, _1950} + {_0, _2941};
  wire [1:0] _29862 = {_0, _4574} + {_0, _6334};
  wire [2:0] _29863 = {_0, _29861} + {_0, _29862};
  wire [1:0] _29864 = {_0, _9342} + {_0, _10877};
  wire [3:0] _29865 = {_0, _29863} + {_0, _0, _29864};
  wire _29866 = _12301 < _29865;
  wire _29867 = r96 ^ _29866;
  wire _29868 = _12298 ? coded_block[96] : r96;
  wire _29869 = _12296 ? _29867 : _29868;
  always @ (posedge reset or posedge clock) if (reset) r96 <= 1'd0; else if (_12300) r96 <= _29869;
  wire [1:0] _29870 = {_0, _1981} + {_0, _2302};
  wire [1:0] _29871 = {_0, _5022} + {_0, _6652};
  wire [2:0] _29872 = {_0, _29870} + {_0, _29871};
  wire [1:0] _29873 = {_0, _8415} + {_0, _11422};
  wire [3:0] _29874 = {_0, _29872} + {_0, _0, _29873};
  wire _29875 = _12301 < _29874;
  wire _29876 = r95 ^ _29875;
  wire _29877 = _12298 ? coded_block[95] : r95;
  wire _29878 = _12296 ? _29876 : _29877;
  always @ (posedge reset or posedge clock) if (reset) r95 <= 1'd0; else if (_12300) r95 <= _29878;
  wire [1:0] _29879 = {_0, _2013} + {_0, _3231};
  wire [1:0] _29880 = {_0, _4384} + {_0, _7100};
  wire [2:0] _29881 = {_0, _29879} + {_0, _29880};
  wire [1:0] _29882 = {_0, _8736} + {_0, _10493};
  wire [3:0] _29883 = {_0, _29881} + {_0, _0, _29882};
  wire _29884 = _12301 < _29883;
  wire _29885 = r94 ^ _29884;
  wire _29886 = _12298 ? coded_block[94] : r94;
  wire _29887 = _12296 ? _29885 : _29886;
  always @ (posedge reset or posedge clock) if (reset) r94 <= 1'd0; else if (_12300) r94 <= _29887;
  wire [1:0] _29888 = {_0, _2044} + {_0, _3325};
  wire [1:0] _29889 = {_0, _5310} + {_0, _6462};
  wire [2:0] _29890 = {_0, _29888} + {_0, _29889};
  wire [1:0] _29891 = {_0, _9181} + {_0, _10814};
  wire [3:0] _29892 = {_0, _29890} + {_0, _0, _29891};
  wire _29893 = _12301 < _29892;
  wire _29894 = r93 ^ _29893;
  wire _29895 = _12298 ? coded_block[93] : r93;
  wire _29896 = _12296 ? _29894 : _29895;
  always @ (posedge reset or posedge clock) if (reset) r93 <= 1'd0; else if (_12300) r93 <= _29896;
  wire [1:0] _29897 = {_0, _97} + {_0, _3037};
  wire [1:0] _29898 = {_0, _4861} + {_0, _7485};
  wire [2:0] _29899 = {_0, _29897} + {_0, _29898};
  wire [1:0] _29900 = {_0, _9469} + {_0, _10621};
  wire [3:0] _29901 = {_0, _29899} + {_0, _0, _29900};
  wire _29902 = _12301 < _29901;
  wire _29903 = r92 ^ _29902;
  wire _29904 = _12298 ? coded_block[92] : r92;
  wire _29905 = _12296 ? _29903 : _29904;
  always @ (posedge reset or posedge clock) if (reset) r92 <= 1'd0; else if (_12300) r92 <= _29905;
  wire [1:0] _29906 = {_0, _128} + {_0, _3933};
  wire [1:0] _29907 = {_0, _5116} + {_0, _6942};
  wire [2:0] _29908 = {_0, _29906} + {_0, _29907};
  wire [1:0] _29909 = {_0, _9566} + {_0, _11550};
  wire [3:0] _29910 = {_0, _29908} + {_0, _0, _29909};
  wire _29911 = _12301 < _29910;
  wire _29912 = r91 ^ _29911;
  wire _29913 = _12298 ? coded_block[91] : r91;
  wire _29914 = _12296 ? _29912 : _29913;
  always @ (posedge reset or posedge clock) if (reset) r91 <= 1'd0; else if (_12300) r91 <= _29914;
  wire [1:0] _29915 = {_0, _161} + {_0, _3580};
  wire [1:0] _29916 = {_0, _6012} + {_0, _7199};
  wire [2:0] _29917 = {_0, _29915} + {_0, _29916};
  wire [1:0] _29918 = {_0, _9022} + {_0, _11644};
  wire [3:0] _29919 = {_0, _29917} + {_0, _0, _29918};
  wire _29920 = _12301 < _29919;
  wire _29921 = r90 ^ _29920;
  wire _29922 = _12298 ? coded_block[90] : r90;
  wire _29923 = _12296 ? _29921 : _29922;
  always @ (posedge reset or posedge clock) if (reset) r90 <= 1'd0; else if (_12300) r90 <= _29923;
  wire [1:0] _29924 = {_0, _192} + {_0, _3805};
  wire [1:0] _29925 = {_0, _5663} + {_0, _8092};
  wire [2:0] _29926 = {_0, _29924} + {_0, _29925};
  wire [1:0] _29927 = {_0, _9279} + {_0, _11101};
  wire [3:0] _29928 = {_0, _29926} + {_0, _0, _29927};
  wire _29929 = _12301 < _29928;
  wire _29930 = r89 ^ _29929;
  wire _29931 = _12298 ? coded_block[89] : r89;
  wire _29932 = _12296 ? _29930 : _29931;
  always @ (posedge reset or posedge clock) if (reset) r89 <= 1'd0; else if (_12300) r89 <= _29932;
  wire [1:0] _29933 = {_0, _224} + {_0, _3678};
  wire [1:0] _29934 = {_0, _5884} + {_0, _7741};
  wire [2:0] _29935 = {_0, _29933} + {_0, _29934};
  wire [1:0] _29936 = {_0, _10172} + {_0, _11358};
  wire [3:0] _29937 = {_0, _29935} + {_0, _0, _29936};
  wire _29938 = _12301 < _29937;
  wire _29939 = r88 ^ _29938;
  wire _29940 = _12298 ? coded_block[88] : r88;
  wire _29941 = _12296 ? _29939 : _29940;
  always @ (posedge reset or posedge clock) if (reset) r88 <= 1'd0; else if (_12300) r88 <= _29941;
  wire [1:0] _29942 = {_0, _255} + {_0, _4028};
  wire [1:0] _29943 = {_0, _5757} + {_0, _7965};
  wire [2:0] _29944 = {_0, _29942} + {_0, _29943};
  wire [1:0] _29945 = {_0, _9822} + {_0, _12251};
  wire [3:0] _29946 = {_0, _29944} + {_0, _0, _29945};
  wire _29947 = _12301 < _29946;
  wire _29948 = r87 ^ _29947;
  wire _29949 = _12298 ? coded_block[87] : r87;
  wire _29950 = _12296 ? _29948 : _29949;
  always @ (posedge reset or posedge clock) if (reset) r87 <= 1'd0; else if (_12300) r87 <= _29950;
  wire [1:0] _29951 = {_0, _320} + {_0, _3359};
  wire [1:0] _29952 = {_0, _4830} + {_0, _8186};
  wire [2:0] _29953 = {_0, _29951} + {_0, _29952};
  wire [1:0] _29954 = {_0, _9917} + {_0, _12124};
  wire [3:0] _29955 = {_0, _29953} + {_0, _0, _29954};
  wire _29956 = _12301 < _29955;
  wire _29957 = r86 ^ _29956;
  wire _29958 = _12298 ? coded_block[86] : r86;
  wire _29959 = _12296 ? _29957 : _29958;
  always @ (posedge reset or posedge clock) if (reset) r86 <= 1'd0; else if (_12300) r86 <= _29959;
  wire [1:0] _29960 = {_0, _352} + {_0, _2910};
  wire [1:0] _29961 = {_0, _5438} + {_0, _6908};
  wire [2:0] _29962 = {_0, _29960} + {_0, _29961};
  wire [1:0] _29963 = {_0, _8256} + {_0, _11996};
  wire [3:0] _29964 = {_0, _29962} + {_0, _0, _29963};
  wire _29965 = _12301 < _29964;
  wire _29966 = r85 ^ _29965;
  wire _29967 = _12298 ? coded_block[85] : r85;
  wire _29968 = _12296 ? _29966 : _29967;
  always @ (posedge reset or posedge clock) if (reset) r85 <= 1'd0; else if (_12300) r85 <= _29968;
  wire [1:0] _29969 = {_0, _383} + {_0, _2526};
  wire [1:0] _29970 = {_0, _4989} + {_0, _7517};
  wire [2:0] _29971 = {_0, _29969} + {_0, _29970};
  wire [1:0] _29972 = {_0, _8991} + {_0, _10335};
  wire [3:0] _29973 = {_0, _29971} + {_0, _0, _29972};
  wire _29974 = _12301 < _29973;
  wire _29975 = r84 ^ _29974;
  wire _29976 = _12298 ? coded_block[84] : r84;
  wire _29977 = _12296 ? _29975 : _29976;
  always @ (posedge reset or posedge clock) if (reset) r84 <= 1'd0; else if (_12300) r84 <= _29977;
  wire [1:0] _29978 = {_0, _416} + {_0, _3549};
  wire [1:0] _29979 = {_0, _4605} + {_0, _7069};
  wire [2:0] _29980 = {_0, _29978} + {_0, _29979};
  wire [1:0] _29981 = {_0, _9597} + {_0, _11069};
  wire [3:0] _29982 = {_0, _29980} + {_0, _0, _29981};
  wire _29983 = _12301 < _29982;
  wire _29984 = r83 ^ _29983;
  wire _29985 = _12298 ? coded_block[83] : r83;
  wire _29986 = _12296 ? _29984 : _29985;
  always @ (posedge reset or posedge clock) if (reset) r83 <= 1'd0; else if (_12300) r83 <= _29986;
  wire [1:0] _29987 = {_0, _447} + {_0, _3964};
  wire [1:0] _29988 = {_0, _5628} + {_0, _6687};
  wire [2:0] _29989 = {_0, _29987} + {_0, _29988};
  wire [1:0] _29990 = {_0, _9149} + {_0, _11677};
  wire [3:0] _29991 = {_0, _29989} + {_0, _0, _29990};
  wire _29992 = _12301 < _29991;
  wire _29993 = r82 ^ _29992;
  wire _29994 = _12298 ? coded_block[82] : r82;
  wire _29995 = _12296 ? _29993 : _29994;
  always @ (posedge reset or posedge clock) if (reset) r82 <= 1'd0; else if (_12300) r82 <= _29995;
  wire [1:0] _29996 = {_0, _479} + {_0, _2430};
  wire [1:0] _29997 = {_0, _6045} + {_0, _7710};
  wire [2:0] _29998 = {_0, _29996} + {_0, _29997};
  wire [1:0] _29999 = {_0, _8767} + {_0, _11228};
  wire [3:0] _30000 = {_0, _29998} + {_0, _0, _29999};
  wire _30001 = _12301 < _30000;
  wire _30002 = r81 ^ _30001;
  wire _30003 = _12298 ? coded_block[81] : r81;
  wire _30004 = _12296 ? _30002 : _30003;
  always @ (posedge reset or posedge clock) if (reset) r81 <= 1'd0; else if (_12300) r81 <= _30004;
  wire [1:0] _30005 = {_0, _510} + {_0, _3870};
  wire [1:0] _30006 = {_0, _4511} + {_0, _8123};
  wire [2:0] _30007 = {_0, _30005} + {_0, _30006};
  wire [1:0] _30008 = {_0, _9790} + {_0, _10846};
  wire [3:0] _30009 = {_0, _30007} + {_0, _0, _30008};
  wire _30010 = _12301 < _30009;
  wire _30011 = r80 ^ _30010;
  wire _30012 = _12298 ? coded_block[80] : r80;
  wire _30013 = _12296 ? _30011 : _30012;
  always @ (posedge reset or posedge clock) if (reset) r80 <= 1'd0; else if (_12300) r80 <= _30013;
  wire [1:0] _30014 = {_0, _576} + {_0, _2847};
  wire [1:0] _30015 = {_0, _5246} + {_0, _8028};
  wire [2:0] _30016 = {_0, _30014} + {_0, _30015};
  wire [1:0] _30017 = {_0, _8670} + {_0, _12282};
  wire [3:0] _30018 = {_0, _30016} + {_0, _0, _30017};
  wire _30019 = _12301 < _30018;
  wire _30020 = r79 ^ _30019;
  wire _30021 = _12298 ? coded_block[79] : r79;
  wire _30022 = _12296 ? _30020 : _30021;
  always @ (posedge reset or posedge clock) if (reset) r79 <= 1'd0; else if (_12300) r79 <= _30022;
  wire [1:0] _30023 = {_0, _608} + {_0, _3005};
  wire [1:0] _30024 = {_0, _4926} + {_0, _7326};
  wire [2:0] _30025 = {_0, _30023} + {_0, _30024};
  wire [1:0] _30026 = {_0, _10108} + {_0, _10748};
  wire [3:0] _30027 = {_0, _30025} + {_0, _0, _30026};
  wire _30028 = _12301 < _30027;
  wire _30029 = r78 ^ _30028;
  wire _30030 = _12298 ? coded_block[78] : r78;
  wire _30031 = _12296 ? _30029 : _30030;
  always @ (posedge reset or posedge clock) if (reset) r78 <= 1'd0; else if (_12300) r78 <= _30031;
  wire [1:0] _30032 = {_0, _639} + {_0, _2813};
  wire [1:0] _30033 = {_0, _5085} + {_0, _7005};
  wire [2:0] _30034 = {_0, _30032} + {_0, _30033};
  wire [1:0] _30035 = {_0, _9406} + {_0, _12188};
  wire [3:0] _30036 = {_0, _30034} + {_0, _0, _30035};
  wire _30037 = _12301 < _30036;
  wire _30038 = r77 ^ _30037;
  wire _30039 = _12298 ? coded_block[77] : r77;
  wire _30040 = _12296 ? _30038 : _30039;
  always @ (posedge reset or posedge clock) if (reset) r77 <= 1'd0; else if (_12300) r77 <= _30040;
  wire [1:0] _30041 = {_0, _672} + {_0, _3198};
  wire [1:0] _30042 = {_0, _4895} + {_0, _7163};
  wire [2:0] _30043 = {_0, _30041} + {_0, _30042};
  wire [1:0] _30044 = {_0, _9085} + {_0, _11485};
  wire [3:0] _30045 = {_0, _30043} + {_0, _0, _30044};
  wire _30046 = _12301 < _30045;
  wire _30047 = r76 ^ _30046;
  wire _30048 = _12298 ? coded_block[76] : r76;
  wire _30049 = _12296 ? _30047 : _30048;
  always @ (posedge reset or posedge clock) if (reset) r76 <= 1'd0; else if (_12300) r76 <= _30049;
  wire [1:0] _30050 = {_0, _703} + {_0, _2336};
  wire [1:0] _30051 = {_0, _5279} + {_0, _6973};
  wire [2:0] _30052 = {_0, _30050} + {_0, _30051};
  wire [1:0] _30053 = {_0, _9248} + {_0, _11165};
  wire [3:0] _30054 = {_0, _30052} + {_0, _0, _30053};
  wire _30055 = _12301 < _30054;
  wire _30056 = r75 ^ _30055;
  wire _30057 = _12298 ? coded_block[75] : r75;
  wire _30058 = _12296 ? _30056 : _30057;
  always @ (posedge reset or posedge clock) if (reset) r75 <= 1'd0; else if (_12300) r75 <= _30058;
  wire [1:0] _30059 = {_0, _735} + {_0, _2112};
  wire [1:0] _30060 = {_0, _4415} + {_0, _7357};
  wire [2:0] _30061 = {_0, _30059} + {_0, _30060};
  wire [1:0] _30062 = {_0, _9054} + {_0, _11326};
  wire [3:0] _30063 = {_0, _30061} + {_0, _0, _30062};
  wire _30064 = _12301 < _30063;
  wire _30065 = r74 ^ _30064;
  wire _30066 = _12298 ? coded_block[74] : r74;
  wire _30067 = _12296 ? _30065 : _30066;
  always @ (posedge reset or posedge clock) if (reset) r74 <= 1'd0; else if (_12300) r74 <= _30067;
  wire [1:0] _30068 = {_0, _766} + {_0, _2686};
  wire [1:0] _30069 = {_0, _4192} + {_0, _6494};
  wire [2:0] _30070 = {_0, _30068} + {_0, _30069};
  wire [1:0] _30071 = {_0, _9438} + {_0, _11132};
  wire [3:0] _30072 = {_0, _30070} + {_0, _0, _30071};
  wire _30073 = _12301 < _30072;
  wire _30074 = r73 ^ _30073;
  wire _30075 = _12298 ? coded_block[73] : r73;
  wire _30076 = _12296 ? _30074 : _30075;
  always @ (posedge reset or posedge clock) if (reset) r73 <= 1'd0; else if (_12300) r73 <= _30076;
  wire [1:0] _30077 = {_0, _800} + {_0, _2623};
  wire [1:0] _30078 = {_0, _4767} + {_0, _6270};
  wire [2:0] _30079 = {_0, _30077} + {_0, _30078};
  wire [1:0] _30080 = {_0, _8574} + {_0, _11516};
  wire [3:0] _30081 = {_0, _30079} + {_0, _0, _30080};
  wire _30082 = _12301 < _30081;
  wire _30083 = r72 ^ _30082;
  wire _30084 = _12298 ? coded_block[72] : r72;
  wire _30085 = _12296 ? _30083 : _30084;
  always @ (posedge reset or posedge clock) if (reset) r72 <= 1'd0; else if (_12300) r72 <= _30085;
  wire [1:0] _30086 = {_0, _831} + {_0, _3742};
  wire [1:0] _30087 = {_0, _4703} + {_0, _6845};
  wire [2:0] _30088 = {_0, _30086} + {_0, _30087};
  wire [1:0] _30089 = {_0, _8352} + {_0, _10654};
  wire [3:0] _30090 = {_0, _30088} + {_0, _0, _30089};
  wire _30091 = _12301 < _30090;
  wire _30092 = r71 ^ _30091;
  wire _30093 = _12298 ? coded_block[71] : r71;
  wire _30094 = _12296 ? _30092 : _30093;
  always @ (posedge reset or posedge clock) if (reset) r71 <= 1'd0; else if (_12300) r71 <= _30094;
  wire [1:0] _30095 = {_0, _863} + {_0, _2399};
  wire [1:0] _30096 = {_0, _5821} + {_0, _6781};
  wire [2:0] _30097 = {_0, _30095} + {_0, _30096};
  wire [1:0] _30098 = {_0, _8926} + {_0, _10430};
  wire [3:0] _30099 = {_0, _30097} + {_0, _0, _30098};
  wire _30100 = _12301 < _30099;
  wire _30101 = r70 ^ _30100;
  wire _30102 = _12298 ? coded_block[70] : r70;
  wire _30103 = _12296 ? _30101 : _30102;
  always @ (posedge reset or posedge clock) if (reset) r70 <= 1'd0; else if (_12300) r70 <= _30103;
  wire [1:0] _30104 = {_0, _894} + {_0, _3997};
  wire [1:0] _30105 = {_0, _4478} + {_0, _7900};
  wire [2:0] _30106 = {_0, _30104} + {_0, _30105};
  wire [1:0] _30107 = {_0, _8863} + {_0, _11004};
  wire [3:0] _30108 = {_0, _30106} + {_0, _0, _30107};
  wire _30109 = _12301 < _30108;
  wire _30110 = r69 ^ _30109;
  wire _30111 = _12298 ? coded_block[69] : r69;
  wire _30112 = _12296 ? _30110 : _30111;
  always @ (posedge reset or posedge clock) if (reset) r69 <= 1'd0; else if (_12300) r69 <= _30112;
  wire [1:0] _30113 = {_0, _927} + {_0, _3709};
  wire [1:0] _30114 = {_0, _6076} + {_0, _6558};
  wire [2:0] _30115 = {_0, _30113} + {_0, _30114};
  wire [1:0] _30116 = {_0, _9980} + {_0, _10941};
  wire [3:0] _30117 = {_0, _30115} + {_0, _0, _30116};
  wire _30118 = _12301 < _30117;
  wire _30119 = r68 ^ _30118;
  wire _30120 = _12298 ? coded_block[68] : r68;
  wire _30121 = _12296 ? _30119 : _30120;
  always @ (posedge reset or posedge clock) if (reset) r68 <= 1'd0; else if (_12300) r68 <= _30121;
  wire [1:0] _30122 = {_0, _958} + {_0, _2655};
  wire [1:0] _30123 = {_0, _5790} + {_0, _8155};
  wire [2:0] _30124 = {_0, _30122} + {_0, _30123};
  wire [1:0] _30125 = {_0, _8638} + {_0, _12061};
  wire [3:0] _30126 = {_0, _30124} + {_0, _0, _30125};
  wire _30127 = _12301 < _30126;
  wire _30128 = r67 ^ _30127;
  wire _30129 = _12298 ? coded_block[67] : r67;
  wire _30130 = _12296 ? _30128 : _30129;
  always @ (posedge reset or posedge clock) if (reset) r67 <= 1'd0; else if (_12300) r67 <= _30130;
  wire [1:0] _30131 = {_0, _990} + {_0, _2144};
  wire [1:0] _30132 = {_0, _4734} + {_0, _7868};
  wire [2:0] _30133 = {_0, _30131} + {_0, _30132};
  wire [1:0] _30134 = {_0, _10235} + {_0, _10717};
  wire [3:0] _30135 = {_0, _30133} + {_0, _0, _30134};
  wire _30136 = _12301 < _30135;
  wire _30137 = r66 ^ _30136;
  wire _30138 = _12298 ? coded_block[66] : r66;
  wire _30139 = _12296 ? _30137 : _30138;
  always @ (posedge reset or posedge clock) if (reset) r66 <= 1'd0; else if (_12300) r66 <= _30139;
  wire [1:0] _30140 = {_0, _1021} + {_0, _3135};
  wire [1:0] _30141 = {_0, _4223} + {_0, _6814};
  wire [2:0] _30142 = {_0, _30140} + {_0, _30141};
  wire [1:0] _30143 = {_0, _9949} + {_0, _10303};
  wire [3:0] _30144 = {_0, _30142} + {_0, _0, _30143};
  wire _30145 = _12301 < _30144;
  wire _30146 = r65 ^ _30145;
  wire _30147 = _12298 ? coded_block[65] : r65;
  wire _30148 = _12296 ? _30146 : _30147;
  always @ (posedge reset or posedge clock) if (reset) r65 <= 1'd0; else if (_12300) r65 <= _30148;
  wire [1:0] _30149 = {_0, _1057} + {_0, _3901};
  wire [1:0] _30150 = {_0, _5215} + {_0, _6303};
  wire [2:0] _30151 = {_0, _30149} + {_0, _30150};
  wire [1:0] _30152 = {_0, _8894} + {_0, _12027};
  wire [3:0] _30153 = {_0, _30151} + {_0, _0, _30152};
  wire _30154 = _12301 < _30153;
  wire _30155 = r64 ^ _30154;
  wire _30156 = _12298 ? coded_block[64] : r64;
  wire _30157 = _12296 ? _30155 : _30156;
  always @ (posedge reset or posedge clock) if (reset) r64 <= 1'd0; else if (_12300) r64 <= _30157;
  wire [1:0] _30158 = {_0, _1088} + {_0, _3068};
  wire [1:0] _30159 = {_0, _5981} + {_0, _7293};
  wire [2:0] _30160 = {_0, _30158} + {_0, _30159};
  wire [1:0] _30161 = {_0, _8383} + {_0, _10973};
  wire [3:0] _30162 = {_0, _30160} + {_0, _0, _30161};
  wire _30163 = _12301 < _30162;
  wire _30164 = r63 ^ _30163;
  wire _30165 = _12298 ? coded_block[63] : r63;
  wire _30166 = _12296 ? _30164 : _30165;
  always @ (posedge reset or posedge clock) if (reset) r63 <= 1'd0; else if (_12300) r63 <= _30166;
  wire [1:0] _30167 = {_0, _1120} + {_0, _2592};
  wire [1:0] _30168 = {_0, _5152} + {_0, _8059};
  wire [2:0] _30169 = {_0, _30167} + {_0, _30168};
  wire [1:0] _30170 = {_0, _9375} + {_0, _10462};
  wire [3:0] _30171 = {_0, _30169} + {_0, _0, _30170};
  wire _30172 = _12301 < _30171;
  wire _30173 = r62 ^ _30172;
  wire _30174 = _12298 ? coded_block[62] : r62;
  wire _30175 = _12296 ? _30173 : _30174;
  always @ (posedge reset or posedge clock) if (reset) r62 <= 1'd0; else if (_12300) r62 <= _30175;
  wire [1:0] _30176 = {_0, _1151} + {_0, _2719};
  wire [1:0] _30177 = {_0, _4671} + {_0, _7230};
  wire [2:0] _30178 = {_0, _30176} + {_0, _30177};
  wire [1:0] _30179 = {_0, _10141} + {_0, _11453};
  wire [3:0] _30180 = {_0, _30178} + {_0, _0, _30179};
  wire _30181 = _12301 < _30180;
  wire _30182 = r61 ^ _30181;
  wire _30183 = _12298 ? coded_block[61] : r61;
  wire _30184 = _12296 ? _30182 : _30183;
  always @ (posedge reset or posedge clock) if (reset) r61 <= 1'd0; else if (_12300) r61 <= _30184;
  wire [1:0] _30185 = {_0, _1184} + {_0, _4060};
  wire [1:0] _30186 = {_0, _4798} + {_0, _6750};
  wire [2:0] _30187 = {_0, _30185} + {_0, _30186};
  wire [1:0] _30188 = {_0, _9311} + {_0, _12219};
  wire [3:0] _30189 = {_0, _30187} + {_0, _0, _30188};
  wire _30190 = _12301 < _30189;
  wire _30191 = r60 ^ _30190;
  wire _30192 = _12298 ? coded_block[60] : r60;
  wire _30193 = _12296 ? _30191 : _30192;
  always @ (posedge reset or posedge clock) if (reset) r60 <= 1'd0; else if (_12300) r60 <= _30193;
  wire [1:0] _30194 = {_0, _1215} + {_0, _3294};
  wire [1:0] _30195 = {_0, _6139} + {_0, _6877};
  wire [2:0] _30196 = {_0, _30194} + {_0, _30195};
  wire [1:0] _30197 = {_0, _8830} + {_0, _11389};
  wire [3:0] _30198 = {_0, _30196} + {_0, _0, _30197};
  wire _30199 = _12301 < _30198;
  wire _30200 = r59 ^ _30199;
  wire _30201 = _12298 ? coded_block[59] : r59;
  wire _30202 = _12296 ? _30200 : _30201;
  always @ (posedge reset or posedge clock) if (reset) r59 <= 1'd0; else if (_12300) r59 <= _30202;
  wire [1:0] _30203 = {_0, _1247} + {_0, _3262};
  wire [1:0] _30204 = {_0, _5373} + {_0, _6207};
  wire [2:0] _30205 = {_0, _30203} + {_0, _30204};
  wire [1:0] _30206 = {_0, _8957} + {_0, _10910};
  wire [3:0] _30207 = {_0, _30205} + {_0, _0, _30206};
  wire _30208 = _12301 < _30207;
  wire _30209 = r58 ^ _30208;
  wire _30210 = _12298 ? coded_block[58] : r58;
  wire _30211 = _12296 ? _30209 : _30210;
  always @ (posedge reset or posedge clock) if (reset) r58 <= 1'd0; else if (_12300) r58 <= _30211;
  wire [1:0] _30212 = {_0, _1278} + {_0, _4091};
  wire [1:0] _30213 = {_0, _5342} + {_0, _7454};
  wire [2:0] _30214 = {_0, _30212} + {_0, _30213};
  wire [1:0] _30215 = {_0, _8288} + {_0, _11038};
  wire [3:0] _30216 = {_0, _30214} + {_0, _0, _30215};
  wire _30217 = _12301 < _30216;
  wire _30218 = r57 ^ _30217;
  wire _30219 = _12298 ? coded_block[57] : r57;
  wire _30220 = _12296 ? _30218 : _30219;
  always @ (posedge reset or posedge clock) if (reset) r57 <= 1'd0; else if (_12300) r57 <= _30220;
  wire [1:0] _30221 = {_0, _1312} + {_0, _2367};
  wire [1:0] _30222 = {_0, _4160} + {_0, _7420};
  wire [2:0] _30223 = {_0, _30221} + {_0, _30222};
  wire [1:0] _30224 = {_0, _9534} + {_0, _10366};
  wire [3:0] _30225 = {_0, _30223} + {_0, _0, _30224};
  wire _30226 = _12301 < _30225;
  wire _30227 = r56 ^ _30226;
  wire _30228 = _12298 ? coded_block[56] : r56;
  wire _30229 = _12296 ? _30227 : _30228;
  always @ (posedge reset or posedge clock) if (reset) r56 <= 1'd0; else if (_12300) r56 <= _30229;
  wire [1:0] _30230 = {_0, _1343} + {_0, _3773};
  wire [1:0] _30231 = {_0, _4447} + {_0, _6239};
  wire [2:0] _30232 = {_0, _30230} + {_0, _30231};
  wire [1:0] _30233 = {_0, _9503} + {_0, _11613};
  wire [3:0] _30234 = {_0, _30232} + {_0, _0, _30233};
  wire _30235 = _12301 < _30234;
  wire _30236 = r55 ^ _30235;
  wire _30237 = _12298 ? coded_block[55] : r55;
  wire _30238 = _12296 ? _30236 : _30237;
  always @ (posedge reset or posedge clock) if (reset) r55 <= 1'd0; else if (_12300) r55 <= _30238;
  wire [1:0] _30239 = {_0, _1375} + {_0, _3615};
  wire [1:0] _30240 = {_0, _5853} + {_0, _6525};
  wire [2:0] _30241 = {_0, _30239} + {_0, _30240};
  wire [1:0] _30242 = {_0, _8319} + {_0, _11581};
  wire [3:0] _30243 = {_0, _30241} + {_0, _0, _30242};
  wire _30244 = _12301 < _30243;
  wire _30245 = r54 ^ _30244;
  wire _30246 = _12298 ? coded_block[54] : r54;
  wire _30247 = _12296 ? _30245 : _30246;
  always @ (posedge reset or posedge clock) if (reset) r54 <= 1'd0; else if (_12300) r54 <= _30247;
  wire [1:0] _30248 = {_0, _34} + {_0, _2081};
  wire [1:0] _30249 = {_0, _4129} + {_0, _6176};
  wire [2:0] _30250 = {_0, _30248} + {_0, _30249};
  wire [1:0] _30251 = {_0, _8225} + {_0, _10272};
  wire [3:0] _30252 = {_0, _30250} + {_0, _0, _30251};
  wire _30253 = _12301 < _30252;
  wire _30254 = r53 ^ _30253;
  wire _30255 = _12298 ? coded_block[53] : r53;
  wire _30256 = _12296 ? _30254 : _30255;
  always @ (posedge reset or posedge clock) if (reset) r53 <= 1'd0; else if (_12300) r53 <= _30256;
  wire [1:0] _30257 = {_0, _2044} + {_0, _4091};
  wire [1:0] _30258 = {_0, _6139} + {_0, _8186};
  wire [2:0] _30259 = {_0, _30257} + {_0, _30258};
  wire [1:0] _30260 = {_0, _10235} + {_0, _12282};
  wire [3:0] _30261 = {_0, _30259} + {_0, _0, _30260};
  wire _30262 = _12301 < _30261;
  wire _30263 = r52 ^ _30262;
  wire _30264 = _12298 ? coded_block[52] : r52;
  wire _30265 = _12296 ? _30263 : _30264;
  always @ (posedge reset or posedge clock) if (reset) r52 <= 1'd0; else if (_12300) r52 <= _30265;
  wire [1:0] _30266 = {_0, _65} + {_0, _2112};
  wire [1:0] _30267 = {_0, _4160} + {_0, _6207};
  wire [2:0] _30268 = {_0, _30266} + {_0, _30267};
  wire [1:0] _30269 = {_0, _8256} + {_0, _10303};
  wire [3:0] _30270 = {_0, _30268} + {_0, _0, _30269};
  wire _30271 = _12301 < _30270;
  wire _30272 = r51 ^ _30271;
  wire _30273 = _12298 ? coded_block[51] : r51;
  wire _30274 = _12296 ? _30272 : _30273;
  always @ (posedge reset or posedge clock) if (reset) r51 <= 1'd0; else if (_12300) r51 <= _30274;
  wire [1:0] _30275 = {_0, _97} + {_0, _2144};
  wire [1:0] _30276 = {_0, _4192} + {_0, _6239};
  wire [2:0] _30277 = {_0, _30275} + {_0, _30276};
  wire [1:0] _30278 = {_0, _8288} + {_0, _10335};
  wire [3:0] _30279 = {_0, _30277} + {_0, _0, _30278};
  wire _30280 = _12301 < _30279;
  wire _30281 = r50 ^ _30280;
  wire _30282 = _12298 ? coded_block[50] : r50;
  wire _30283 = _12296 ? _30281 : _30282;
  always @ (posedge reset or posedge clock) if (reset) r50 <= 1'd0; else if (_12300) r50 <= _30283;
  wire [1:0] _30284 = {_0, _161} + {_0, _2208};
  wire [1:0] _30285 = {_0, _4256} + {_0, _6303};
  wire [2:0] _30286 = {_0, _30284} + {_0, _30285};
  wire [1:0] _30287 = {_0, _8352} + {_0, _10399};
  wire [3:0] _30288 = {_0, _30286} + {_0, _0, _30287};
  wire _30289 = _12301 < _30288;
  wire _30290 = r49 ^ _30289;
  wire _30291 = _12298 ? coded_block[49] : r49;
  wire _30292 = _12296 ? _30290 : _30291;
  always @ (posedge reset or posedge clock) if (reset) r49 <= 1'd0; else if (_12300) r49 <= _30292;
  wire [1:0] _30293 = {_0, _192} + {_0, _2239};
  wire [1:0] _30294 = {_0, _4287} + {_0, _6334};
  wire [2:0] _30295 = {_0, _30293} + {_0, _30294};
  wire [1:0] _30296 = {_0, _8383} + {_0, _10430};
  wire [3:0] _30297 = {_0, _30295} + {_0, _0, _30296};
  wire _30298 = _12301 < _30297;
  wire _30299 = r48 ^ _30298;
  wire _30300 = _12298 ? coded_block[48] : r48;
  wire _30301 = _12296 ? _30299 : _30300;
  always @ (posedge reset or posedge clock) if (reset) r48 <= 1'd0; else if (_12300) r48 <= _30301;
  wire [1:0] _30302 = {_0, _224} + {_0, _2271};
  wire [1:0] _30303 = {_0, _4319} + {_0, _6366};
  wire [2:0] _30304 = {_0, _30302} + {_0, _30303};
  wire [1:0] _30305 = {_0, _8415} + {_0, _10462};
  wire [3:0] _30306 = {_0, _30304} + {_0, _0, _30305};
  wire _30307 = _12301 < _30306;
  wire _30308 = r47 ^ _30307;
  wire _30309 = _12298 ? coded_block[47] : r47;
  wire _30310 = _12296 ? _30308 : _30309;
  always @ (posedge reset or posedge clock) if (reset) r47 <= 1'd0; else if (_12300) r47 <= _30310;
  wire [1:0] _30311 = {_0, _255} + {_0, _2302};
  wire [1:0] _30312 = {_0, _4350} + {_0, _6397};
  wire [2:0] _30313 = {_0, _30311} + {_0, _30312};
  wire [1:0] _30314 = {_0, _8446} + {_0, _10493};
  wire [3:0] _30315 = {_0, _30313} + {_0, _0, _30314};
  wire _30316 = _12301 < _30315;
  wire _30317 = r46 ^ _30316;
  wire _30318 = _12298 ? coded_block[46] : r46;
  wire _30319 = _12296 ? _30317 : _30318;
  always @ (posedge reset or posedge clock) if (reset) r46 <= 1'd0; else if (_12300) r46 <= _30319;
  wire [1:0] _30320 = {_0, _289} + {_0, _2336};
  wire [1:0] _30321 = {_0, _4384} + {_0, _6431};
  wire [2:0] _30322 = {_0, _30320} + {_0, _30321};
  wire [1:0] _30323 = {_0, _8480} + {_0, _10527};
  wire [3:0] _30324 = {_0, _30322} + {_0, _0, _30323};
  wire _30325 = _12301 < _30324;
  wire _30326 = r45 ^ _30325;
  wire _30327 = _12298 ? coded_block[45] : r45;
  wire _30328 = _12296 ? _30326 : _30327;
  always @ (posedge reset or posedge clock) if (reset) r45 <= 1'd0; else if (_12300) r45 <= _30328;
  wire [1:0] _30329 = {_0, _320} + {_0, _2367};
  wire [1:0] _30330 = {_0, _4415} + {_0, _6462};
  wire [2:0] _30331 = {_0, _30329} + {_0, _30330};
  wire [1:0] _30332 = {_0, _8511} + {_0, _10558};
  wire [3:0] _30333 = {_0, _30331} + {_0, _0, _30332};
  wire _30334 = _12301 < _30333;
  wire _30335 = r44 ^ _30334;
  wire _30336 = _12298 ? coded_block[44] : r44;
  wire _30337 = _12296 ? _30335 : _30336;
  always @ (posedge reset or posedge clock) if (reset) r44 <= 1'd0; else if (_12300) r44 <= _30337;
  wire [1:0] _30338 = {_0, _352} + {_0, _2399};
  wire [1:0] _30339 = {_0, _4447} + {_0, _6494};
  wire [2:0] _30340 = {_0, _30338} + {_0, _30339};
  wire [1:0] _30341 = {_0, _8543} + {_0, _10590};
  wire [3:0] _30342 = {_0, _30340} + {_0, _0, _30341};
  wire _30343 = _12301 < _30342;
  wire _30344 = r43 ^ _30343;
  wire _30345 = _12298 ? coded_block[43] : r43;
  wire _30346 = _12296 ? _30344 : _30345;
  always @ (posedge reset or posedge clock) if (reset) r43 <= 1'd0; else if (_12300) r43 <= _30346;
  wire [1:0] _30347 = {_0, _383} + {_0, _2430};
  wire [1:0] _30348 = {_0, _4478} + {_0, _6525};
  wire [2:0] _30349 = {_0, _30347} + {_0, _30348};
  wire [1:0] _30350 = {_0, _8574} + {_0, _10621};
  wire [3:0] _30351 = {_0, _30349} + {_0, _0, _30350};
  wire _30352 = _12301 < _30351;
  wire _30353 = r42 ^ _30352;
  wire _30354 = _12298 ? coded_block[42] : r42;
  wire _30355 = _12296 ? _30353 : _30354;
  always @ (posedge reset or posedge clock) if (reset) r42 <= 1'd0; else if (_12300) r42 <= _30355;
  wire [1:0] _30356 = {_0, _416} + {_0, _2463};
  wire [1:0] _30357 = {_0, _4511} + {_0, _6558};
  wire [2:0] _30358 = {_0, _30356} + {_0, _30357};
  wire [1:0] _30359 = {_0, _8607} + {_0, _10654};
  wire [3:0] _30360 = {_0, _30358} + {_0, _0, _30359};
  wire _30361 = _12301 < _30360;
  wire _30362 = r41 ^ _30361;
  wire _30363 = _12298 ? coded_block[41] : r41;
  wire _30364 = _12296 ? _30362 : _30363;
  always @ (posedge reset or posedge clock) if (reset) r41 <= 1'd0; else if (_12300) r41 <= _30364;
  wire [1:0] _30365 = {_0, _479} + {_0, _2526};
  wire [1:0] _30366 = {_0, _4574} + {_0, _6621};
  wire [2:0] _30367 = {_0, _30365} + {_0, _30366};
  wire [1:0] _30368 = {_0, _8670} + {_0, _10717};
  wire [3:0] _30369 = {_0, _30367} + {_0, _0, _30368};
  wire _30370 = _12301 < _30369;
  wire _30371 = r40 ^ _30370;
  wire _30372 = _12298 ? coded_block[40] : r40;
  wire _30373 = _12296 ? _30371 : _30372;
  always @ (posedge reset or posedge clock) if (reset) r40 <= 1'd0; else if (_12300) r40 <= _30373;
  wire [1:0] _30374 = {_0, _510} + {_0, _2557};
  wire [1:0] _30375 = {_0, _4605} + {_0, _6652};
  wire [2:0] _30376 = {_0, _30374} + {_0, _30375};
  wire [1:0] _30377 = {_0, _8701} + {_0, _10748};
  wire [3:0] _30378 = {_0, _30376} + {_0, _0, _30377};
  wire _30379 = _12301 < _30378;
  wire _30380 = r39 ^ _30379;
  wire _30381 = _12298 ? coded_block[39] : r39;
  wire _30382 = _12296 ? _30380 : _30381;
  always @ (posedge reset or posedge clock) if (reset) r39 <= 1'd0; else if (_12300) r39 <= _30382;
  wire [1:0] _30383 = {_0, _545} + {_0, _2592};
  wire [1:0] _30384 = {_0, _4640} + {_0, _6687};
  wire [2:0] _30385 = {_0, _30383} + {_0, _30384};
  wire [1:0] _30386 = {_0, _8736} + {_0, _10783};
  wire [3:0] _30387 = {_0, _30385} + {_0, _0, _30386};
  wire _30388 = _12301 < _30387;
  wire _30389 = r38 ^ _30388;
  wire _30390 = _12298 ? coded_block[38] : r38;
  wire _30391 = _12296 ? _30389 : _30390;
  always @ (posedge reset or posedge clock) if (reset) r38 <= 1'd0; else if (_12300) r38 <= _30391;
  wire [1:0] _30392 = {_0, _576} + {_0, _2623};
  wire [1:0] _30393 = {_0, _4671} + {_0, _6718};
  wire [2:0] _30394 = {_0, _30392} + {_0, _30393};
  wire [1:0] _30395 = {_0, _8767} + {_0, _10814};
  wire [3:0] _30396 = {_0, _30394} + {_0, _0, _30395};
  wire _30397 = _12301 < _30396;
  wire _30398 = r37 ^ _30397;
  wire _30399 = _12298 ? coded_block[37] : r37;
  wire _30400 = _12296 ? _30398 : _30399;
  always @ (posedge reset or posedge clock) if (reset) r37 <= 1'd0; else if (_12300) r37 <= _30400;
  wire [1:0] _30401 = {_0, _608} + {_0, _2655};
  wire [1:0] _30402 = {_0, _4703} + {_0, _6750};
  wire [2:0] _30403 = {_0, _30401} + {_0, _30402};
  wire [1:0] _30404 = {_0, _8799} + {_0, _10846};
  wire [3:0] _30405 = {_0, _30403} + {_0, _0, _30404};
  wire _30406 = _12301 < _30405;
  wire _30407 = r36 ^ _30406;
  wire _30408 = _12298 ? coded_block[36] : r36;
  wire _30409 = _12296 ? _30407 : _30408;
  always @ (posedge reset or posedge clock) if (reset) r36 <= 1'd0; else if (_12300) r36 <= _30409;
  wire [1:0] _30410 = {_0, _639} + {_0, _2686};
  wire [1:0] _30411 = {_0, _4734} + {_0, _6781};
  wire [2:0] _30412 = {_0, _30410} + {_0, _30411};
  wire [1:0] _30413 = {_0, _8830} + {_0, _10877};
  wire [3:0] _30414 = {_0, _30412} + {_0, _0, _30413};
  wire _30415 = _12301 < _30414;
  wire _30416 = r35 ^ _30415;
  wire _30417 = _12298 ? coded_block[35] : r35;
  wire _30418 = _12296 ? _30416 : _30417;
  always @ (posedge reset or posedge clock) if (reset) r35 <= 1'd0; else if (_12300) r35 <= _30418;
  wire [1:0] _30419 = {_0, _672} + {_0, _2719};
  wire [1:0] _30420 = {_0, _4767} + {_0, _6814};
  wire [2:0] _30421 = {_0, _30419} + {_0, _30420};
  wire [1:0] _30422 = {_0, _8863} + {_0, _10910};
  wire [3:0] _30423 = {_0, _30421} + {_0, _0, _30422};
  wire _30424 = _12301 < _30423;
  wire _30425 = r34 ^ _30424;
  wire _30426 = _12298 ? coded_block[34] : r34;
  wire _30427 = _12296 ? _30425 : _30426;
  always @ (posedge reset or posedge clock) if (reset) r34 <= 1'd0; else if (_12300) r34 <= _30427;
  wire [1:0] _30428 = {_0, _703} + {_0, _2750};
  wire [1:0] _30429 = {_0, _4798} + {_0, _6845};
  wire [2:0] _30430 = {_0, _30428} + {_0, _30429};
  wire [1:0] _30431 = {_0, _8894} + {_0, _10941};
  wire [3:0] _30432 = {_0, _30430} + {_0, _0, _30431};
  wire _30433 = _12301 < _30432;
  wire _30434 = r33 ^ _30433;
  wire _30435 = _12298 ? coded_block[33] : r33;
  wire _30436 = _12296 ? _30434 : _30435;
  always @ (posedge reset or posedge clock) if (reset) r33 <= 1'd0; else if (_12300) r33 <= _30436;
  wire [1:0] _30437 = {_0, _735} + {_0, _2782};
  wire [1:0] _30438 = {_0, _4830} + {_0, _6877};
  wire [2:0] _30439 = {_0, _30437} + {_0, _30438};
  wire [1:0] _30440 = {_0, _8926} + {_0, _10973};
  wire [3:0] _30441 = {_0, _30439} + {_0, _0, _30440};
  wire _30442 = _12301 < _30441;
  wire _30443 = r32 ^ _30442;
  wire _30444 = _12298 ? coded_block[32] : r32;
  wire _30445 = _12296 ? _30443 : _30444;
  always @ (posedge reset or posedge clock) if (reset) r32 <= 1'd0; else if (_12300) r32 <= _30445;
  wire [1:0] _30446 = {_0, _766} + {_0, _2813};
  wire [1:0] _30447 = {_0, _4861} + {_0, _6908};
  wire [2:0] _30448 = {_0, _30446} + {_0, _30447};
  wire [1:0] _30449 = {_0, _8957} + {_0, _11004};
  wire [3:0] _30450 = {_0, _30448} + {_0, _0, _30449};
  wire _30451 = _12301 < _30450;
  wire _30452 = r31 ^ _30451;
  wire _30453 = _12298 ? coded_block[31] : r31;
  wire _30454 = _12296 ? _30452 : _30453;
  always @ (posedge reset or posedge clock) if (reset) r31 <= 1'd0; else if (_12300) r31 <= _30454;
  wire [1:0] _30455 = {_0, _800} + {_0, _2847};
  wire [1:0] _30456 = {_0, _4895} + {_0, _6942};
  wire [2:0] _30457 = {_0, _30455} + {_0, _30456};
  wire [1:0] _30458 = {_0, _8991} + {_0, _11038};
  wire [3:0] _30459 = {_0, _30457} + {_0, _0, _30458};
  wire _30460 = _12301 < _30459;
  wire _30461 = r30 ^ _30460;
  wire _30462 = _12298 ? coded_block[30] : r30;
  wire _30463 = _12296 ? _30461 : _30462;
  always @ (posedge reset or posedge clock) if (reset) r30 <= 1'd0; else if (_12300) r30 <= _30463;
  wire [1:0] _30464 = {_0, _831} + {_0, _2878};
  wire [1:0] _30465 = {_0, _4926} + {_0, _6973};
  wire [2:0] _30466 = {_0, _30464} + {_0, _30465};
  wire [1:0] _30467 = {_0, _9022} + {_0, _11069};
  wire [3:0] _30468 = {_0, _30466} + {_0, _0, _30467};
  wire _30469 = _12301 < _30468;
  wire _30470 = r29 ^ _30469;
  wire _30471 = _12298 ? coded_block[29] : r29;
  wire _30472 = _12296 ? _30470 : _30471;
  always @ (posedge reset or posedge clock) if (reset) r29 <= 1'd0; else if (_12300) r29 <= _30472;
  wire [1:0] _30473 = {_0, _863} + {_0, _2910};
  wire [1:0] _30474 = {_0, _4958} + {_0, _7005};
  wire [2:0] _30475 = {_0, _30473} + {_0, _30474};
  wire [1:0] _30476 = {_0, _9054} + {_0, _11101};
  wire [3:0] _30477 = {_0, _30475} + {_0, _0, _30476};
  wire _30478 = _12301 < _30477;
  wire _30479 = r28 ^ _30478;
  wire _30480 = _12298 ? coded_block[28] : r28;
  wire _30481 = _12296 ? _30479 : _30480;
  always @ (posedge reset or posedge clock) if (reset) r28 <= 1'd0; else if (_12300) r28 <= _30481;
  wire [1:0] _30482 = {_0, _894} + {_0, _2941};
  wire [1:0] _30483 = {_0, _4989} + {_0, _7036};
  wire [2:0] _30484 = {_0, _30482} + {_0, _30483};
  wire [1:0] _30485 = {_0, _9085} + {_0, _11132};
  wire [3:0] _30486 = {_0, _30484} + {_0, _0, _30485};
  wire _30487 = _12301 < _30486;
  wire _30488 = r27 ^ _30487;
  wire _30489 = _12298 ? coded_block[27] : r27;
  wire _30490 = _12296 ? _30488 : _30489;
  always @ (posedge reset or posedge clock) if (reset) r27 <= 1'd0; else if (_12300) r27 <= _30490;
  wire [1:0] _30491 = {_0, _927} + {_0, _2974};
  wire [1:0] _30492 = {_0, _5022} + {_0, _7069};
  wire [2:0] _30493 = {_0, _30491} + {_0, _30492};
  wire [1:0] _30494 = {_0, _9118} + {_0, _11165};
  wire [3:0] _30495 = {_0, _30493} + {_0, _0, _30494};
  wire _30496 = _12301 < _30495;
  wire _30497 = r26 ^ _30496;
  wire _30498 = _12298 ? coded_block[26] : r26;
  wire _30499 = _12296 ? _30497 : _30498;
  always @ (posedge reset or posedge clock) if (reset) r26 <= 1'd0; else if (_12300) r26 <= _30499;
  wire [1:0] _30500 = {_0, _958} + {_0, _3005};
  wire [1:0] _30501 = {_0, _5053} + {_0, _7100};
  wire [2:0] _30502 = {_0, _30500} + {_0, _30501};
  wire [1:0] _30503 = {_0, _9149} + {_0, _11196};
  wire [3:0] _30504 = {_0, _30502} + {_0, _0, _30503};
  wire _30505 = _12301 < _30504;
  wire _30506 = r25 ^ _30505;
  wire _30507 = _12298 ? coded_block[25] : r25;
  wire _30508 = _12296 ? _30506 : _30507;
  always @ (posedge reset or posedge clock) if (reset) r25 <= 1'd0; else if (_12300) r25 <= _30508;
  wire [1:0] _30509 = {_0, _990} + {_0, _3037};
  wire [1:0] _30510 = {_0, _5085} + {_0, _7132};
  wire [2:0] _30511 = {_0, _30509} + {_0, _30510};
  wire [1:0] _30512 = {_0, _9181} + {_0, _11228};
  wire [3:0] _30513 = {_0, _30511} + {_0, _0, _30512};
  wire _30514 = _12301 < _30513;
  wire _30515 = r24 ^ _30514;
  wire _30516 = _12298 ? coded_block[24] : r24;
  wire _30517 = _12296 ? _30515 : _30516;
  always @ (posedge reset or posedge clock) if (reset) r24 <= 1'd0; else if (_12300) r24 <= _30517;
  wire [1:0] _30518 = {_0, _1021} + {_0, _3068};
  wire [1:0] _30519 = {_0, _5116} + {_0, _7163};
  wire [2:0] _30520 = {_0, _30518} + {_0, _30519};
  wire [1:0] _30521 = {_0, _9212} + {_0, _11259};
  wire [3:0] _30522 = {_0, _30520} + {_0, _0, _30521};
  wire _30523 = _12301 < _30522;
  wire _30524 = r23 ^ _30523;
  wire _30525 = _12298 ? coded_block[23] : r23;
  wire _30526 = _12296 ? _30524 : _30525;
  always @ (posedge reset or posedge clock) if (reset) r23 <= 1'd0; else if (_12300) r23 <= _30526;
  wire [1:0] _30527 = {_0, _1057} + {_0, _3104};
  wire [1:0] _30528 = {_0, _5152} + {_0, _7199};
  wire [2:0] _30529 = {_0, _30527} + {_0, _30528};
  wire [1:0] _30530 = {_0, _9248} + {_0, _11295};
  wire [3:0] _30531 = {_0, _30529} + {_0, _0, _30530};
  wire _30532 = _12301 < _30531;
  wire _30533 = r22 ^ _30532;
  wire _30534 = _12298 ? coded_block[22] : r22;
  wire _30535 = _12296 ? _30533 : _30534;
  always @ (posedge reset or posedge clock) if (reset) r22 <= 1'd0; else if (_12300) r22 <= _30535;
  wire [1:0] _30536 = {_0, _1088} + {_0, _3135};
  wire [1:0] _30537 = {_0, _5183} + {_0, _7230};
  wire [2:0] _30538 = {_0, _30536} + {_0, _30537};
  wire [1:0] _30539 = {_0, _9279} + {_0, _11326};
  wire [3:0] _30540 = {_0, _30538} + {_0, _0, _30539};
  wire _30541 = _12301 < _30540;
  wire _30542 = r21 ^ _30541;
  wire _30543 = _12298 ? coded_block[21] : r21;
  wire _30544 = _12296 ? _30542 : _30543;
  always @ (posedge reset or posedge clock) if (reset) r21 <= 1'd0; else if (_12300) r21 <= _30544;
  wire [1:0] _30545 = {_0, _1120} + {_0, _3167};
  wire [1:0] _30546 = {_0, _5215} + {_0, _7262};
  wire [2:0] _30547 = {_0, _30545} + {_0, _30546};
  wire [1:0] _30548 = {_0, _9311} + {_0, _11358};
  wire [3:0] _30549 = {_0, _30547} + {_0, _0, _30548};
  wire _30550 = _12301 < _30549;
  wire _30551 = r20 ^ _30550;
  wire _30552 = _12298 ? coded_block[20] : r20;
  wire _30553 = _12296 ? _30551 : _30552;
  always @ (posedge reset or posedge clock) if (reset) r20 <= 1'd0; else if (_12300) r20 <= _30553;
  wire [1:0] _30554 = {_0, _1151} + {_0, _3198};
  wire [1:0] _30555 = {_0, _5246} + {_0, _7293};
  wire [2:0] _30556 = {_0, _30554} + {_0, _30555};
  wire [1:0] _30557 = {_0, _9342} + {_0, _11389};
  wire [3:0] _30558 = {_0, _30556} + {_0, _0, _30557};
  wire _30559 = _12301 < _30558;
  wire _30560 = r19 ^ _30559;
  wire _30561 = _12298 ? coded_block[19] : r19;
  wire _30562 = _12296 ? _30560 : _30561;
  always @ (posedge reset or posedge clock) if (reset) r19 <= 1'd0; else if (_12300) r19 <= _30562;
  wire [1:0] _30563 = {_0, _1184} + {_0, _3231};
  wire [1:0] _30564 = {_0, _5279} + {_0, _7326};
  wire [2:0] _30565 = {_0, _30563} + {_0, _30564};
  wire [1:0] _30566 = {_0, _9375} + {_0, _11422};
  wire [3:0] _30567 = {_0, _30565} + {_0, _0, _30566};
  wire _30568 = _12301 < _30567;
  wire _30569 = r18 ^ _30568;
  wire _30570 = _12298 ? coded_block[18] : r18;
  wire _30571 = _12296 ? _30569 : _30570;
  always @ (posedge reset or posedge clock) if (reset) r18 <= 1'd0; else if (_12300) r18 <= _30571;
  wire [1:0] _30572 = {_0, _1215} + {_0, _3262};
  wire [1:0] _30573 = {_0, _5310} + {_0, _7357};
  wire [2:0] _30574 = {_0, _30572} + {_0, _30573};
  wire [1:0] _30575 = {_0, _9406} + {_0, _11453};
  wire [3:0] _30576 = {_0, _30574} + {_0, _0, _30575};
  wire _30577 = _12301 < _30576;
  wire _30578 = r17 ^ _30577;
  wire _30579 = _12298 ? coded_block[17] : r17;
  wire _30580 = _12296 ? _30578 : _30579;
  always @ (posedge reset or posedge clock) if (reset) r17 <= 1'd0; else if (_12300) r17 <= _30580;
  wire [1:0] _30581 = {_0, _1247} + {_0, _3294};
  wire [1:0] _30582 = {_0, _5342} + {_0, _7389};
  wire [2:0] _30583 = {_0, _30581} + {_0, _30582};
  wire [1:0] _30584 = {_0, _9438} + {_0, _11485};
  wire [3:0] _30585 = {_0, _30583} + {_0, _0, _30584};
  wire _30586 = _12301 < _30585;
  wire _30587 = r16 ^ _30586;
  wire _30588 = _12298 ? coded_block[16] : r16;
  wire _30589 = _12296 ? _30587 : _30588;
  always @ (posedge reset or posedge clock) if (reset) r16 <= 1'd0; else if (_12300) r16 <= _30589;
  wire [1:0] _30590 = {_0, _1278} + {_0, _3325};
  wire [1:0] _30591 = {_0, _5373} + {_0, _7420};
  wire [2:0] _30592 = {_0, _30590} + {_0, _30591};
  wire [1:0] _30593 = {_0, _9469} + {_0, _11516};
  wire [3:0] _30594 = {_0, _30592} + {_0, _0, _30593};
  wire _30595 = _12301 < _30594;
  wire _30596 = r15 ^ _30595;
  wire _30597 = _12298 ? coded_block[15] : r15;
  wire _30598 = _12296 ? _30596 : _30597;
  always @ (posedge reset or posedge clock) if (reset) r15 <= 1'd0; else if (_12300) r15 <= _30598;
  wire [1:0] _30599 = {_0, _1312} + {_0, _3359};
  wire [1:0] _30600 = {_0, _5407} + {_0, _7454};
  wire [2:0] _30601 = {_0, _30599} + {_0, _30600};
  wire [1:0] _30602 = {_0, _9503} + {_0, _11550};
  wire [3:0] _30603 = {_0, _30601} + {_0, _0, _30602};
  wire _30604 = _12301 < _30603;
  wire _30605 = r14 ^ _30604;
  wire _30606 = _12298 ? coded_block[14] : r14;
  wire _30607 = _12296 ? _30605 : _30606;
  always @ (posedge reset or posedge clock) if (reset) r14 <= 1'd0; else if (_12300) r14 <= _30607;
  wire [1:0] _30608 = {_0, _1343} + {_0, _3390};
  wire [1:0] _30609 = {_0, _5438} + {_0, _7485};
  wire [2:0] _30610 = {_0, _30608} + {_0, _30609};
  wire [1:0] _30611 = {_0, _9534} + {_0, _11581};
  wire [3:0] _30612 = {_0, _30610} + {_0, _0, _30611};
  wire _30613 = _12301 < _30612;
  wire _30614 = r13 ^ _30613;
  wire _30615 = _12298 ? coded_block[13] : r13;
  wire _30616 = _12296 ? _30614 : _30615;
  always @ (posedge reset or posedge clock) if (reset) r13 <= 1'd0; else if (_12300) r13 <= _30616;
  wire [1:0] _30617 = {_0, _1375} + {_0, _3422};
  wire [1:0] _30618 = {_0, _5470} + {_0, _7517};
  wire [2:0] _30619 = {_0, _30617} + {_0, _30618};
  wire [1:0] _30620 = {_0, _9566} + {_0, _11613};
  wire [3:0] _30621 = {_0, _30619} + {_0, _0, _30620};
  wire _30622 = _12301 < _30621;
  wire _30623 = r12 ^ _30622;
  wire _30624 = _12298 ? coded_block[12] : r12;
  wire _30625 = _12296 ? _30623 : _30624;
  always @ (posedge reset or posedge clock) if (reset) r12 <= 1'd0; else if (_12300) r12 <= _30625;
  wire [1:0] _30626 = {_0, _1439} + {_0, _3486};
  wire [1:0] _30627 = {_0, _5534} + {_0, _7581};
  wire [2:0] _30628 = {_0, _30626} + {_0, _30627};
  wire [1:0] _30629 = {_0, _9630} + {_0, _11677};
  wire [3:0] _30630 = {_0, _30628} + {_0, _0, _30629};
  wire _30631 = _12301 < _30630;
  wire _30632 = r11 ^ _30631;
  wire _30633 = _12298 ? coded_block[11] : r11;
  wire _30634 = _12296 ? _30632 : _30633;
  always @ (posedge reset or posedge clock) if (reset) r11 <= 1'd0; else if (_12300) r11 <= _30634;
  wire [1:0] _30635 = {_0, _1470} + {_0, _3517};
  wire [1:0] _30636 = {_0, _5565} + {_0, _7612};
  wire [2:0] _30637 = {_0, _30635} + {_0, _30636};
  wire [1:0] _30638 = {_0, _9661} + {_0, _11708};
  wire [3:0] _30639 = {_0, _30637} + {_0, _0, _30638};
  wire _30640 = _12301 < _30639;
  wire _30641 = r10 ^ _30640;
  wire _30642 = _12298 ? coded_block[10] : r10;
  wire _30643 = _12296 ? _30641 : _30642;
  always @ (posedge reset or posedge clock) if (reset) r10 <= 1'd0; else if (_12300) r10 <= _30643;
  wire [1:0] _30644 = {_0, _1502} + {_0, _3549};
  wire [1:0] _30645 = {_0, _5597} + {_0, _7644};
  wire [2:0] _30646 = {_0, _30644} + {_0, _30645};
  wire [1:0] _30647 = {_0, _9693} + {_0, _11740};
  wire [3:0] _30648 = {_0, _30646} + {_0, _0, _30647};
  wire _30649 = _12301 < _30648;
  wire _30650 = r9 ^ _30649;
  wire _30651 = _12298 ? coded_block[9] : r9;
  wire _30652 = _12296 ? _30650 : _30651;
  always @ (posedge reset or posedge clock) if (reset) r9 <= 1'd0; else if (_12300) r9 <= _30652;
  wire [1:0] _30653 = {_0, _1533} + {_0, _3580};
  wire [1:0] _30654 = {_0, _5628} + {_0, _7675};
  wire [2:0] _30655 = {_0, _30653} + {_0, _30654};
  wire [1:0] _30656 = {_0, _9724} + {_0, _11771};
  wire [3:0] _30657 = {_0, _30655} + {_0, _0, _30656};
  wire _30658 = _12301 < _30657;
  wire _30659 = r8 ^ _30658;
  wire _30660 = _12298 ? coded_block[8] : r8;
  wire _30661 = _12296 ? _30659 : _30660;
  always @ (posedge reset or posedge clock) if (reset) r8 <= 1'd0; else if (_12300) r8 <= _30661;
  wire [1:0] _30662 = {_0, _1568} + {_0, _3615};
  wire [1:0] _30663 = {_0, _5663} + {_0, _7710};
  wire [2:0] _30664 = {_0, _30662} + {_0, _30663};
  wire [1:0] _30665 = {_0, _9759} + {_0, _11806};
  wire [3:0] _30666 = {_0, _30664} + {_0, _0, _30665};
  wire _30667 = _12301 < _30666;
  wire _30668 = r7 ^ _30667;
  wire _30669 = _12298 ? coded_block[7] : r7;
  wire _30670 = _12296 ? _30668 : _30669;
  always @ (posedge reset or posedge clock) if (reset) r7 <= 1'd0; else if (_12300) r7 <= _30670;
  wire [1:0] _30671 = {_0, _1599} + {_0, _3646};
  wire [1:0] _30672 = {_0, _5694} + {_0, _7741};
  wire [2:0] _30673 = {_0, _30671} + {_0, _30672};
  wire [1:0] _30674 = {_0, _9790} + {_0, _11837};
  wire [3:0] _30675 = {_0, _30673} + {_0, _0, _30674};
  wire _30676 = _12301 < _30675;
  wire _30677 = r6 ^ _30676;
  wire _30678 = _12298 ? coded_block[6] : r6;
  wire _30679 = _12296 ? _30677 : _30678;
  always @ (posedge reset or posedge clock) if (reset) r6 <= 1'd0; else if (_12300) r6 <= _30679;
  wire [1:0] _30680 = {_0, _1631} + {_0, _3678};
  wire [1:0] _30681 = {_0, _5726} + {_0, _7773};
  wire [2:0] _30682 = {_0, _30680} + {_0, _30681};
  wire [1:0] _30683 = {_0, _9822} + {_0, _11869};
  wire [3:0] _30684 = {_0, _30682} + {_0, _0, _30683};
  wire _30685 = _12301 < _30684;
  wire _30686 = r5 ^ _30685;
  wire _30687 = _12298 ? coded_block[5] : r5;
  wire _30688 = _12296 ? _30686 : _30687;
  always @ (posedge reset or posedge clock) if (reset) r5 <= 1'd0; else if (_12300) r5 <= _30688;
  wire [1:0] _30689 = {_0, _1662} + {_0, _3709};
  wire [1:0] _30690 = {_0, _5757} + {_0, _7804};
  wire [2:0] _30691 = {_0, _30689} + {_0, _30690};
  wire [1:0] _30692 = {_0, _9853} + {_0, _11900};
  wire [3:0] _30693 = {_0, _30691} + {_0, _0, _30692};
  wire _30694 = _12301 < _30693;
  wire _30695 = r4 ^ _30694;
  wire _30696 = _12298 ? coded_block[4] : r4;
  wire _30697 = _12296 ? _30695 : _30696;
  always @ (posedge reset or posedge clock) if (reset) r4 <= 1'd0; else if (_12300) r4 <= _30697;
  wire [1:0] _30698 = {_0, _1726} + {_0, _3773};
  wire [1:0] _30699 = {_0, _5821} + {_0, _7868};
  wire [2:0] _30700 = {_0, _30698} + {_0, _30699};
  wire [1:0] _30701 = {_0, _9917} + {_0, _11964};
  wire [3:0] _30702 = {_0, _30700} + {_0, _0, _30701};
  wire _30703 = _12301 < _30702;
  wire _30704 = r3 ^ _30703;
  wire _30705 = _12298 ? coded_block[3] : r3;
  wire _30706 = _12296 ? _30704 : _30705;
  always @ (posedge reset or posedge clock) if (reset) r3 <= 1'd0; else if (_12300) r3 <= _30706;
  wire [1:0] _30707 = {_0, _1758} + {_0, _3805};
  wire [1:0] _30708 = {_0, _5853} + {_0, _7900};
  wire [2:0] _30709 = {_0, _30707} + {_0, _30708};
  wire [1:0] _30710 = {_0, _9949} + {_0, _11996};
  wire [3:0] _30711 = {_0, _30709} + {_0, _0, _30710};
  wire _30712 = _12301 < _30711;
  wire _30713 = r2 ^ _30712;
  wire _30714 = _12298 ? coded_block[2] : r2;
  wire _30715 = _12296 ? _30713 : _30714;
  always @ (posedge reset or posedge clock) if (reset) r2 <= 1'd0; else if (_12300) r2 <= _30715;
  wire [1:0] _30716 = {_0, _1789} + {_0, _3836};
  wire [1:0] _30717 = {_0, _5884} + {_0, _7931};
  wire [2:0] _30718 = {_0, _30716} + {_0, _30717};
  wire [1:0] _30719 = {_0, _9980} + {_0, _12027};
  wire [3:0] _30720 = {_0, _30718} + {_0, _0, _30719};
  wire _30721 = _12301 < _30720;
  wire _30722 = r1 ^ _30721;
  wire _30723 = _12298 ? coded_block[1] : r1;
  wire _30724 = _12296 ? _30722 : _30723;
  always @ (posedge reset or posedge clock) if (reset) r1 <= 1'd0; else if (_12300) r1 <= _30724;
  wire [1:0] _30725 = {_0, _1823} + {_0, _3870};
  wire [1:0] _30726 = {_0, _5918} + {_0, _7965};
  wire [2:0] _30727 = {_0, _30725} + {_0, _30726};
  wire [1:0] _30728 = {_0, _10014} + {_0, _12061};
  wire [3:0] _30729 = {_0, _30727} + {_0, _0, _30728};
  wire _30730 = _12301 < _30729;
  wire _30731 = r0 ^ _30730;
  wire _30732 = _12298 ? coded_block[0] : r0;
  wire _30733 = _12296 ? _30731 : _30732;
  always @ (posedge reset or posedge clock) if (reset) r0 <= 1'd0; else if (_12300) r0 <= _30733;
  assign decoded = _12291;
  assign decoded_block = {r2047, r2046, r2045, r2044, r2043, r2042, r2041, r2040, r2039, r2038, r2037, r2036, r2035, r2034, r2033, r2032, r2031, r2030, r2029, r2028, r2027, r2026, r2025, r2024, r2023, r2022, r2021, r2020, r2019, r2018, r2017, r2016, r2015, r2014, r2013, r2012, r2011, r2010, r2009, r2008, r2007, r2006, r2005, r2004, r2003, r2002, r2001, r2000, r1999, r1998, r1997, r1996, r1995, r1994, r1993, r1992, r1991, r1990, r1989, r1988, r1987, r1986, r1985, r1984, r1983, r1982, r1981, r1980, r1979, r1978, r1977, r1976, r1975, r1974, r1973, r1972, r1971, r1970, r1969, r1968, r1967, r1966, r1965, r1964, r1963, r1962, r1961, r1960, r1959, r1958, r1957, r1956, r1955, r1954, r1953, r1952, r1951, r1950, r1949, r1948, r1947, r1946, r1945, r1944, r1943, r1942, r1941, r1940, r1939, r1938, r1937, r1936, r1935, r1934, r1933, r1932, r1931, r1930, r1929, r1928, r1927, r1926, r1925, r1924, r1923, r1922, r1921, r1920, r1919, r1918, r1917, r1916, r1915, r1914, r1913, r1912, r1911, r1910, r1909, r1908, r1907, r1906, r1905, r1904, r1903, r1902, r1901, r1900, r1899, r1898, r1897, r1896, r1895, r1894, r1893, r1892, r1891, r1890, r1889, r1888, r1887, r1886, r1885, r1884, r1883, r1882, r1881, r1880, r1879, r1878, r1877, r1876, r1875, r1874, r1873, r1872, r1871, r1870, r1869, r1868, r1867, r1866, r1865, r1864, r1863, r1862, r1861, r1860, r1859, r1858, r1857, r1856, r1855, r1854, r1853, r1852, r1851, r1850, r1849, r1848, r1847, r1846, r1845, r1844, r1843, r1842, r1841, r1840, r1839, r1838, r1837, r1836, r1835, r1834, r1833, r1832, r1831, r1830, r1829, r1828, r1827, r1826, r1825, r1824, r1823, r1822, r1821, r1820, r1819, r1818, r1817, r1816, r1815, r1814, r1813, r1812, r1811, r1810, r1809, r1808, r1807, r1806, r1805, r1804, r1803, r1802, r1801, r1800, r1799, r1798, r1797, r1796, r1795, r1794, r1793, r1792, r1791, r1790, r1789, r1788, r1787, r1786, r1785, r1784, r1783, r1782, r1781, r1780, r1779, r1778, r1777, r1776, r1775, r1774, r1773, r1772, r1771, r1770, r1769, r1768, r1767, r1766, r1765, r1764, r1763, r1762, r1761, r1760, r1759, r1758, r1757, r1756, r1755, r1754, r1753, r1752, r1751, r1750, r1749, r1748, r1747, r1746, r1745, r1744, r1743, r1742, r1741, r1740, r1739, r1738, r1737, r1736, r1735, r1734, r1733, r1732, r1731, r1730, r1729, r1728, r1727, r1726, r1725, r1724, r1723, r1722, r1721, r1720, r1719, r1718, r1717, r1716, r1715, r1714, r1713, r1712, r1711, r1710, r1709, r1708, r1707, r1706, r1705, r1704, r1703, r1702, r1701, r1700, r1699, r1698, r1697, r1696, r1695, r1694, r1693, r1692, r1691, r1690, r1689, r1688, r1687, r1686, r1685, r1684, r1683, r1682, r1681, r1680, r1679, r1678, r1677, r1676, r1675, r1674, r1673, r1672, r1671, r1670, r1669, r1668, r1667, r1666, r1665, r1664, r1663, r1662, r1661, r1660, r1659, r1658, r1657, r1656, r1655, r1654, r1653, r1652, r1651, r1650, r1649, r1648, r1647, r1646, r1645, r1644, r1643, r1642, r1641, r1640, r1639, r1638, r1637, r1636, r1635, r1634, r1633, r1632, r1631, r1630, r1629, r1628, r1627, r1626, r1625, r1624, r1623, r1622, r1621, r1620, r1619, r1618, r1617, r1616, r1615, r1614, r1613, r1612, r1611, r1610, r1609, r1608, r1607, r1606, r1605, r1604, r1603, r1602, r1601, r1600, r1599, r1598, r1597, r1596, r1595, r1594, r1593, r1592, r1591, r1590, r1589, r1588, r1587, r1586, r1585, r1584, r1583, r1582, r1581, r1580, r1579, r1578, r1577, r1576, r1575, r1574, r1573, r1572, r1571, r1570, r1569, r1568, r1567, r1566, r1565, r1564, r1563, r1562, r1561, r1560, r1559, r1558, r1557, r1556, r1555, r1554, r1553, r1552, r1551, r1550, r1549, r1548, r1547, r1546, r1545, r1544, r1543, r1542, r1541, r1540, r1539, r1538, r1537, r1536, r1535, r1534, r1533, r1532, r1531, r1530, r1529, r1528, r1527, r1526, r1525, r1524, r1523, r1522, r1521, r1520, r1519, r1518, r1517, r1516, r1515, r1514, r1513, r1512, r1511, r1510, r1509, r1508, r1507, r1506, r1505, r1504, r1503, r1502, r1501, r1500, r1499, r1498, r1497, r1496, r1495, r1494, r1493, r1492, r1491, r1490, r1489, r1488, r1487, r1486, r1485, r1484, r1483, r1482, r1481, r1480, r1479, r1478, r1477, r1476, r1475, r1474, r1473, r1472, r1471, r1470, r1469, r1468, r1467, r1466, r1465, r1464, r1463, r1462, r1461, r1460, r1459, r1458, r1457, r1456, r1455, r1454, r1453, r1452, r1451, r1450, r1449, r1448, r1447, r1446, r1445, r1444, r1443, r1442, r1441, r1440, r1439, r1438, r1437, r1436, r1435, r1434, r1433, r1432, r1431, r1430, r1429, r1428, r1427, r1426, r1425, r1424, r1423, r1422, r1421, r1420, r1419, r1418, r1417, r1416, r1415, r1414, r1413, r1412, r1411, r1410, r1409, r1408, r1407, r1406, r1405, r1404, r1403, r1402, r1401, r1400, r1399, r1398, r1397, r1396, r1395, r1394, r1393, r1392, r1391, r1390, r1389, r1388, r1387, r1386, r1385, r1384, r1383, r1382, r1381, r1380, r1379, r1378, r1377, r1376, r1375, r1374, r1373, r1372, r1371, r1370, r1369, r1368, r1367, r1366, r1365, r1364, r1363, r1362, r1361, r1360, r1359, r1358, r1357, r1356, r1355, r1354, r1353, r1352, r1351, r1350, r1349, r1348, r1347, r1346, r1345, r1344, r1343, r1342, r1341, r1340, r1339, r1338, r1337, r1336, r1335, r1334, r1333, r1332, r1331, r1330, r1329, r1328, r1327, r1326, r1325, r1324, r1323, r1322, r1321, r1320, r1319, r1318, r1317, r1316, r1315, r1314, r1313, r1312, r1311, r1310, r1309, r1308, r1307, r1306, r1305, r1304, r1303, r1302, r1301, r1300, r1299, r1298, r1297, r1296, r1295, r1294, r1293, r1292, r1291, r1290, r1289, r1288, r1287, r1286, r1285, r1284, r1283, r1282, r1281, r1280, r1279, r1278, r1277, r1276, r1275, r1274, r1273, r1272, r1271, r1270, r1269, r1268, r1267, r1266, r1265, r1264, r1263, r1262, r1261, r1260, r1259, r1258, r1257, r1256, r1255, r1254, r1253, r1252, r1251, r1250, r1249, r1248, r1247, r1246, r1245, r1244, r1243, r1242, r1241, r1240, r1239, r1238, r1237, r1236, r1235, r1234, r1233, r1232, r1231, r1230, r1229, r1228, r1227, r1226, r1225, r1224, r1223, r1222, r1221, r1220, r1219, r1218, r1217, r1216, r1215, r1214, r1213, r1212, r1211, r1210, r1209, r1208, r1207, r1206, r1205, r1204, r1203, r1202, r1201, r1200, r1199, r1198, r1197, r1196, r1195, r1194, r1193, r1192, r1191, r1190, r1189, r1188, r1187, r1186, r1185, r1184, r1183, r1182, r1181, r1180, r1179, r1178, r1177, r1176, r1175, r1174, r1173, r1172, r1171, r1170, r1169, r1168, r1167, r1166, r1165, r1164, r1163, r1162, r1161, r1160, r1159, r1158, r1157, r1156, r1155, r1154, r1153, r1152, r1151, r1150, r1149, r1148, r1147, r1146, r1145, r1144, r1143, r1142, r1141, r1140, r1139, r1138, r1137, r1136, r1135, r1134, r1133, r1132, r1131, r1130, r1129, r1128, r1127, r1126, r1125, r1124, r1123, r1122, r1121, r1120, r1119, r1118, r1117, r1116, r1115, r1114, r1113, r1112, r1111, r1110, r1109, r1108, r1107, r1106, r1105, r1104, r1103, r1102, r1101, r1100, r1099, r1098, r1097, r1096, r1095, r1094, r1093, r1092, r1091, r1090, r1089, r1088, r1087, r1086, r1085, r1084, r1083, r1082, r1081, r1080, r1079, r1078, r1077, r1076, r1075, r1074, r1073, r1072, r1071, r1070, r1069, r1068, r1067, r1066, r1065, r1064, r1063, r1062, r1061, r1060, r1059, r1058, r1057, r1056, r1055, r1054, r1053, r1052, r1051, r1050, r1049, r1048, r1047, r1046, r1045, r1044, r1043, r1042, r1041, r1040, r1039, r1038, r1037, r1036, r1035, r1034, r1033, r1032, r1031, r1030, r1029, r1028, r1027, r1026, r1025, r1024, r1023, r1022, r1021, r1020, r1019, r1018, r1017, r1016, r1015, r1014, r1013, r1012, r1011, r1010, r1009, r1008, r1007, r1006, r1005, r1004, r1003, r1002, r1001, r1000, r999, r998, r997, r996, r995, r994, r993, r992, r991, r990, r989, r988, r987, r986, r985, r984, r983, r982, r981, r980, r979, r978, r977, r976, r975, r974, r973, r972, r971, r970, r969, r968, r967, r966, r965, r964, r963, r962, r961, r960, r959, r958, r957, r956, r955, r954, r953, r952, r951, r950, r949, r948, r947, r946, r945, r944, r943, r942, r941, r940, r939, r938, r937, r936, r935, r934, r933, r932, r931, r930, r929, r928, r927, r926, r925, r924, r923, r922, r921, r920, r919, r918, r917, r916, r915, r914, r913, r912, r911, r910, r909, r908, r907, r906, r905, r904, r903, r902, r901, r900, r899, r898, r897, r896, r895, r894, r893, r892, r891, r890, r889, r888, r887, r886, r885, r884, r883, r882, r881, r880, r879, r878, r877, r876, r875, r874, r873, r872, r871, r870, r869, r868, r867, r866, r865, r864, r863, r862, r861, r860, r859, r858, r857, r856, r855, r854, r853, r852, r851, r850, r849, r848, r847, r846, r845, r844, r843, r842, r841, r840, r839, r838, r837, r836, r835, r834, r833, r832, r831, r830, r829, r828, r827, r826, r825, r824, r823, r822, r821, r820, r819, r818, r817, r816, r815, r814, r813, r812, r811, r810, r809, r808, r807, r806, r805, r804, r803, r802, r801, r800, r799, r798, r797, r796, r795, r794, r793, r792, r791, r790, r789, r788, r787, r786, r785, r784, r783, r782, r781, r780, r779, r778, r777, r776, r775, r774, r773, r772, r771, r770, r769, r768, r767, r766, r765, r764, r763, r762, r761, r760, r759, r758, r757, r756, r755, r754, r753, r752, r751, r750, r749, r748, r747, r746, r745, r744, r743, r742, r741, r740, r739, r738, r737, r736, r735, r734, r733, r732, r731, r730, r729, r728, r727, r726, r725, r724, r723, r722, r721, r720, r719, r718, r717, r716, r715, r714, r713, r712, r711, r710, r709, r708, r707, r706, r705, r704, r703, r702, r701, r700, r699, r698, r697, r696, r695, r694, r693, r692, r691, r690, r689, r688, r687, r686, r685, r684, r683, r682, r681, r680, r679, r678, r677, r676, r675, r674, r673, r672, r671, r670, r669, r668, r667, r666, r665, r664, r663, r662, r661, r660, r659, r658, r657, r656, r655, r654, r653, r652, r651, r650, r649, r648, r647, r646, r645, r644, r643, r642, r641, r640, r639, r638, r637, r636, r635, r634, r633, r632, r631, r630, r629, r628, r627, r626, r625, r624, r623, r622, r621, r620, r619, r618, r617, r616, r615, r614, r613, r612, r611, r610, r609, r608, r607, r606, r605, r604, r603, r602, r601, r600, r599, r598, r597, r596, r595, r594, r593, r592, r591, r590, r589, r588, r587, r586, r585, r584, r583, r582, r581, r580, r579, r578, r577, r576, r575, r574, r573, r572, r571, r570, r569, r568, r567, r566, r565, r564, r563, r562, r561, r560, r559, r558, r557, r556, r555, r554, r553, r552, r551, r550, r549, r548, r547, r546, r545, r544, r543, r542, r541, r540, r539, r538, r537, r536, r535, r534, r533, r532, r531, r530, r529, r528, r527, r526, r525, r524, r523, r522, r521, r520, r519, r518, r517, r516, r515, r514, r513, r512, r511, r510, r509, r508, r507, r506, r505, r504, r503, r502, r501, r500, r499, r498, r497, r496, r495, r494, r493, r492, r491, r490, r489, r488, r487, r486, r485, r484, r483, r482, r481, r480, r479, r478, r477, r476, r475, r474, r473, r472, r471, r470, r469, r468, r467, r466, r465, r464, r463, r462, r461, r460, r459, r458, r457, r456, r455, r454, r453, r452, r451, r450, r449, r448, r447, r446, r445, r444, r443, r442, r441, r440, r439, r438, r437, r436, r435, r434, r433, r432, r431, r430, r429, r428, r427, r426, r425, r424, r423, r422, r421, r420, r419, r418, r417, r416, r415, r414, r413, r412, r411, r410, r409, r408, r407, r406, r405, r404, r403, r402, r401, r400, r399, r398, r397, r396, r395, r394, r393, r392, r391, r390, r389, r388, r387, r386, r385, r384, r383, r382, r381, r380, r379, r378, r377, r376, r375, r374, r373, r372, r371, r370, r369, r368, r367, r366, r365, r364, r363, r362, r361, r360, r359, r358, r357, r356, r355, r354, r353, r352, r351, r350, r349, r348, r347, r346, r345, r344, r343, r342, r341, r340, r339, r338, r337, r336, r335, r334, r333, r332, r331, r330, r329, r328, r327, r326, r325, r324, r323, r322, r321, r320, r319, r318, r317, r316, r315, r314, r313, r312, r311, r310, r309, r308, r307, r306, r305, r304, r303, r302, r301, r300, r299, r298, r297, r296, r295, r294, r293, r292, r291, r290, r289, r288, r287, r286, r285, r284, r283, r282, r281, r280, r279, r278, r277, r276, r275, r274, r273, r272, r271, r270, r269, r268, r267, r266, r265, r264, r263, r262, r261, r260, r259, r258, r257, r256, r255, r254, r253, r252, r251, r250, r249, r248, r247, r246, r245, r244, r243, r242, r241, r240, r239, r238, r237, r236, r235, r234, r233, r232, r231, r230, r229, r228, r227, r226, r225, r224, r223, r222, r221, r220, r219, r218, r217, r216, r215, r214, r213, r212, r211, r210, r209, r208, r207, r206, r205, r204, r203, r202, r201, r200, r199, r198, r197, r196, r195, r194, r193, r192, r191, r190, r189, r188, r187, r186, r185, r184, r183, r182, r181, r180, r179, r178, r177, r176, r175, r174, r173, r172, r171, r170, r169, r168, r167, r166, r165, r164, r163, r162, r161, r160, r159, r158, r157, r156, r155, r154, r153, r152, r151, r150, r149, r148, r147, r146, r145, r144, r143, r142, r141, r140, r139, r138, r137, r136, r135, r134, r133, r132, r131, r130, r129, r128, r127, r126, r125, r124, r123, r122, r121, r120, r119, r118, r117, r116, r115, r114, r113, r112, r111, r110, r109, r108, r107, r106, r105, r104, r103, r102, r101, r100, r99, r98, r97, r96, r95, r94, r93, r92, r91, r90, r89, r88, r87, r86, r85, r84, r83, r82, r81, r80, r79, r78, r77, r76, r75, r74, r73, r72, r71, r70, r69, r68, r67, r66, r65, r64, r63, r62, r61, r60, r59, r58, r57, r56, r55, r54, r53, r52, r51, r50, r49, r48, r47, r46, r45, r44, r43, r42, r41, r40, r39, r38, r37, r36, r35, r34, r33, r32, r31, r30, r29, r28, r27, r26, r25, r24, r23, r22, r21, r20, r19, r18, r17, r16, r15, r14, r13, r12, r11, r10, r9, r8, r7, r6, r5, r4, r3, r2, r1, r0};
endmodule

